PK
     ˡ�Z�`�* *    cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_0":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_0":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_1":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_1":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_2":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_2":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_3":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_3":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_4":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_4":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_5":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_5":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_6":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_6":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_7":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_7":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_8":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_8":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_9":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_9":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_10":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_10":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_11":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_11":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_12":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_12":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_13":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_13":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_14":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_14":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_15":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_15":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_16":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_16":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_17":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_17":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_18":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_18":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_19":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_19":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_20":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_20":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_21":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_21":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_22":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_22":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_23":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_23":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_24":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_24":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_25":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_25":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_26":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_26":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_27":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_27":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_28":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_28":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_29":[],"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_29":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_0_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_0_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_0_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_0_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_1_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_1_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_1_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_1_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_2_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_2_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_2_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_2_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_3_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_3_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_3_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_3_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_4_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_4_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_4_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_4_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_5_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_5_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_5_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_5_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_6_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_6_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_6_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_6_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_7_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_7_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_7_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_7_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_8_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_8_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_8_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_8_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_9_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_9_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_9_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_9_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_10_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_10_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_10_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_10_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_11_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_11_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_11_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_11_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_12_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_12_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_12_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_12_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_13_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_13_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_13_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_13_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_14_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_14_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_14_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_14_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_15_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_15_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_15_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_15_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_16_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_16_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_16_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_16_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_17_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_17_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_17_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_17_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_18_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_18_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_18_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_18_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_19_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_19_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_19_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_19_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_20_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_20_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_20_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_20_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_21_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_21_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_21_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_21_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_22_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_22_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_22_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_22_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_23_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_23_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_23_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_23_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_24_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_24_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_24_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_24_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_25_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_25_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_25_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_25_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_26_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_26_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_26_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_26_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_27_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_27_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_27_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_27_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_28_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_28_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_28_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_28_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_29_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_29_polarity-neg":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_29_polarity-pos":[],"pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_29_polarity-neg":[],"pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_0":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_0"],"pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_1":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_1"],"pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_0":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_5"],"pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_1":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_6"],"pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_0":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_5"],"pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_1":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_6"],"pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_0":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_0"],"pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_1":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_1"],"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_0":["pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_0","pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_0"],"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_1":["pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_1","pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_1"],"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_2":["pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_1"],"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_3":["pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_0","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_18"],"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_4":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19"],"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_5":["pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_0","pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_0"],"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_6":["pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_1","pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_1"],"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_7":[],"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_8":[],"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_9":[],"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_10":[],"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_11":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_15"],"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_12":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_14"],"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_13":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_13"],"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_14":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_11"],"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_15":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_10"],"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_16":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_12"],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_0":[],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_1":[],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_2":[],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_3":[],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_4":[],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_5":[],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_6":[],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_7":[],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_8":[],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_9":[],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_10":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_15"],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_11":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_14"],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_12":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_16"],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_13":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_13"],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_14":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_12"],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_15":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_11"],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_16":[],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_17":[],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_18":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_3"],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_4","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_0","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_1"],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_20":[],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_21":[],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_22":[],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_23":[],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_24":[],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_25":["pin-type-component_362ae36f-3285-42bd-a265-880763af6269_2"],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_26":["pin-type-component_362ae36f-3285-42bd-a265-880763af6269_1"],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_27":["pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_0"],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28":["pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_2","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_3"],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_29":[],"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_30":[],"pin-type-component_362ae36f-3285-42bd-a265-880763af6269_0":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19"],"pin-type-component_362ae36f-3285-42bd-a265-880763af6269_1":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_26"],"pin-type-component_362ae36f-3285-42bd-a265-880763af6269_2":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_25"],"pin-type-component_362ae36f-3285-42bd-a265-880763af6269_3":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28"],"pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_0":[],"pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_1":[],"pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_2":[],"pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_3":[],"pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_4":[],"pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_5":[],"pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_6":[],"pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_7":[],"pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_8":[],"pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_9":[],"pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_10":[],"pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_11":[],"pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_12":[],"pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_13":[],"pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_14":[],"pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_15":[],"pin-type-component_c4a184a4-3697-449d-9903-a666adf64026_0":[],"pin-type-component_c4a184a4-3697-449d-9903-a666adf64026_1":[],"pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_0":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_27"],"pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_1":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19"],"pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_2":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28"],"pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_0":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_3"],"pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_1":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_2"]},"pin_to_color":{"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_0":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_0":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_1":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_1":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_2":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_2":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_3":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_3":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_4":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_4":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_5":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_5":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_6":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_6":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_7":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_7":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_8":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_8":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_9":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_9":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_10":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_10":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_11":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_11":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_12":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_12":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_13":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_13":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_14":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_14":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_15":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_15":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_16":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_16":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_17":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_17":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_18":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_18":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_19":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_19":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_20":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_20":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_21":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_21":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_22":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_22":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_23":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_23":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_24":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_24":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_25":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_25":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_26":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_26":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_27":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_27":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_28":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_28":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_29":"#000000","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_29":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_0_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_0_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_0_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_0_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_1_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_1_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_1_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_1_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_2_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_2_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_2_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_2_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_3_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_3_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_3_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_3_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_4_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_4_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_4_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_4_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_5_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_5_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_5_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_5_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_6_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_6_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_6_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_6_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_7_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_7_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_7_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_7_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_8_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_8_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_8_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_8_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_9_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_9_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_9_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_9_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_10_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_10_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_10_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_10_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_11_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_11_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_11_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_11_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_12_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_12_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_12_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_12_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_13_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_13_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_13_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_13_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_14_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_14_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_14_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_14_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_15_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_15_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_15_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_15_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_16_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_16_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_16_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_16_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_17_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_17_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_17_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_17_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_18_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_18_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_18_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_18_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_19_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_19_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_19_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_19_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_20_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_20_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_20_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_20_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_21_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_21_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_21_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_21_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_22_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_22_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_22_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_22_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_23_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_23_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_23_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_23_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_24_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_24_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_24_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_24_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_25_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_25_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_25_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_25_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_26_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_26_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_26_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_26_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_27_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_27_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_27_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_27_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_28_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_28_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_28_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_28_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_29_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_29_polarity-neg":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_29_polarity-pos":"#000000","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_29_polarity-neg":"#000000","pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_0":"#010067","pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_1":"#9E008E","pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_0":"#0E4CA1","pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_1":"#FFE502","pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_0":"#0E4CA1","pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_1":"#FFE502","pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_0":"#010067","pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_1":"#9E008E","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_0":"#010067","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_1":"#9E008E","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_2":"#B500FF","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_3":"#FF74A3","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_4":"#968AE8","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_5":"#0E4CA1","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_6":"#FFE502","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_7":"#000000","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_8":"#000000","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_9":"#000000","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_10":"#000000","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_11":"#98FF52","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_12":"#A75740","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_13":"#01FFFE","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_14":"#FE8900","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_15":"#BDC6FF","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_16":"#BB8800","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_0":"#000000","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_1":"#000000","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_2":"#000000","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_3":"#000000","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_4":"#000000","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_5":"#000000","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_6":"#000000","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_7":"#000000","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_8":"#000000","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_9":"#000000","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_10":"#BDC6FF","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_11":"#FE8900","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_12":"#BB8800","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_13":"#01FFFE","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_14":"#A75740","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_15":"#98FF52","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_16":"#000000","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_17":"#000000","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_18":"#FF74A3","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19":"#968AE8","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_20":"#000000","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_21":"#000000","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_22":"#000000","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_23":"#000000","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_24":"#000000","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_25":"#FFA6FE","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_26":"#A5FFD2","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_27":"#774D00","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28":"#7544B1","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_29":"#000000","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_30":"#000000","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_0":"#968AE8","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_1":"#A5FFD2","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_2":"#FFA6FE","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_3":"#7544B1","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_0":"#000000","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_1":"#000000","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_2":"#000000","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_3":"#000000","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_4":"#000000","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_5":"#000000","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_6":"#000000","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_7":"#000000","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_8":"#000000","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_9":"#000000","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_10":"#000000","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_11":"#000000","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_12":"#000000","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_13":"#000000","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_14":"#000000","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_15":"#000000","pin-type-component_c4a184a4-3697-449d-9903-a666adf64026_0":"#000000","pin-type-component_c4a184a4-3697-449d-9903-a666adf64026_1":"#000000","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_0":"#774D00","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_1":"#968AE8","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_2":"#7544B1","pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_0":"#FF74A3","pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_1":"#B500FF"},"pin_to_state":{"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_0":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_0":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_1":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_1":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_2":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_2":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_3":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_3":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_4":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_4":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_5":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_5":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_6":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_6":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_7":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_7":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_8":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_8":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_9":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_9":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_10":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_10":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_11":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_11":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_12":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_12":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_13":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_13":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_14":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_14":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_15":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_15":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_16":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_16":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_17":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_17":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_18":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_18":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_19":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_19":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_20":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_20":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_21":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_21":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_22":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_22":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_23":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_23":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_24":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_24":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_25":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_25":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_26":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_26":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_27":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_27":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_28":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_28":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_29":"neutral","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_29":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_0_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_0_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_0_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_0_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_1_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_1_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_1_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_1_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_2_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_2_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_2_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_2_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_3_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_3_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_3_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_3_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_4_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_4_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_4_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_4_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_5_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_5_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_5_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_5_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_6_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_6_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_6_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_6_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_7_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_7_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_7_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_7_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_8_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_8_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_8_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_8_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_9_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_9_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_9_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_9_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_10_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_10_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_10_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_10_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_11_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_11_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_11_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_11_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_12_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_12_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_12_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_12_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_13_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_13_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_13_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_13_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_14_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_14_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_14_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_14_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_15_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_15_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_15_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_15_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_16_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_16_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_16_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_16_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_17_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_17_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_17_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_17_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_18_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_18_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_18_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_18_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_19_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_19_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_19_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_19_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_20_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_20_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_20_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_20_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_21_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_21_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_21_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_21_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_22_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_22_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_22_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_22_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_23_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_23_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_23_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_23_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_24_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_24_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_24_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_24_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_25_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_25_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_25_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_25_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_26_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_26_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_26_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_26_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_27_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_27_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_27_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_27_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_28_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_28_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_28_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_28_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_29_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_29_polarity-neg":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_29_polarity-pos":"neutral","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_29_polarity-neg":"neutral","pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_0":"neutral","pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_1":"neutral","pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_0":"neutral","pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_1":"neutral","pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_0":"neutral","pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_1":"neutral","pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_0":"neutral","pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_1":"neutral","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_0":"neutral","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_1":"neutral","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_2":"neutral","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_3":"neutral","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_4":"neutral","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_5":"neutral","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_6":"neutral","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_7":"neutral","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_8":"neutral","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_9":"neutral","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_10":"neutral","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_11":"neutral","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_12":"neutral","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_13":"neutral","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_14":"neutral","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_15":"neutral","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_16":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_0":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_1":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_2":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_3":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_4":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_5":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_6":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_7":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_8":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_9":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_10":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_11":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_12":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_13":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_14":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_15":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_16":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_17":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_18":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_20":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_21":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_22":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_23":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_24":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_25":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_26":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_27":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_29":"neutral","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_30":"neutral","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_0":"neutral","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_1":"neutral","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_2":"neutral","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_3":"neutral","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_0":"neutral","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_1":"neutral","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_2":"neutral","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_3":"neutral","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_4":"neutral","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_5":"neutral","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_6":"neutral","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_7":"neutral","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_8":"neutral","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_9":"neutral","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_10":"neutral","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_11":"neutral","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_12":"neutral","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_13":"neutral","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_14":"neutral","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_15":"neutral","pin-type-component_c4a184a4-3697-449d-9903-a666adf64026_0":"neutral","pin-type-component_c4a184a4-3697-449d-9903-a666adf64026_1":"neutral","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_0":"neutral","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_1":"neutral","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_2":"neutral","pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_0":"neutral","pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_1":"neutral"},"next_color_idx":32,"wires_placed_in_order":[["pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_0","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_0"],["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_0","pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_0"],["pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_1","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_1"],["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_1","pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_1"],["pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_0","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_5"],["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_5","pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_0"],["pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_1","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_6"],["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_6","pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_1"],["pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_1","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_2"],["pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_0","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28"],["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_3"],["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_4","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_0"],["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_4","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19"],["pin-type-component_362ae36f-3285-42bd-a265-880763af6269_0","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_1"],["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_11","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_15"],["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_12","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_14"],["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_13","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_13"],["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_14","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_11"],["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_15","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_10"],["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_16","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_12"],["pin-type-component_362ae36f-3285-42bd-a265-880763af6269_1","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_26"],["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_25","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_2"],["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_27","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_3"],["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_27","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_2"],["pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_2","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_0"],["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_27","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_0"],["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_2"],["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_2","pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_1"],["pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_0","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_3"],["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_4","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19"],["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_0"],["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_1"],["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_15","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_11"],["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_14","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_12"],["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_13","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_13"],["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_11","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_14"],["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_15","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_10"],["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_12","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_16"],["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_3","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_18"],["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_2"],["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_3"],["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_26","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_1"],["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_25","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_2"],["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_27","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_0"],["pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_1","pin-type-component_5c94b46d-7fef-4bd1-a0eb-c5c4156d6d12_0"],["pin-type-component_5c94b46d-7fef-4bd1-a0eb-c5c4156d6d12_1","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_2"],["pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_1","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_2"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_0","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_0"]]],[[],[["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_0","pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_0"]]],[[],[["pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_1","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_1"]]],[[],[["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_1","pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_1"]]],[[],[["pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_0","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_5"]]],[[],[["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_5","pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_0"]]],[[],[["pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_1","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_6"]]],[[],[["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_6","pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_1"]]],[[],[["pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_1","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_2"]]],[[],[["pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_0","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28"]]],[[],[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_3"]]],[[],[["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_4","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_0"]]],[[],[["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_4","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19"]]],[[],[["pin-type-component_362ae36f-3285-42bd-a265-880763af6269_0","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_1"]]],[[],[["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_11","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_15"]]],[[],[["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_12","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_14"]]],[[],[["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_13","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_13"]]],[[],[["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_14","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_11"]]],[[],[["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_15","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_10"]]],[[],[["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_16","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_12"]]],[[],[["pin-type-component_362ae36f-3285-42bd-a265-880763af6269_1","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_26"]]],[[],[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_25","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_2"]]],[[],[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_27","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_3"]]],[[],[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_27","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_2"]]],[[],[["pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_2","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_0"]]],[[["pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_0","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_2"]],[]],[[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_27","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_2"]],[]],[[],[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_27","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_0"]]],[[],[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_2"]]],[[["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_2","pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_1"]],[]],[[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_3"]],[]],[[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_4"]],[]],[[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_15","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_11"]],[]],[[["pin-type-component_362ae36f-3285-42bd-a265-880763af6269_0","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_4"]],[]],[[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_14","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_12"]],[]],[[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_13","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_13"]],[]],[[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_11","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_14"]],[]],[[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_10","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_15"]],[]],[[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_12","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_16"]],[]],[[["pin-type-component_362ae36f-3285-42bd-a265-880763af6269_2","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_25"]],[]],[[["pin-type-component_362ae36f-3285-42bd-a265-880763af6269_1","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_26"]],[]],[[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_27","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_0"]],[]],[[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_2"]],[]],[[["pin-type-component_362ae36f-3285-42bd-a265-880763af6269_3","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_27"]],[]],[[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28","pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_0"]],[]],[[["pin-type-component_362ae36f-3285-42bd-a265-880763af6269_0","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_1"]],[]],[[],[["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_2","pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_1"]]],[[],[["pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_0","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_3"]]],[[],[["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_4","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19"]]],[[],[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_0"]]],[[],[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_1"]]],[[],[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_15","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_11"]]],[[],[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_14","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_12"]]],[[],[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_13","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_13"]]],[[],[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_11","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_14"]]],[[],[["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_15","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_10"]]],[[],[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_12","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_16"]]],[[],[["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_3","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_18"]]],[[],[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_2"]]],[[],[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_3"]]],[[],[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_26","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_1"]]],[[],[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_25","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_2"]]],[[],[["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_27","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_0"]]],[[["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_2","pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_1"]],[]],[[],[["pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_1","pin-type-component_5c94b46d-7fef-4bd1-a0eb-c5c4156d6d12_0"]]],[[],[["pin-type-component_5c94b46d-7fef-4bd1-a0eb-c5c4156d6d12_1","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_2"]]],[[["pin-type-component_5c94b46d-7fef-4bd1-a0eb-c5c4156d6d12_0","pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_1"]],[]],[[["pin-type-component_5c94b46d-7fef-4bd1-a0eb-c5c4156d6d12_1","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_2"]],[]],[[],[["pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_1","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_2"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_0":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_0":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_1":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_1":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_2":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_2":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_3":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_3":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_4":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_4":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_5":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_5":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_6":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_6":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_7":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_7":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_8":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_8":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_9":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_9":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_10":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_10":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_11":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_11":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_12":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_12":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_13":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_13":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_14":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_14":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_15":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_15":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_16":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_16":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_17":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_17":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_18":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_18":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_19":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_19":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_20":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_20":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_21":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_21":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_22":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_22":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_23":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_23":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_24":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_24":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_25":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_25":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_26":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_26":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_27":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_27":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_28":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_28":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_0_29":"_","pin-type-breadboard_913a444f-47d6-41b6-8ff5-260cf7862a45_1_29":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_0_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_0_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_0_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_0_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_1_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_1_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_1_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_1_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_2_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_2_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_2_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_2_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_3_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_3_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_3_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_3_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_4_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_4_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_4_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_4_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_5_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_5_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_5_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_5_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_6_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_6_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_6_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_6_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_7_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_7_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_7_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_7_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_8_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_8_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_8_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_8_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_9_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_9_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_9_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_9_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_10_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_10_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_10_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_10_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_11_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_11_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_11_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_11_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_12_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_12_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_12_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_12_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_13_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_13_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_13_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_13_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_14_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_14_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_14_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_14_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_15_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_15_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_15_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_15_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_16_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_16_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_16_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_16_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_17_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_17_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_17_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_17_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_18_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_18_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_18_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_18_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_19_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_19_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_19_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_19_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_20_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_20_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_20_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_20_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_21_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_21_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_21_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_21_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_22_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_22_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_22_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_22_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_23_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_23_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_23_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_23_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_24_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_24_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_24_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_24_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_25_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_25_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_25_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_25_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_26_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_26_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_26_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_26_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_27_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_27_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_27_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_27_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_28_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_28_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_28_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_28_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_29_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_0_29_polarity-neg":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_29_polarity-pos":"_","pin-type-power-rail_913a444f-47d6-41b6-8ff5-260cf7862a45_1_29_polarity-neg":"_","pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_0":"0000000000000000","pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_1":"0000000000000001","pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_0":"0000000000000002","pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_1":"0000000000000003","pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_0":"0000000000000002","pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_1":"0000000000000003","pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_0":"0000000000000000","pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_1":"0000000000000001","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_0":"0000000000000000","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_1":"0000000000000001","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_2":"0000000000000004","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_3":"0000000000000005","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_4":"0000000000000006","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_5":"0000000000000002","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_6":"0000000000000003","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_7":"_","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_8":"_","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_9":"_","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_10":"_","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_11":"0000000000000007","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_12":"0000000000000008","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_13":"0000000000000009","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_14":"0000000000000010","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_15":"0000000000000011","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_16":"0000000000000012","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_0":"_","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_1":"_","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_2":"_","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_3":"_","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_4":"_","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_5":"_","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_6":"_","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_7":"_","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_8":"_","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_9":"_","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_10":"0000000000000011","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_11":"0000000000000010","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_12":"0000000000000012","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_13":"0000000000000009","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_14":"0000000000000008","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_15":"0000000000000007","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_16":"_","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_17":"_","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_18":"0000000000000005","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19":"0000000000000006","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_20":"_","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_21":"_","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_22":"_","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_23":"_","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_24":"_","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_25":"0000000000000015","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_26":"0000000000000014","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_27":"0000000000000016","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28":"0000000000000013","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_29":"_","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_30":"_","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_0":"0000000000000006","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_1":"0000000000000014","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_2":"0000000000000015","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_3":"0000000000000013","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_0":"_","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_1":"_","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_2":"_","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_3":"_","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_4":"_","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_5":"_","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_6":"_","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_7":"_","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_8":"_","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_9":"_","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_10":"_","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_11":"_","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_12":"_","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_13":"_","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_14":"_","pin-type-component_d91a83ea-e231-409e-8f49-9762e6d4f502_15":"_","pin-type-component_c4a184a4-3697-449d-9903-a666adf64026_0":"_","pin-type-component_c4a184a4-3697-449d-9903-a666adf64026_1":"_","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_0":"0000000000000016","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_1":"0000000000000006","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_2":"0000000000000013","pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_0":"0000000000000005","pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_1":"0000000000000004"},"component_id_to_pins":{"5e61949a-dd1f-4cfe-9b29-fea363a0c649":["0","1"],"34171893-90ec-4951-ae00-a62c978f62fc":["0","1"],"d7127ed3-03cf-4499-ad9a-c6fe05f81bde":["0","1"],"eb17a8e7-d287-4e59-9b8e-c4e99b281459":["0","1"],"902e1a76-96d0-4e30-b844-467374c96eb5":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16"],"59a6712b-40c1-463b-b0f1-94aaa93b70cf":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30"],"362ae36f-3285-42bd-a265-880763af6269":["0","1","2","3"],"d91a83ea-e231-409e-8f49-9762e6d4f502":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15"],"c4a184a4-3697-449d-9903-a666adf64026":["0","1"],"5db64a13-4092-4d7a-8a10-1591adc773bd":["0","1","2"],"d0a22dfe-53da-4559-b65d-0afb70497422":["0","1"]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_0","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_0","pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_0"],"0000000000000001":["pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_1","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_1","pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_1"],"0000000000000002":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_5","pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_0","pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_0"],"0000000000000003":["pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_1","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_6","pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_1"],"0000000000000005":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_3","pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_0","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_18"],"0000000000000006":["pin-type-component_362ae36f-3285-42bd-a265-880763af6269_0","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_4","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_1"],"0000000000000007":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_15","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_11"],"0000000000000008":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_14","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_12"],"0000000000000009":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_13","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_13"],"0000000000000010":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_11","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_14"],"0000000000000011":["pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_15","pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_10"],"0000000000000012":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_12","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_16"],"0000000000000013":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_2","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_3"],"0000000000000014":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_26","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_1"],"0000000000000015":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_25","pin-type-component_362ae36f-3285-42bd-a265-880763af6269_2"],"0000000000000016":["pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_27","pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_0"],"0000000000000004":["pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_1","pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_2"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000005":"Net 5","0000000000000006":"Net 6","0000000000000007":"Net 7","0000000000000008":"Net 8","0000000000000009":"Net 9","0000000000000010":"Net 10","0000000000000011":"Net 11","0000000000000012":"Net 12","0000000000000013":"Net 13","0000000000000014":"Net 14","0000000000000015":"Net 15","0000000000000016":"Net 16","0000000000000004":"Net 4"},"all_breadboard_info_list":["913a444f-47d6-41b6-8ff5-260cf7862a45_30_2_True_910_70.00000000000003_up"],"breadboard_info_list":["913a444f-47d6-41b6-8ff5-260cf7862a45_30_2_True_910_70.00000000000003_up"],"componentsData":[{"compProperties":{},"position":[-278.9124575000003,-546.5998644999999],"typeId":"aa3e6a7d-1852-40d5-bd6a-bf11ddb1f8b8","componentVersion":1,"instanceId":"5e61949a-dd1f-4cfe-9b29-fea363a0c649","orientation":"down","circleData":[[-162.5,-565.0000000000001],[-163.96533350000004,-537.067]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[418.9124575000001,-208.40013550000003],"typeId":"aa3e6a7d-1852-40d5-bd6a-bf11ddb1f8b8","componentVersion":1,"instanceId":"34171893-90ec-4951-ae00-a62c978f62fc","orientation":"up","circleData":[[302.5,-190],[303.96533349999993,-217.93300000000005]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[388.9124575000002,-553.4001355],"typeId":"aa3e6a7d-1852-40d5-bd6a-bf11ddb1f8b8","componentVersion":1,"instanceId":"d7127ed3-03cf-4499-ad9a-c6fe05f81bde","orientation":"up","circleData":[[272.5,-535],[273.96533350000004,-562.9330000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-293.9124574999997,-156.59986450000022],"typeId":"aa3e6a7d-1852-40d5-bd6a-bf11ddb1f8b8","componentVersion":1,"instanceId":"eb17a8e7-d287-4e59-9b8e-c4e99b281459","orientation":"down","circleData":[[-177.5,-175.00000000000006],[-178.9653334999996,-147.06700000000015]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"DRI0002","displayFormat":"input","showOnComp":false,"isVisibleToUser":false},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"DFRobot","displayFormat":"input","showOnComp":false,"isVisibleToUser":false}},"position":[51.54879849999996,-295.4565850000001],"typeId":"7deca677-57aa-869d-46fd-8698e7333ef9","componentVersion":1,"instanceId":"902e1a76-96d0-4e30-b844-467374c96eb5","orientation":"up","circleData":[[-72.5,-265],[-72.5,-236.96472099999997],[-22.28202950000002,-171.1770084999998],[5.7537115000000085,-171.1770084999998],[33.78944949999993,-171.1770084999998],[176.03949099999997,-242.4648279999999],[176.03949099999997,-270.5008105000001],[-0.2796650000000227,-240.40810599999986],[14.720291499999917,-240.40826649999985],[65.00821599999998,-201.51485649999984],[140.00812600000003,-201.51485649999984],[65.00832549999998,-186.5146494999999],[80.00823100000005,-186.5146494999999],[95.00822800000005,-186.5146494999999],[110.0082534999999,-186.5146494999999],[125.00814399999999,-186.5146494999999],[140.00812600000003,-186.5146494999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[166.7528155,125.60992550000023],"typeId":"518495d5-e179-49dc-aafe-d7d40a222bea","componentVersion":1,"instanceId":"59a6712b-40c1-463b-b0f1-94aaa93b70cf","orientation":"left","circleData":[[47.50000000000003,50.000000000000014],[48.339376000000044,202.79000000000008],[63.1315000000001,51.225500000000025],[77.39650000000009,50.51300000000016],[91.66300000000004,50.51300000000013],[62.48228200000008,203.65909399999998],[79.66656400000002,202.94509400000004],[93.868282,202.94509400000004],[107.07581200000001,201.45381200000014],[107.13429550000004,51.137886500000135],[122.41781800000005,50.41070450000005],[138.4285,50.41100000000003],[153.71259100000006,51.138795499999986],[168.26800000000006,49.681999999999874],[183.55179550000003,50.410091000000165],[198.83649999999997,50.409795499999944],[213.3924999999999,51.138182000000114],[228.6759999999999,51.13849999999999],[243.23199999999986,51.13759100000013],[259.24359099999987,51.13788650000018],[122.27799999999999,203.2985],[138.18490600000004,201.80750000000006],[154.09209400000006,201.3101240000001],[169.00450000000004,202.80200000000008],[184.911376,202.80200000000008],[198.8304999999999,203.29850000000005],[214.73799999999991,203.29850000000005],[229.41249999999988,203.29850000000005],[244.8225939999999,203.29909400000014],[261.2272179999998,203.29878200000013],[307.60749999999945,126.89900000000014]],"code":"496,folder,{\"name\":\"sketch\",\"id\":\"227e2f43-4ab3-4da3-9ba0-ccc4512a3a7a\",\"explorerHtmlId\":\"2891ad08-2dbb-4e4f-9439-0c08f504d9a9\",\"nameHtmlId\":\"2b296b16-9ce7-4a06-bd0b-9c72c6f4cb5f\",\"nameInputHtmlId\":\"d2a72738-34a3-47fa-a99b-55fa2c4931b0\",\"explorerChildHtmlId\":\"d17dc3a5-e9f4-4771-b8cd-a2c25443db84\",\"explorerCarrotOpenHtmlId\":\"56ff546a-a8db-48ff-8799-613c7fe8cd12\",\"explorerCarrotClosedHtmlId\":\"77c85943-1122-4f6b-a18f-8f45d99a0917\",\"arduinoBoardFqbn\":\"\",\"arduinoBoardName\":\"\",\"arduinoPortAddress\":\"\"},2,16964,file,{\"name\":\"sketch.ino\",\"id\":\"1c723573-fe01-4b50-8611-0c22be2c8ef9\",\"explorerHtmlId\":\"eb8f6fcc-4cb4-4876-a50a-d47701e5c42c\",\"nameHtmlId\":\"be697b69-9b50-474c-8e0c-26145ab74931\",\"nameInputHtmlId\":\"a3cf0ed3-2636-47dc-90dd-a634532bf636\",\"code\":\"#include <Robojax_L298N_DC_motor.h> \\n#include <BluetoothSerial.h> \\n#include <ESP32Servo.h> \\n//---------Flag structure-----------------------------------------\\ntypedef  struct  _vFlag\\n{\\n  uint8_t BTFlag =  0 ;\\n  uint8_t L298NFlag =  0 ;\\n  uint8_t HCSR04Flag = 1 ; \\n  uint8_t LEDFlag =  1 ;\\n  uint8_t ServoFlag =  0 ;\\n  uint8_t initial_Flag =  0 ;\\n  uint8_t FunctionFlag =  0 ;\\n  uint8_t back_light_Flag =  0 ;\\n  uint8_t front_light_Flag =  0 ;\\n} vFlag ;\\nvFlag * flag_Ptr;\\nvFlag flag;\\n//---------BT------------------------\\nBluetoothSerial SerialBT;\\n//------------------servo---------------------------------\\nServo myservo;   // create servo object to control a servo\\n// Recommended PWM GPIO pins on the ESP32 include 2,4,12-19,21-23,25-27,32-33\\n#define servoPin 13\\n//------LED------------------\\n#define LED_BUILTIN 2\\n//-------------L298--------------------------------------------------\\n// motor 1 settings\\n#define CHA 0\\n#define ENA 4 // this pin must be PWM enabled pin if Arduino board is used\\n#define IN1 16\\n#define IN2 17\\n// motor 2 settings\\n#define IN3 18\\n#define IN4 19\\n#define ENB 5 // this pin must be PWM enabled pin if Arduino board is used\\n#define CHB 1\\n\\nconst  int CCW =  2 ; // do not change\\nconst  int CW   =  1 ; // do not change\\n\\n#define motor1 1 // do not change\\n#define motor2 2 // do not change\\n\\n// for two motors without debug information // Watch video instruciton for this line: https://youtu.be/2JTMqURJTwg\\nRobojax_L298N_DC_motor  motors ( IN1 , IN2 , ENA , CHA ,   IN3 , IN4 , ENB , CHB );\\n//------Bluetooth RC Controller Define ----\\n#define back_light 21\\n#define front_light 22\\n//-----hcsr04 sensor------------------\\n#define TRIGPIN_PIN 12\\n#define ECHO_PIN 14 \\nlong duration;\\nunsigned  long currentMillis =  0 ;\\n//----------global ---------------------\\n#define MAX_DISTANCE 200\\n#define MAX_SPEED 190 // Sets speed of DC motors\\nint speedSet =  0 ;\\nint distance =  60 ;\\nint distanceR =  0 ;\\nint distanceL =  0 ;\\n//--------- uart structure -----------------------------------------------\\n//----------uart--------------\\n#define LINE_BUFFER_LENGTH 64\\ntypedef  struct  _vUart\\n{\\n  char c;\\n  int lineIndex =  0 ;\\n  int line1Index =  0 ;\\n  int BTlineIndex =  0 ;\\n  bool lineIsComment;\\n  bool lineSemiColon;\\n  //char *line;\\n  char  line [ 128 ];\\n  //char line1[128];\\n  char  BTline [ 20 ];\\n  //char R_line[20];\\n  //char L_line[20];\\n  String inputString;\\n  String BTinputString;\\n  String S1inputString;\\n  int  V [ 16 ];\\n  char  ctemp [ 30 ];\\n  char  I2C_Data [ 80 ];\\n  int DC_Spped =  50 ;\\n  float  Voltage [ 16 ];\\n  int  Buffer [ 128 ];\\n  int StartCnt =  0 ;\\n  int ReadCnt =  0 ;\\n  int sensorValue =  0 ;\\n} vUart ;\\nvUart * Uart_Ptr;\\nvUart Uart;\\n//-------------------------------------\\nTaskHandle_t huart;\\nTaskHandle_t hfunction;\\n\\nvoid  vUARTTask ( void  * pvParameters );\\nvoid  vFunctionTask ( void  * pvParameters );\\n//------------------------------------------------------------------------------\\nvoid  initial ()\\n{\\n  Serial . println ( F ( \\\"Create Task\\\" ));\\n  //----------------------------------------------------------------------\\n  xTaskCreatePinnedToCore (\\n    vUARTTask, \\\"UARTTask\\\" // A name just for humans\\n    ,\\n    1024 // This stack size can be checked & adjusted by reading the Stack Highwater\\n    ,\\n    NULL , 3 // Priority, with 3 (configMAX_PRIORITIES - 1) being the highest, and 0 being the lowest.\\n    ,\\n    & huart //handle\\n    ,\\n    0 );\\n\\n  xTaskCreatePinnedToCore (\\n    vFunctionTask, \\\"FunctionTask\\\"\\n    ,\\n    1024 // Stack size\\n    ,\\n    NULL , 1 // Priority\\n    ,\\n    & hfunction\\n    ,\\n    1 );\\n\\n  //----------------------------------------------------------------------\\n\\n  //----------------------------------------------------------------------\\n}\\n\\nvoid  Forward ()\\n{  \\n  //motors.rotate(motor1, 60, CCW);\\n  //motors.rotate(motor2, 60, CCW);\\n  digitalWrite (IN1, LOW);\\n  digitalWrite (IN2, HIGH);\\n  analogWrite (ENA, 100 );\\n  digitalWrite (IN3, LOW);\\n  digitalWrite (IN4, HIGH);\\n  analogWrite (ENB, 100 );\\n}\\n\\nvoid  Reverse () {\\n  //motors.rotate(motor2, 70, CW);\\n  //motors.rotate(motor1, 70, CW);\\n  digitalWrite (IN1, HIGH);\\n  digitalWrite (IN2, LOW);\\n  analogWrite (ENA, 100 );\\n  digitalWrite (IN3, HIGH);\\n  digitalWrite (IN4, LOW);\\n  analogWrite (ENB, 100 );\\n}\\nvoid  Left ()\\n{\\n  //motors.rotate(motor1, 70, CW);\\n  //motors.rotate(motor2, 70, CCW); //LF\\n  digitalWrite (IN1, LOW);\\n  digitalWrite (IN2, HIGH);\\n  analogWrite (ENA, 100 );\\n}\\nvoid  Right ()\\n{\\n  digitalWrite (IN3, LOW);\\n  digitalWrite (IN4, HIGH);\\n  analogWrite (ENB, 100 );\\n  //motors.rotate(motor1, 70, CCW); //RF\\n  //motors.rotate(motor2, 70, CW);\\n}\\nvoid  Stop ()\\n{\\n  motors . brake ( 1 );\\n  motors . brake ( 2 );\\n  //myservo.detach();\\n}\\n//-------------------------------------------------\\nvoid  setup ()\\n{\\n  Serial.begin ( 9600 ) ;​\\n  Serial . println ( F ( \\\"init\\\" ));\\n  initial ();\\n  SerialBT .begin ( \\\"BT_L298N\\\" ) ;\\n  myservo.setPeriodHertz ( 50 )     ;​\\n  myservo . attach (servoPin, 500 , 2400 );\\n  pinMode (LED_BUILTIN, OUTPUT);\\n  pinMode (TRIGPIN_PIN, OUTPUT);\\n  pinMode (ECHO_PIN, INPUT);\\n  pinMode (IN1, OUTPUT);\\n  pinMode (IN2, OUTPUT);\\n  pinMode (IN3, OUTPUT);\\n  pinMode (IN4, OUTPUT);\\n  pinMode (ENA, OUTPUT);\\n  pinMode (ENB, OUTPUT);\\n  pinMode (back_light, OUTPUT);\\n  pinMode (front_light, OUTPUT);\\n  motors.begin ( ) ;\\n  myservo . write ( 90 );\\n}\\n//-----------------------------------------\\nvoid  loop ()\\n{\\n  Serial .print ( F ( \\\"Main at core:\\\" ) );\\n  Serial .println ( xPortGetCoreID ()) ;\\n  while ( 1 )\\n  {\\n    if ( flag . HCSR04Flag == 1 )\\n    {\\n      if (distance <= 35 )\\n      {\\n        Stop ();\\n        delay ( 200 );\\n        Reverse ();\\n        delay ( 400 );\\n        Stop ();\\n        delay ( 100 );\\n        flag . HCSR04Flag = 2 ;\\n        delay ( 2000 );\\n        flag . HCSR04Flag = 3 ;\\n        delay ( 2000 );\\n        flag . HCSR04Flag = 1 ;\\n        if ((distanceR >= distanceL) )\\n        {\\n          Left ();\\n          delay ( 700 );\\n          Stop ();\\n          delay ( 200 );\\n          flag . HCSR04Flag = 1 ;\\n        }\\n        else \\n        {\\n          Right ();\\n          delay ( 700 );\\n          Stop ();\\n          delay ( 200 );\\n          flag . HCSR04Flag = 1 ;\\n        }\\n        myservo . write ( 90 );\\n        delay ( 1000 );\\n      }\\n      else \\n      {\\n        flag . HCSR04Flag = 1 ;\\n        Forward ();\\n        delay ( 100 );\\n        Stop ();\\n        delay ( 30 );\\n      }      \\n    }\\n    vTaskDelay ( 1 );\\n  }\\n}\\n//----------------------------------------\\nvoid  processCommand ( char  * data )\\n{\\n  int len, xlen, ylen, zlen, alen;\\n  int tempDIO;\\n  String stemp;\\n\\n  len =  Uart . inputString . length ();\\n  //---------------------------------------\\n  if ( strstr (data, \\\"VER\\\" ) !=  NULL )\\n  {\\n    Serial . println ( F ( \\\"ESP32_20230710\\\" ));\\n  }\\n  //-------------- HCSR04 --------------------\\n  if ( strstr (data, \\\"HCSR04_ON\\\" ) !=  NULL )\\n  {\\n    flag . HCSR04Flag  =  1 ;\\n    Serial . println ( F ( \\\"HCSR04_ON\\\" ));\\n  }\\n  if ( strstr (data, \\\"HCSR04_OFF\\\" ) !=  NULL )\\n  {\\n    flag . HCSR04Flag  =  0 ;\\n    Serial . println ( F ( \\\"HCSR04_OFF\\\" ));\\n  }  \\n  //----------------L298N----------\\n  if ( strstr (data, \\\"F\\\" ) !=  NULL )\\n  {\\n    Serial .println ( F ( \\\"Forward\\\" )) ;\\n    Forward ();\\n    //forward();\\n    \\n  }\\n  if ( strstr (data, \\\"L\\\" ) !=  NULL )\\n  {\\n    Serial .println ( F ( \\\"Left\\\" ) );\\n    Left ();\\n  }\\n  if ( strstr (data, \\\"R\\\" ) !=  NULL )\\n  {\\n    Serial .println ( F ( \\\"Right\\\" )) ;\\n    Right ();\\n  }\\n  if ( strstr (data, \\\"B\\\" ) !=  NULL )\\n  {\\n    Serial . println ( F ( \\\"Reverse\\\" ));\\n    Reverse ();\\n    //backward();\\n  }\\n  if ( strstr (data, \\\"S\\\" ) !=  NULL )\\n  {\\n    Serial .println ( F ( \\\"Stop\\\" ) );\\n    Stop ();\\n  }\\n  //-----------------servo---------\\n  //-------------- Servo --------------------\\n  if ( strstr (data, \\\"SERVO_5\\\" ) !=  NULL )\\n  {\\n    Serial . println ( F ( \\\"SERVO_5\\\" ));\\n    myservo . write ( 5 );\\n    //myservo.detach();\\n  }\\n  if ( strstr (data, \\\"SERVO_10\\\" ) !=  NULL )\\n  {\\n    Serial . println ( F ( \\\"SERVO_10\\\" ));\\n    myservo . write ( 10 );\\n  }\\n  if ( strstr (data, \\\"SERVO_20\\\" ) !=  NULL )\\n  {\\n    Serial . println ( F ( \\\"SERVO_20\\\" ));\\n    myservo . write ( 20 );\\n  }\\n  if ( strstr (data, \\\"SERVO_30\\\" ) !=  NULL )\\n  {\\n    Serial . println ( F ( \\\"SERVO_30\\\" ));\\n    myservo . write ( 30 );\\n  }\\n  if ( strstr (data, \\\"SERVO_50\\\" ) !=  NULL )\\n  {\\n    Serial . println ( F ( \\\"SERVO_50\\\" ));\\n    myservo . write ( 50 );\\n  }\\n  if ( strstr (data, \\\"SERVO_80\\\" ) !=  NULL )\\n  {\\n    Serial . println ( F ( \\\"SERVO_80\\\" ));\\n    myservo . write ( 80 );\\n  }\\n  if ( strstr (data, \\\"SERVO_90\\\" ) !=  NULL )\\n  {\\n    Serial . println ( F ( \\\"SERVO_90\\\" ));\\n    myservo . write ( 90 );\\n  }\\n  if ( strstr (data, \\\"SERVO_100\\\" ) !=  NULL )\\n  {\\n    Serial . println ( F ( \\\"SERVO_100\\\" ));\\n    myservo . write ( 100 );\\n  }\\n  if ( strstr (data, \\\"SERVO_120\\\" ) !=  NULL )\\n  {\\n    Serial . println ( F ( \\\"SERVO_120\\\" ));\\n    myservo . write ( 120 );\\n  }\\n  if ( strstr (data, \\\"SERVO_140\\\" ) !=  NULL )\\n  {\\n    Serial . println ( F ( \\\"SERVO_140\\\" ));\\n    myservo . write ( 140 );\\n  }\\n  if ( strstr (data, \\\"SERVO_150\\\" ) !=  NULL )\\n  {\\n    Serial . println ( F ( \\\"SERVO_150\\\" ));\\n    myservo . write ( 150 );\\n  }\\n}\\n//-----------------------------------------\\n//------------------BT-----------------\\nvoid  BTprocessCommand ( String  data )\\n{\\n  if (data == \\\"FS\\\" )\\n  {\\n    Serial .println ( F ( \\\"Forward\\\" )) ;\\n    Forward ();\\n  }\\n  if (data ==  \\\"LS\\\" )\\n  {\\n    Serial .println ( F ( \\\"Left\\\" ) );\\n    Left ();\\n  }\\n  if (data ==  \\\"RS\\\" )\\n  {\\n    Serial .println ( F ( \\\"Right\\\" )) ;\\n    Right ();\\n  }\\n  if (data ==  \\\"BS\\\" )\\n  {\\n    Serial . println ( F ( \\\"Reverse\\\" ));\\n    Reverse ();\\n  }\\n  if (data ==  \\\"S\\\" )\\n  {\\n    Serial .println ( F ( \\\"Stop\\\" ) );\\n    Stop ();\\n  }\\n  if (data ==  \\\"X\\\" )\\n  {\\n    flag . HCSR04Flag = 0 ;\\n    Serial .println ( F ( \\\"Stop\\\" ) );\\n    Stop ();\\n    flag . back_light_Flag = 2 ;\\n    flag . HCSR04Flag = 0 ;\\n  }\\n  if (data ==  \\\"x\\\" )\\n  {\\n    Serial .println ( F ( \\\"Stop\\\" ) );\\n    Stop ();\\n    flag . back_light_Flag = 0 ;\\n    flag . HCSR04Flag = 1 ;\\n  }\\n  if (data ==  \\\"FGFS\\\" )\\n  {\\n    //LF\\n    motors . rotate (motor1, 60 , CCW);\\n    motors . rotate (motor2, 100 , CCW);\\n  }\\n  if (data ==  \\\"FIFS\\\" )\\n  {\\n    //RF\\n    motors . rotate (motor1, 100 , CCW);\\n    motors . rotate (motor2, 60 , CCW);\\n  }\\n  if (data ==  \\\"BHBS\\\" )\\n  {\\n    //LB\\n    motors . rotate (motor1, 60 , CW);\\n    motors . rotate (motor2, 100 , CW);\\n  }\\n  if (data ==  \\\"BJBS\\\" )\\n  {\\n    //RB\\n    motors . rotate (motor1, 100 , CW);\\n    motors . rotate (motor2, 60 , CW);\\n  }\\n  if (data ==  \\\"U\\\" )\\n  {\\n    //backlight\\n    digitalWrite (back_light, HIGH);  \\n    flag . back_light_Flag = 1 ;\\n    //Serial.println(F(\\\"light\\\"));\\n  }\\n  if (data ==  \\\"u\\\" )\\n  {\\n    //backlight\\n    digitalWrite (back_light, LOW);\\n    flag . back_light_Flag = 0 ;\\n    //Serial.println(F(\\\"lightoff\\\"));\\n  }\\n  if (data ==  \\\"W\\\" )\\n  {\\n    digitalWrite (front_light, HIGH);  \\n    flag . front_light_Flag = 1 ;\\n    //Serial.println(F(\\\"light\\\"));\\n  }\\n  if (data ==  \\\"w\\\" )\\n  {\\n    digitalWrite (front_light, LOW);\\n    flag . front_light_Flag = 0 ;\\n    //Serial.println(F(\\\"lightoff\\\"));\\n  }\\n}\\n//-------------------------------------------\\nvoid  vUARTTask ( void  * pvParameters )\\n{\\n  ( void )pvParameters;\\n\\n  Serial . print ( F ( \\\"UARTTask at core:\\\" ));\\n  Serial .println ( xPortGetCoreID ()) ;\\n  for (;;)\\n  {\\n    while ( Serial . available () >  0 )\\n    {\\n      Uart.c = Serial.read ( ) ;​​  \\n  \\n      if (( Uart . c  ==  ' \\\\n ' ) || ( Uart . c  ==  ' \\\\r ' ))\\n      { // End of line reached\\n        if ( Uart . lineIndex  >  0 )\\n        { // Line is complete. Then execute!\\n          Uart . line [ Uart . lineIndex ] =  ' \\\\0 ' ; // Terminate string\\n          //Serial.println( F(\\\"Debug\\\") );\\n          //Serial.println( Uart.inputString );\\n          processCommand ( Uart . line );\\n          Uart . lineIndex  =  0 ;\\n          Uart . inputString  =  \\\"\\\" ;\\n        }\\n        else\\n        {\\n          // Empty or comment line. Skip block.\\n        }\\n        Uart.lineIsComment = false ;​​  \\n        Uart.lineSemiColon = false ;​​  \\n        Serial . println ( F ( \\\"ok>\\\" ));\\n      }\\n      else\\n      {\\n        //Serial.println( c );\\n        if (( Uart . lineIsComment ) || ( Uart . lineSemiColon ))\\n        {\\n          if ( Uart . c  ==  ')' )\\n            Uart . lineIsComment  =  false ; // End of comment. Resume line.\\n        }\\n        else\\n        {\\n          if ( Uart . c  ==  '/' )\\n          { // Block delete not supported. Ignore character.\\n          }\\n          else  if ( Uart . c  ==  '~' )\\n          { // Enable comments flag and ignore all characters until ')' or EOL.\\n            Uart . lineIsComment  =  true ;\\n          }\\n          else  if ( Uart . c  ==  ';' )\\n          {\\n            Uart . lineSemiColon  =  true ;\\n          }\\n          else  if ( Uart . lineIndex  >= LINE_BUFFER_LENGTH -  1 )\\n          {\\n            Serial . println ( \\\"ERROR - lineBuffer overflow\\\" );\\n            Uart.lineIsComment = false ;​​  \\n            Uart.lineSemiColon = false ;​​  \\n          }\\n          else  if ( Uart . c  >=  'a'  &&  Uart . c  <=  'z' )\\n          { // Upcase lowercase\\n            Uart . line [ Uart . lineIndex ] =  Uart . c  -  'a'  +  'A' ;\\n            Uart . lineIndex  =  Uart . lineIndex  +  1 ;\\n            Uart . inputString  += ( char )( Uart . c  -  'a'  +  'A' );\\n          }\\n          else\\n          {\\n            Uart . line [ Uart . lineIndex ] =  Uart . c ;\\n            Uart . lineIndex  =  Uart . lineIndex  +  1 ;\\n            Uart . inputString  +=  Uart . c ;\\n          }\\n        }\\n      }\\n    } //while (Serial.available() > 0)\\n    while ( SerialBT . available ())\\n    {\\n      flag . L298NFlag = 1 ;\\n      String BTdata =  SerialBT . readString ();\\n      Stop ();\\n      Serial.println (BTdata ) ;\\n      BTprocessCommand (BTdata); // do something with the command\\n    } //while (BT.available())\\n    vTaskDelay ( 1 );\\n  }\\n}\\nvoid  vFunctionTask ( void  * pvParameters )\\n{\\n  ( void )pvParameters;\\n\\n  Serial . print ( F ( \\\"FunctionTask at core:\\\" ));\\n  Serial .println ( xPortGetCoreID ()) ;\\n  for (;;) // A Task shall never return or exit.\\n  {\\n    if ( flag . HCSR04Flag == 1 )\\n    {\\n      currentMillis =  millis ();\\n      myservo . write ( 90 );\\n      digitalWrite (TRIGPIN_PIN, LOW);  \\n      delayMicroseconds ( 2 );  \\n      digitalWrite (TRIGPIN_PIN, HIGH);\\n      delayMicroseconds ( 10 );\\n      digitalWrite (TRIGPIN_PIN, LOW);  \\n      duration =  pulseIn (ECHO_PIN, HIGH);\\n      distance = duration / 29 / 2 ;\\n      if (duration == 0 )\\n      {\\n        Serial .println ( \\\" No pulse is from sensor\\\" );\\n      }\\n      else \\n      {\\n        Serial .print ( \\\"Ultrasonic sensor is shown distance:\\\" );\\n        Serial . print ( distance );\\n        Serial . println ( \\\"cm\\\" );\\n        Serial .print (distanceR - distanceL) ;\\n        Serial . println ( \\\"cm\\\" );\\n      }\\n    }\\n    if ( flag . HCSR04Flag == 2 )   //lookRight\\n    {\\n      myservo . write ( 20 );\\n      digitalWrite (TRIGPIN_PIN, LOW);  \\n      delayMicroseconds ( 2 );  \\n      digitalWrite (TRIGPIN_PIN, HIGH);\\n      delayMicroseconds ( 10 );  \\n      digitalWrite (TRIGPIN_PIN, LOW);  \\n      duration =  pulseIn (ECHO_PIN, HIGH);\\n      distanceR = duration / 29 / 2 ;\\n      if (duration == 0 )\\n      {\\n        Serial .println ( \\\" No pulse is from sensor\\\" );\\n      }\\n      else \\n      {\\n        //Serial.print(\\\"Ultrasonic sensor is shown distanceR:\\\");\\n        //Serial.print(distanceR);\\n        //Serial.println(\\\"cm\\\");\\n      }\\n    }\\n    if ( flag . HCSR04Flag == 3 )   //lookLeft\\n    {\\n      myservo . write ( 160 );\\n      digitalWrite (TRIGPIN_PIN, LOW);  \\n      delayMicroseconds ( 2 );  \\n      digitalWrite (TRIGPIN_PIN, HIGH);\\n      delayMicroseconds ( 10 );  \\n      digitalWrite (TRIGPIN_PIN, LOW);  \\n      duration =  pulseIn (ECHO_PIN, HIGH);\\n      distanceL = duration / 29 / 2 ;\\n      if (duration == 0 )\\n      {\\n        Serial .println ( \\\" No pulse is from sensor\\\" );\\n      }\\n      else \\n      {\\n        //Serial.print(\\\"Ultrasonic sensor is shown distanceL:\\\");\\n        //Serial.print(distanceL);\\n        //Serial.println(\\\"cm\\\");\\n      }\\n    }\\n    vTaskDelay ( 1 );\\n  }\\n}\\n\\n\\n\"},0,252,file,{\"name\":\"documentation.txt\",\"id\":\"976f74aa-852e-4922-ac9f-2ffeeda25571\",\"explorerHtmlId\":\"e6cefdc9-8f70-4d36-a023-8fec4ebddba2\",\"nameHtmlId\":\"fcaaf6fc-647c-40db-8e7b-3d809a4abbde\",\"nameInputHtmlId\":\"89afa26c-60de-43c2-b8f2-93269e4cae2e\",\"code\":\"\"},0,","codeLabelPosition":[166.75281549999994,41.34585050000021],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"SEN-15569","displayFormat":"input","showOnComp":false,"isVisibleToUser":false},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"SparkFun","displayFormat":"input","showOnComp":false,"isVisibleToUser":false}},"position":[522.0136135,13.496435000000133],"typeId":"f7a95729-a811-496b-83f5-7789de376adf","componentVersion":2,"instanceId":"362ae36f-3285-42bd-a265-880763af6269","orientation":"up","circleData":[[497.5,79.99999999999997],[512.4992245000001,79.99999999999997],[527.4999985000002,79.99530950000005],[542.4984445,79.99374950000012]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[974.3166684999998,-246.74021950000002],"typeId":"3b4a66b1-0d1b-40c2-92f7-ec286f5c89ab","componentVersion":2,"instanceId":"d91a83ea-e231-409e-8f49-9762e6d4f502","orientation":"up","circleData":[[887.5000000000001,-370.00000000000006],[885.7465000000003,-349.4826235000001],[887.5000000000001,-326.90602900000005],[888.6390625,-307.2204955],[886.0537195000003,-289.2899620000001],[886.3609390000003,-266.4046480000001],[887.8072195000001,-247.33505350000013],[887.8072195000001,-225.89602000000014],[1073.2501705000004,-371.7535000000001],[1073.5573885000003,-350.92890400000005],[1073.8646080000003,-329.79859000000005],[1073.8646080000003,-308.97399550000006],[1073.5573885000003,-290.7362440000001],[1073.5573885000003,-269.6044300000001],[1073.5573885000003,-247.02783400000015],[1072.1111080000005,-229.40302000000014]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1260.6234745000002,-617.8651329999999],"typeId":"d749d278-6a0d-4deb-825c-1b35ffc56ae5","componentVersion":1,"instanceId":"c4a184a4-3697-449d-9903-a666adf64026","orientation":"up","circleData":[[1247.5,-700.0000000000001],[1226.3215,-700.0000000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[85.0307214999997,332.2454],"typeId":"437e01f5-4fa2-4201-ac70-cfe748b41bde","componentVersion":1,"instanceId":"5db64a13-4092-4d7a-8a10-1591adc773bd","orientation":"up","circleData":[[182.5,365],[176.77668700000004,381.1663985000001],[173.06546049999997,394.8784985000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1321","displayFormat":"input","showOnComp":false,"isVisibleToUser":false},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Adafruit Industries","displayFormat":"input","showOnComp":false,"isVisibleToUser":false}},"position":[-427.4864915000003,231.41439200000005],"typeId":"7dbe2b3d-2053-a5aa-7735-837175ae747c","componentVersion":1,"instanceId":"d0a22dfe-53da-4559-b65d-0afb70497422","orientation":"up","circleData":[[-327.5,110],[-327.5,95.00210750000006]],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-714.00000","left":"-536.72507","width":"1917.70752","height":"1236.50000","x":"-536.72507","y":"-714.00000"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_0\",\"endPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_0\",\"rawStartPinId\":\"pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_0\",\"rawEndPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-162.5000000000_-565.0000000000\\\",\\\"-117.5000000000_-565.0000000000\\\",\\\"-117.5000000000_-265.0000000000\\\",\\\"-72.5000000000_-265.0000000000\\\"]}\"}","{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_0\",\"endPinId\":\"pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_0\",\"rawStartPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_0\",\"rawEndPinId\":\"pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-72.5000000000_-265.0000000000\\\",\\\"-125.0000000000_-265.0000000000\\\",\\\"-125.0000000000_-175.0000000000\\\",\\\"-177.5000000000_-175.0000000000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_1\",\"endPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_1\",\"rawStartPinId\":\"pin-type-component_5e61949a-dd1f-4cfe-9b29-fea363a0c649_1\",\"rawEndPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-163.9653335000_-537.0670000000\\\",\\\"-118.2326667500_-537.0670000000\\\",\\\"-118.2326667500_-236.9647210000\\\",\\\"-72.5000000000_-236.9647210000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_1\",\"endPinId\":\"pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_1\",\"rawStartPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_1\",\"rawEndPinId\":\"pin-type-component_eb17a8e7-d287-4e59-9b8e-c4e99b281459_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-72.5000000000_-236.9647210000\\\",\\\"-125.7326667500_-236.9647210000\\\",\\\"-125.7326667500_-147.0670000000\\\",\\\"-178.9653335000_-147.0670000000\\\"]}\"}","{\"color\":\"#0E4CA1\",\"startPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_5\",\"endPinId\":\"pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_0\",\"rawStartPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_5\",\"rawEndPinId\":\"pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"176.0394910000_-242.4648280000\\\",\\\"224.2697455000_-242.4648280000\\\",\\\"224.2697455000_-535.0000000000\\\",\\\"272.5000000000_-535.0000000000\\\"]}\"}","{\"color\":\"#0E4CA1\",\"startPinId\":\"pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_0\",\"endPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_5\",\"rawStartPinId\":\"pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_0\",\"rawEndPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"302.5000000000_-190.0000000000\\\",\\\"212.5000000000_-190.0000000000\\\",\\\"212.5000000000_-242.4648280000\\\",\\\"176.0394910000_-242.4648280000\\\"]}\"}","{\"color\":\"#FFE502\",\"startPinId\":\"pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_1\",\"endPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_6\",\"rawStartPinId\":\"pin-type-component_34171893-90ec-4951-ae00-a62c978f62fc_1\",\"rawEndPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"303.9653335000_-217.9330000000\\\",\\\"212.5000000000_-217.9330000000\\\",\\\"212.5000000000_-270.5008105000\\\",\\\"176.0394910000_-270.5008105000\\\"]}\"}","{\"color\":\"#FFE502\",\"startPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_6\",\"endPinId\":\"pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_1\",\"rawStartPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_6\",\"rawEndPinId\":\"pin-type-component_d7127ed3-03cf-4499-ad9a-c6fe05f81bde_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"176.0394910000_-270.5008105000\\\",\\\"225.0024122500_-270.5008105000\\\",\\\"225.0024122500_-562.9330000000\\\",\\\"273.9653335000_-562.9330000000\\\"]}\"}","{\"color\":\"#FF74A3\",\"startPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_3\",\"endPinId\":\"pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_0\",\"rawStartPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_3\",\"rawEndPinId\":\"pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"5.7537115000_-171.1770085000\\\",\\\"5.7537115000_-10.0000000000\\\",\\\"-282.5000000000_-10.0000000000\\\",\\\"-282.5000000000_110.0000000000\\\",\\\"-327.5000000000_110.0000000000\\\"]}\"}","{\"color\":\"#FF74A3\",\"startPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_18\",\"endPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_3\",\"rawStartPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_18\",\"rawEndPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"243.2320000000_51.1375910000\\\",\\\"243.2320000000_-70.0000000000\\\",\\\"5.7537115000_-70.0000000000\\\",\\\"5.7537115000_-171.1770085000\\\"]}\"}","{\"color\":\"#968AE8\",\"startPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19\",\"endPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_4\",\"rawStartPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19\",\"rawEndPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"259.2435910000_51.1378865000\\\",\\\"259.2435910000_-70.0000000000\\\",\\\"33.7894495000_-70.0000000000\\\",\\\"33.7894495000_-171.1770085000\\\"]}\"}","{\"color\":\"#968AE8\",\"startPinId\":\"pin-type-component_362ae36f-3285-42bd-a265-880763af6269_0\",\"endPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19\",\"rawStartPinId\":\"pin-type-component_362ae36f-3285-42bd-a265-880763af6269_0\",\"rawEndPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"497.5000000000_80.0000000000\\\",\\\"497.5000000000_95.0000000000\\\",\\\"362.5000000000_95.0000000000\\\",\\\"362.5000000000_20.0000000000\\\",\\\"259.2435910000_20.0000000000\\\",\\\"259.2435910000_51.1378865000\\\"]}\"}","{\"color\":\"#968AE8\",\"startPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19\",\"endPinId\":\"pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_1\",\"rawStartPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_19\",\"rawEndPinId\":\"pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"259.2435910000_51.1378865000\\\",\\\"259.2435910000_20.0000000000\\\",\\\"347.5000000000_20.0000000000\\\",\\\"347.5000000000_381.1663985000\\\",\\\"176.7766870000_381.1663985000\\\"]}\"}","{\"color\":\"#98FF52\",\"startPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_15\",\"endPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_11\",\"rawStartPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_15\",\"rawEndPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_11\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"198.8365000000_50.4097955000\\\",\\\"198.8365000000_-70.0000000000\\\",\\\"65.0083255000_-70.0000000000\\\",\\\"65.0083255000_-186.5146495000\\\"]}\"}","{\"color\":\"#A75740\",\"startPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_14\",\"endPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_12\",\"rawStartPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_14\",\"rawEndPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_12\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"183.5517955000_50.4100910000\\\",\\\"183.5517955000_-70.0000000000\\\",\\\"80.0082310000_-70.0000000000\\\",\\\"80.0082310000_-186.5146495000\\\"]}\"}","{\"color\":\"#01FFFE\",\"startPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_13\",\"endPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_13\",\"rawStartPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_13\",\"rawEndPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_13\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"168.2680000000_49.6820000000\\\",\\\"168.2680000000_-70.0000000000\\\",\\\"95.0082280000_-70.0000000000\\\",\\\"95.0082280000_-186.5146495000\\\"]}\"}","{\"color\":\"#FE8900\",\"startPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_11\",\"endPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_14\",\"rawStartPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_11\",\"rawEndPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_14\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"138.4285000000_50.4110000000\\\",\\\"138.4285000000_-70.0000000000\\\",\\\"110.0082535000_-70.0000000000\\\",\\\"110.0082535000_-186.5146495000\\\"]}\"}","{\"color\":\"#BDC6FF\",\"startPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_10\",\"endPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_15\",\"rawStartPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_10\",\"rawEndPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_15\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"122.4178180000_50.4107045000\\\",\\\"122.4178180000_-70.0000000000\\\",\\\"125.0081440000_-70.0000000000\\\",\\\"125.0081440000_-186.5146495000\\\"]}\"}","{\"color\":\"#BB8800\",\"startPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_12\",\"endPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_16\",\"rawStartPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_12\",\"rawEndPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_16\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"153.7125910000_51.1387955000\\\",\\\"153.7125910000_-70.0000000000\\\",\\\"140.0081260000_-70.0000000000\\\",\\\"140.0081260000_-186.5146495000\\\"]}\"}","{\"color\":\"#7544B1\",\"startPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28\",\"endPinId\":\"pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_2\",\"rawStartPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28\",\"rawEndPinId\":\"pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"244.8225940000_203.2990940000\\\",\\\"244.8225940000_394.8784985000\\\",\\\"173.0654605000_394.8784985000\\\"]}\"}","{\"color\":\"#7544B1\",\"startPinId\":\"pin-type-component_362ae36f-3285-42bd-a265-880763af6269_3\",\"endPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28\",\"rawStartPinId\":\"pin-type-component_362ae36f-3285-42bd-a265-880763af6269_3\",\"rawEndPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_28\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"542.4984445000_79.9937495000\\\",\\\"542.4984445000_230.0000000000\\\",\\\"244.8225940000_230.0000000000\\\",\\\"244.8225940000_203.2990940000\\\"]}\"}","{\"color\":\"#A5FFD2\",\"startPinId\":\"pin-type-component_362ae36f-3285-42bd-a265-880763af6269_1\",\"endPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_26\",\"rawStartPinId\":\"pin-type-component_362ae36f-3285-42bd-a265-880763af6269_1\",\"rawEndPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_26\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"512.4992245000_80.0000000000\\\",\\\"512.4992245000_230.0000000000\\\",\\\"214.7380000000_230.0000000000\\\",\\\"214.7380000000_203.2985000000\\\"]}\"}","{\"color\":\"#FFA6FE\",\"startPinId\":\"pin-type-component_362ae36f-3285-42bd-a265-880763af6269_2\",\"endPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_25\",\"rawStartPinId\":\"pin-type-component_362ae36f-3285-42bd-a265-880763af6269_2\",\"rawEndPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_25\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"527.4999985000_79.9953095000\\\",\\\"527.4999985000_230.0000000000\\\",\\\"198.8305000000_230.0000000000\\\",\\\"198.8305000000_203.2985000000\\\"]}\"}","{\"color\":\"#774D00\",\"startPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_27\",\"endPinId\":\"pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_0\",\"rawStartPinId\":\"pin-type-component_59a6712b-40c1-463b-b0f1-94aaa93b70cf_27\",\"rawEndPinId\":\"pin-type-component_5db64a13-4092-4d7a-8a10-1591adc773bd_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"229.4125000000_203.2985000000\\\",\\\"229.4125000000_365.0000000000\\\",\\\"182.5000000000_365.0000000000\\\"]}\"}","{\"color\":\"#B500FF\",\"startPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_2\",\"endPinId\":\"pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_1\",\"rawStartPinId\":\"pin-type-component_902e1a76-96d0-4e30-b844-467374c96eb5_2\",\"rawEndPinId\":\"pin-type-component_d0a22dfe-53da-4559-b65d-0afb70497422_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-22.2820295000_-171.1770085000\\\",\\\"-22.2820295000_95.0021075000\\\",\\\"-327.5000000000_95.0021075000\\\"]}\"}"],"projectDescription":""}PK
     ˡ�Z               jsons/PK
     ˡ�Z1٭<7  <7     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"gear motor","category":["User Defined"],"id":"aa3e6a7d-1852-40d5-bd6a-bf11ddb1f8b8","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"e575fc9c-d7f1-4841-924b-9061a1257de8.png","iconPic":"b905cced-8669-4310-a345-cc026e3fb08c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"27.19180","numDisplayRows":"16.15562","pins":[{"uniquePinIdString":"0","positionMil":"583.50695,685.11343","isAnchorPin":true,"label":"+"},{"uniquePinIdString":"1","positionMil":"593.27584,871.33343","isAnchorPin":false,"label":"-"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"gear motor","category":["User Defined"],"id":"aa3e6a7d-1852-40d5-bd6a-bf11ddb1f8b8","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"e575fc9c-d7f1-4841-924b-9061a1257de8.png","iconPic":"b905cced-8669-4310-a345-cc026e3fb08c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"27.19180","numDisplayRows":"16.15562","pins":[{"uniquePinIdString":"0","positionMil":"583.50695,685.11343","isAnchorPin":true,"label":"+"},{"uniquePinIdString":"1","positionMil":"593.27584,871.33343","isAnchorPin":false,"label":"-"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"gear motor","category":["User Defined"],"id":"aa3e6a7d-1852-40d5-bd6a-bf11ddb1f8b8","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"e575fc9c-d7f1-4841-924b-9061a1257de8.png","iconPic":"b905cced-8669-4310-a345-cc026e3fb08c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"27.19180","numDisplayRows":"16.15562","pins":[{"uniquePinIdString":"0","positionMil":"583.50695,685.11343","isAnchorPin":true,"label":"+"},{"uniquePinIdString":"1","positionMil":"593.27584,871.33343","isAnchorPin":false,"label":"-"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"gear motor","category":["User Defined"],"id":"aa3e6a7d-1852-40d5-bd6a-bf11ddb1f8b8","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"e575fc9c-d7f1-4841-924b-9061a1257de8.png","iconPic":"b905cced-8669-4310-a345-cc026e3fb08c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"27.19180","numDisplayRows":"16.15562","pins":[{"uniquePinIdString":"0","positionMil":"583.50695,685.11343","isAnchorPin":true,"label":"+"},{"uniquePinIdString":"1","positionMil":"593.27584,871.33343","isAnchorPin":false,"label":"-"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"L298N DC motor driver","category":["Output"],"userDefined":false,"id":"7deca677-57aa-869d-46fd-8698e7333ef9","subtypeDescription":"","subtypePic":"dd9bac2c-35cc-4be2-808f-eb026b88f611.png","iconPic":"a657ee5f-a898-4bcf-bee9-a045b7cf922a.png","pinInfo":{"numDisplayCols":"16.92906","numDisplayRows":"16.92906","pins":[{"uniquePinIdString":"0","positionMil":"19.46101,643.40910","isAnchorPin":true,"label":"OUT1"},{"uniquePinIdString":"1","positionMil":"19.46101,456.50724","isAnchorPin":false,"label":"OUT2"},{"uniquePinIdString":"2","positionMil":"354.24748,17.92249","isAnchorPin":false,"label":"12V"},{"uniquePinIdString":"3","positionMil":"541.15242,17.92249","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"4","positionMil":"728.05734,17.92249","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"5","positionMil":"1676.39095,493.17462","isAnchorPin":false,"label":"OUT3"},{"uniquePinIdString":"6","positionMil":"1676.39095,680.08117","isAnchorPin":false,"label":"OUT4"},{"uniquePinIdString":"7","positionMil":"500.92991,479.46314","isAnchorPin":false,"label":"5V-ENA-JMP-I"},{"uniquePinIdString":"8","positionMil":"600.92962,479.46421","isAnchorPin":false,"label":"5V-ENA-JMP-O"},{"uniquePinIdString":"9","positionMil":"936.18245,220.17481","isAnchorPin":false,"label":"+5V-J1"},{"uniquePinIdString":"10","positionMil":"1436.18185,220.17481","isAnchorPin":false,"label":"+5V-J2"},{"uniquePinIdString":"11","positionMil":"936.18318,120.17343","isAnchorPin":false,"label":"ENA"},{"uniquePinIdString":"12","positionMil":"1036.18255,120.17343","isAnchorPin":false,"label":"IN1"},{"uniquePinIdString":"13","positionMil":"1136.18253,120.17343","isAnchorPin":false,"label":"IN2"},{"uniquePinIdString":"14","positionMil":"1236.18270,120.17343","isAnchorPin":false,"label":"IN3"},{"uniquePinIdString":"15","positionMil":"1336.18197,120.17343","isAnchorPin":false,"label":"IN4"},{"uniquePinIdString":"16","positionMil":"1436.18185,120.17343","isAnchorPin":false,"label":"ENB"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"DRI0002","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"DFRobot","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"ESP32 DEV KIT V1","category":["User Defined"],"id":"518495d5-e179-49dc-aafe-d7d40a222bea","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"dfc5a72c-0224-4495-b3b7-0d06b4ba9157.png","iconPic":"f159b6d4-7cee-4dce-98d3-76d280a06797.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"11.23521","numDisplayRows":"21.36983","pins":[{"uniquePinIdString":"0","positionMil":"1065.82667,1863.51027","isAnchorPin":true,"label":"GPI023"},{"uniquePinIdString":"1","positionMil":"47.22667,1857.91443","isAnchorPin":false,"label":"EN"},{"uniquePinIdString":"2","positionMil":"1057.65667,1759.30027","isAnchorPin":false,"label":"GPI022"},{"uniquePinIdString":"3","positionMil":"1062.40667,1664.20027","isAnchorPin":false,"label":"GPI01"},{"uniquePinIdString":"4","positionMil":"1062.40667,1569.09027","isAnchorPin":false,"label":"GPI03"},{"uniquePinIdString":"5","positionMil":"41.43271,1763.62839","isAnchorPin":false,"label":"GPI036"},{"uniquePinIdString":"6","positionMil":"46.19271,1649.06651","isAnchorPin":false,"label":"GPI039"},{"uniquePinIdString":"7","positionMil":"46.19271,1554.38839","isAnchorPin":false,"label":"GPI034"},{"uniquePinIdString":"8","positionMil":"56.13459,1466.33819","isAnchorPin":false,"label":"GPI035"},{"uniquePinIdString":"9","positionMil":"1058.24076,1465.94830","isAnchorPin":false,"label":"GPI021"},{"uniquePinIdString":"10","positionMil":"1063.08864,1364.05815","isAnchorPin":false,"label":"GPI19"},{"uniquePinIdString":"11","positionMil":"1063.08667,1257.32027","isAnchorPin":false,"label":"GPI018"},{"uniquePinIdString":"12","positionMil":"1058.23470,1155.42633","isAnchorPin":false,"label":"GPI05"},{"uniquePinIdString":"13","positionMil":"1067.94667,1058.39027","isAnchorPin":false,"label":"GPI017"},{"uniquePinIdString":"14","positionMil":"1063.09273,956.49830","isAnchorPin":false,"label":"GPI016"},{"uniquePinIdString":"15","positionMil":"1063.09470,854.60027","isAnchorPin":false,"label":"GPI04"},{"uniquePinIdString":"16","positionMil":"1058.23879,757.56027","isAnchorPin":false,"label":"GPI02"},{"uniquePinIdString":"17","positionMil":"1058.23667,655.67027","isAnchorPin":false,"label":"GPI015"},{"uniquePinIdString":"18","positionMil":"1058.24273,558.63027","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"19","positionMil":"1058.24076,451.88633","isAnchorPin":false,"label":"3,3V"},{"uniquePinIdString":"20","positionMil":"43.83667,1364.99027","isAnchorPin":false,"label":"GPI032"},{"uniquePinIdString":"21","positionMil":"53.77667,1258.94423","isAnchorPin":false,"label":"GPI033"},{"uniquePinIdString":"22","positionMil":"57.09251,1152.89631","isAnchorPin":false,"label":"GPI025"},{"uniquePinIdString":"23","positionMil":"47.14667,1053.48027","isAnchorPin":false,"label":"GPI026"},{"uniquePinIdString":"24","positionMil":"47.14667,947.43443","isAnchorPin":false,"label":"GPI027"},{"uniquePinIdString":"25","positionMil":"43.83667,854.64027","isAnchorPin":false,"label":"GPI014"},{"uniquePinIdString":"26","positionMil":"43.83667,748.59027","isAnchorPin":false,"label":"GPI012"},{"uniquePinIdString":"27","positionMil":"43.83667,650.76027","isAnchorPin":false,"label":"GPI013"},{"uniquePinIdString":"28","positionMil":"43.83271,548.02631","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"29","positionMil":"43.83479,438.66215","isAnchorPin":false,"label":"VIN"},{"uniquePinIdString":"30","positionMil":"553.16667,129.46027","isAnchorPin":false,"label":"Power Supply"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"HC-SR04 Ultrasonic Sensor","category":["User Defined"],"userDefined":true,"id":"f7a95729-a811-496b-83f5-7789de376adf","subtypeDescription":"","subtypePic":"5a738b76-89aa-4728-b8e5-f09c859dbb14.png","pinInfo":{"numDisplayCols":"17.75472","numDisplayRows":"9.29339","pins":[{"uniquePinIdString":"0","positionMil":"724.31191,21.31240","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"824.30674,21.31240","isAnchorPin":false,"label":"TRIG"},{"uniquePinIdString":"2","positionMil":"924.31190,21.34367","isAnchorPin":false,"label":"ECHO"},{"uniquePinIdString":"3","positionMil":"1024.30154,21.35407","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"SEN-15569","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"SparkFun","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"ba153158-cccd-4fb1-9320-38bebad1b7f9.png","componentVersion":2,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"ESP32-CAM","category":["User Defined"],"id":"3b4a66b1-0d1b-40c2-92f7-ec286f5c89ab","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"53de2a41-b288-4dfc-9a43-3e5c75810bf2.png","iconPic":"6590c6c2-4084-4043-8677-a67706af7572.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"28.68255","numDisplayRows":"28.68255","pins":[{"uniquePinIdString":"0","positionMil":"855.34971,2255.85937","isAnchorPin":true,"label":"5V"},{"uniquePinIdString":"1","positionMil":"843.65971,2119.07686","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"855.34971,1968.56623","isAnchorPin":false,"label":"OI12"},{"uniquePinIdString":"3","positionMil":"862.94346,1837.32934","isAnchorPin":false,"label":"OI13"},{"uniquePinIdString":"4","positionMil":"845.70784,1717.79245","isAnchorPin":false,"label":"IO15"},{"uniquePinIdString":"5","positionMil":"847.75597,1565.22369","isAnchorPin":false,"label":"IO14"},{"uniquePinIdString":"6","positionMil":"857.39784,1438.09306","isAnchorPin":false,"label":"IO2"},{"uniquePinIdString":"7","positionMil":"857.39784,1295.16617","isAnchorPin":false,"label":"IO1"},{"uniquePinIdString":"8","positionMil":"2093.68418,2267.54937","isAnchorPin":false,"label":"3V3"},{"uniquePinIdString":"9","positionMil":"2095.73230,2128.71873","isAnchorPin":false,"label":"IO16"},{"uniquePinIdString":"10","positionMil":"2097.78043,1987.84997","isAnchorPin":false,"label":"IO0"},{"uniquePinIdString":"11","positionMil":"2097.78043,1849.01934","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"12","positionMil":"2095.73230,1727.43433","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"13","positionMil":"2095.73230,1586.55557","isAnchorPin":false,"label":"UOR"},{"uniquePinIdString":"14","positionMil":"2095.73230,1436.04493","isAnchorPin":false,"label":"UOT"},{"uniquePinIdString":"15","positionMil":"2086.09043,1318.54617","isAnchorPin":false,"label":"GND/R"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"battery with holder","category":["User Defined"],"id":"d749d278-6a0d-4deb-825c-1b35ffc56ae5","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"f2dbd413-946a-4dd4-beb8-9b389826ae17.png","iconPic":"685e2fcc-e73c-46e4-a7b3-171ef11b9715.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"14.71453","numDisplayRows":"11.04227","pins":[{"uniquePinIdString":"0","positionMil":"648.23667,1099.67928","isAnchorPin":true,"label":"positive"},{"uniquePinIdString":"1","positionMil":"507.04667,1099.67928","isAnchorPin":false,"label":"negative"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"SG90 Servo Motr","category":["User Defined"],"id":"437e01f5-4fa2-4201-ac70-cfe748b41bde","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"7485d96b-ebc9-4409-ad2f-5f0bda14de1d.png","iconPic":"544a1249-aa5b-4970-8b42-188baf88f36b.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"13.63979","numDisplayRows":"10.67730","pins":[{"uniquePinIdString":"0","positionMil":"1331.78469,315.50100","isAnchorPin":true,"label":"PWM"},{"uniquePinIdString":"1","positionMil":"1293.62927,207.72501","isAnchorPin":false,"label":"+5V"},{"uniquePinIdString":"2","positionMil":"1268.88776,116.31101","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"9V Battery","category":["Power"],"userDefined":false,"id":"7dbe2b3d-2053-a5aa-7735-837175ae747c","subtypeDescription":"","subtypePic":"2cd57c9b-7217-4a6b-8577-1769ce4bee7a.png","iconPic":"1251016d-b52c-4e05-b483-3027638d0c75.png","pinInfo":{"numDisplayCols":"13.23181","numDisplayRows":"21.09330","pins":[{"uniquePinIdString":"0","positionMil":"1328.16711,1864.09428","isAnchorPin":true,"label":"-"},{"uniquePinIdString":"1","positionMil":"1328.16711,1964.08023","isAnchorPin":false,"label":"+"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"1321","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Adafruit Industries","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     ˡ�Z               images/PK
     ˡ�Z��7��$ �$ /   images/e575fc9c-d7f1-4841-924b-9061a1257de8.png�PNG

   IHDR  �  �   �@�   	pHYs  �  ��+  ��IDATx��y�wu�k<ӝ�fْeK��ll�I̐`g���4YiD�B^B&V֣��a�?������&@�JҴ	!1� ��`�X6�l�� ɒ5�,�^��5�������;�se����ֹ���U���=� �D"�H$Y@�D"�H$�H Q$�D"�H�#D�H$�D"Q�E"�H$�D=@�D"�H$�H Q$�D"�H�#D�H$�D"Q�E"�H$�D=@�D"�H$�H Q$�D"�H�#D�H$�D"Q�E"�H$�D=@�D"�H$�H Q$�D"�H�#D�H$�D"Q�E"�H$�D=@�D"�H$�H Q$�D"�H�#D�H$�D"Q�E"�H$�D=@�D"�H$�H Q$�D"�H�#D�H$�D"Q�E"�H$�D=@�D"�H$�H Q$�D"�H�#D�H$�D"Q�E"�H$�D=@�D"�H$�H Q$�D"�H�#D�H$�D"Q�E"�H$�D=@�D"�H$�H Q$�D"�H�#D�H$�D"Q�E"�H$�D=@�D"�H$�H Q$�D"�H�#D�H$�D"Q�E"�H$�D=@�D"�H$�H Q$�D"�H�#D�H$�D"Q�E"���Dy����w�;88��j5'C��}��ɓ���ܜ�C���$Ir����8Η/_��<3�(����j�}~���g��d �^�@�D�W� �ݻw{�O�vڼv����u?�cǎ�ɟ������`���� ��C��;�N��4w�ф�rp�+�J��%8E�Q�ZM�,K�&� TfN�g�}v��_��n���-[��g��Ț�fF y�5פ�"�k[�"�H�#�����*���'>�5gΜYv����X��y������*�w!n2��j�� �2D�>q}��s]�p ������	�b�pH�d%t]܆��|���:��Ɠ��g��h4	T;�N��n��9����˗O-Y��u���x�7ܐ�H$zMH Q$�^Amٲś��� @5ph�ZY�iU���_����ӧ�?~|�ɓ'��uW�:�8��J"�y�YC���É\����p]>�G��ef>�'L�8�u	(q��������du��E�?��Ab�Z��mO9�t��I����?���ccc�|nhh����6oޜ�H$��� �H$��2A��ھ}�F�n�z�s�=���FH[�����Q����UCت{�7�S�,��A����9�'�-�9\�?	�h9� }'!|������ş�M�Z��i��h����F��r�I� <f���iE	Yq~���D�xj``���z�~z���Go��ck֬�D�l�:ц:4�H$zUK Q$�~@=��C�_|qp�Ν+��/��
�NLL,E [�@u	��
�j� ���\J:�XA5�4���h�}_Lf;��w���-헎a�k�c���(-��i��x�.^M�]�y#�:�h��3F��p�������<.[���G>��,Y��Moz��KS��"ѫO�"�H�]�`���}g푣�,=y���?cAT���/.C@\s�رu�gggG��v+��j!��g`��qF:F���!�d��d��f���6�l8��m�Oے�of]�朌���q�SWA ���1H��n�����h������=���}�c;444t��?��?j��'b�H�C� �H$���l�R{�F>�O\|`߾�<x��ɉ3�4F&�"<���BU��@�E��k � ��$�r�]LZ�ܙ��@φK0�2�Umֱ!�>�_{�2��[�vAp����X�dj�O�sD���3�3�s��)��4�իW�ڻw�#�����������E��E"�����ʎ;F8��O�S?5qfb]��!�C�) d.C�@���i;��1$�NdY3Pe�І<X�z���A{]̌lˡ�r��b[+���U�>'��|�<�uȚ}W������A\P&�_���#8�ejj��zꩣ������_��W��'?�s�ƍ��7o��H�C� �H$i�t�M�fsb���ӗ�S��-�3�W�����̙3k���B.-C�L�/]��o@Ge�2�� H�ݶv��.�]9��Ӷ���m��g��bV��~͹���5 J2q���dm��q�����m�_C�^:==}���Bsvv����������o����+V�x�����|�Cj�H$zE%�(�^�ڶm����۽���n���33W��-N,�:I�
Q����`�����,e𡉀� "Y	��������A�i]ڏ��b��`i/' 3@Z�B.'����`jæQ��[f{��Rj�QޏNh)������O�iL	��;������}��l��>}zéS�~�?s���=ǎ��#��7���#��gA$�"@�D�;Q���ݻ���k�����}Ǔ۟����+�]~���x^�l��8ǢW��3d��}v��Y�$��D{2�h���n6pf��Ҷ�cmb?ˢ���V6�~��1�6�m�7.w�/S�qvv����un#��]����ɵ�o{��>��3�|�����������Ǐ��_}*1�"��#D�H����9|�p��/~q�#>��w����c�bnnv%BJ����j21�v	�<�t4��i�Ģ��y��A�����Ō�����3���G2�m뢙_�,��W?��g�����������Fc4�躌�_�5A��M���@�9����|4cd�ͳ �����\��Ol8q�Ļ~��=�F�Yʧn���?��O���祫�H�I Q$��Eū������g.9���C�����_wz����3U�;y�� �̷!���k�Ǭc2�� g����'�u�>������|�goS�K,�_>���Ěs7 l[!�q�����M�;!�t�1�l\�e�)�"Y'&&.k6��0|W�Z�:}��>Խ�<�̃�g����nڴ)�H�=K Q$�&En������=��GX��s{�޵s�N�<y����ҹ��j� b��m7��0��lH���N��l/�TR�9$����$�>��b�|�/{?���� �߾͹�a�V{L�}�w��6d�kٺj$�t:u���Z��G������۳gϽ���۾��/?�v�ډ����R2G$�$�(�^SB��v��]��׿��{�~�޽{~���ޜ�مK����� �����9	&.�'H6����-'��� R�rqj[�,|������~�5�([$�����l(>�ճ��ʙ�v���F�]��@ڀ�OI�Ënc8����[n�����G֬Y�q���~������tn�^B�"��5!�F>s����O�i����8v�صǏ��'O\�020<<욞��j��+4PH2�r4߆���v������g���c����ŀ����s����藥L����lA4��춗������Ff}ݽŀ�3;;;���aq=�}É'��ر�;۷o߁��Aq�<� ��J Q$�X�On��%����w>s���1==����f�I�M���A��X����DVąf�(^MR I0i�{���ed����v��Pc[��ֵ>�������/�g�^
(˖Ǘ:��� �VS#S��#�cc�`�.i{,ͽ�y�M�O��֥�i� ��ƙ���v���'�9�u�޽�oݺ����Լ��Ε �H$��Ֆ-[�>�_�k�s7�9}�����03|�N&vB��Zf��Ui�n�qe.��x���4�V�uZV9��e7tYeX;�;����\���g��}}�m��T.�c���8��0��@���.6N?
�}�:�u\}���Ĳ�~������駟~tժU�|�s��;:::%�(u%�(�~�t���{�o�ԧ��ϝ��|k�ռad��дw���/���;Y���H.L�f�� "m��;'��X���-4ꗌB*�ٙ�,��]�5l�}71���~����l`=��f]{������e'�ۺhog�OpH��Ʒ!��J����n�Z�KN�8���ѣ��1~����/���n��w��/J��H Q$���#�۷oͭ�����٧����or=o��hT��Ƹv��9d�"ˠ��ԪKh�g�T�Ԋ�C�ѣ8f
m���D��e��W���J[�ę$���u�p�VA�\�/'��w�K��,w�y#���x���=��>N�Ua�S��V�纜�h4 g,����/k��7�f����FQ�Ѫ�Hŷ�i�Zs�:��5y�knf걣���>������'@$zK Q$��e�_�K�����gv�����8=qf�|�;��'�"�@A��,�l��ƴ9E+�~ dbK�0I����ӂ�~�ī�l=ǳ��ŏ�u��Ҿz��6$�۝�D��m�����w��w�^@,[�� �j1����bD��,7!���UπS��*�z}I�#��x��񟜜:{�����������͛����u)D�H���֭[����'���S;~��p~~�b|����ǽɳg#����d[�������C�0a,wv����-�d��HE�\��X��J���\	
����-�/�SX��S�S�Z��&�d�N̘�zR�fT�%Ϙlnk'��1�����<edيXޟ���E�t�1?
�}WaAPڰo,ʔ���O�j���8�*����Ϝ�د���q������k��u'D�H��Ԯ-[�[�|r�g?�7�r���w�;���E>��E�C��l��Ohb���pv�D�g��R��$��r�]9�Ў�[�vf�����G�9�rb��.@9s�)����|����*/x@VD�]�s��q1�����]��;�sk=��ؖ��:f�]~��W�m=7*�.�u͏^�S��[299��;��ƥO=��}�����.������ߝ��u"D�H������<����g�z��;~�'�s#��fg�~��(J��V#���l`+[�H&�I�\�6$�K�0���$�,�Y��_��Z����ؾ�u�����y�q#;ʦ�(�!�z�9`���\�0���n2��6�S_�����.��K)������s\,�����n�ж��i�ݽŶ�EpTggg�<}�ԆCG_����������k�^z�s��׃E"ѫB���<x���}����}Ͽ_������<R�ՊVl&����k�X�+��.Z��R��B#�z�\��|��ﶵ��Nz]����D�~�WےXfK3[&�P}���뉊1TVB�Yώ��~���܅�b�.��U��]��8K�ɞ8�E���:�ޙ���o����?H��T$+u��r�Y��3x����]�w߸|�#���������ޱ�}�{߬#ŶE�Q	 �D��v���r�-���sϻ�o�ff����j���p}�p�Tǔ��E�D)��Q���\?���B������o_x0@�X�� ��Ьg��T�!w��l[݊$��}�y�]˼e�z��d������KYԹ�f���:خi�� ]ލ~,V3q�fl5����\+��b���������]�ű  �*������G�C����)�3�^����V���ٹ�oݱ����{�������w~G���^s@�D?2��������m��z�S�<����qnnv���03� h���N�^Q/���5%gʮIcI4 g�#��1�f]�YD3��ͬ�}?w4�K�Y��7�������$b��ʊXާ�^6�gΣ���s�}�λ|}����|	+��.vO�m�g�|�K��-&Ԁ���mS}L�ixnv�N��aaz�g����w�b�>��7A$z�H Q$�HDVÿ����?���z���:{���_a�`��E,Ya	r(���h��^F��X2��E4�h�����O��jϷu�ze}7�dg:�몘�n�@���b-v�lt܌׵ύ/�������:���Zs0�Knn�HFQך��Az��)�K�_c%��Z�瞶�=�����b�{3ߎ���!zV�4�珬�a���4q�nI#\�e�d�����LMM\~�С�.������/�eۇ�����5 D�H�CY��o��w_��z��_8q�SgϮƗu`�8�Y�
.�@����.^#h����$��B�fy?���,f�]�ZnovsY���[�P����e6g=��OU�:�9��s6����e�ۆІB>�r�N���r�8�t����o1��b�-fy-èy6Hvr���`�Q���q����a�kZ���С�������?���>vD�s	 �D���j�?�����#^�g��LLM]���F�H�L�n�mm�u��b^�vV2oc�x�e�.�4���炇��^h,,TE�r��Y&3!zy7���r��K�dY�1�E��7�0��NYSU��QVE���v�h��ME�S�y�kK~�-��}QVG�{ea,�!�'��ӹ�f^)-v?�}7�gci���Y4�h��ϙI�JS��4���{ӳ���X��n��g��{��i�9O��H�*� �H$��衇��×�x��o�˯<t��q�ڠV'�a�	�.S���W��ۛq�XF�b��d�C?�^?���r�a(����45u�z�om����)<����5-v�ݷ9����Mlbnܻ%W.��c�IN4�9הW����斫�Xվ{ǲw�R�ɺ.�e?����������17[fP�f[�cÁf����g�f/ۻw�G*����|m۶m������U�"���p��|�+�_���߱��G���C?�j.,C*���rñ�A�@Y�tF���V;U��٬c\��Ɲ3�n��q��|���������W���
"M�M��L1E�*�����R�$7�sn�X�[�-��sA��]:Nz{B�27����8z�鱬&�H�)��9��y)�17VQ x	<�U���@y|�Y{�����T�a��%�LQ���9��7�jnؽk�LOM-��:���u�nh�H�c&D�H�i۶m��7����m�v�s{��onv�j�=�%:[�Jh0n�nW�^�*���Y���~�`܄����e�pR����s��&��9�ˡ:�����z��@6��u�D���d���+����d�̻�h��r=gNyJ�Hu5��<Vp��z��Յ�{FL_�U�ⶶ-�/�����}y����1`[�U{=3U�5��Rt��+!=�����ڃ����ܲ(�����w?pջ߽ "я�E"�+��۷[��z�SO<���xW��!�TȢH "\,�c�"��ϸ�e�R����l�Լ��U�^ˠmq*�{y���_��X����䥬V� gf������CkaLr����z�0��B�ϰ�����)`ת�U�N���d�<]G��7�5%	A�?Ms��lx�\C�]�r@�XUt����X�`.���軁�~���T��$;��n�G���2�/M�~�1��:^��^��ٍ[�~k��c#[�|~��Ϳ'�+�	 �D��][�l	o������֝87��N����Z��(s6�E�iv��ś�@]O����xI�\����</���K�ap���M�ky,��nY���I�k��?1��ΔU��SYv���|B��K��T�0_W������\pXp��(��A�gT �� *�=�S+8�Op^���~���✠�S��v�,�>��d�4���N
�k5[�>$��' j�gn����G�5�c�`���@6s��Lh���+��3�I�(��;)�%�e�4���vQ���GF��l��吺�PXY���^�t��vg������ԩǏ�xr�S���^x�͛7����^�@�D/����x�}����g��� �QnE��p i8T�&�~���䑕
��D�R �a����U��
�<)���2�e�
'��D:��B�$�>ˣyԭ��]O�0�c�i�2ܹ:�#�D�GwB��d��Gn[�N��@vg*C����6�n�|��r��FGFGG*P�;P�.�^u5��!���趯S�A1n�,
P6q�Q�!�eG�0�@'Bhl,, �3��!H���L�9�#�:4R�m�'!$N�ڇ���
�K��ǮV�K�1A�oz"�Z�sN\7�U�r*�����<N�c��b"��@Y:5 �v���c@��U�<8�N�a �Bu�u"�@�ݾπ$����vR}g8>
9�6��z�1p�ԙk^�x`�̙�5?�S������w_{�1�D�b	 �D��M��z������xj�P��
N�GY�TJ$�&����4/T�%K�*zm����5�z3���%�mn[��.7uu=;���P�.Zͭ�<O�2�u�E]k���t�*>��J]� eZ�-��(��CE|�1�@�ˠZq���d$��F�k0<R���
Bac#>�j4j)4�~���.� �W�Q�1�J�ףd�������H����D#����qU���,pݐ?�b�8%ޛAH�Y=�[�Lu`j.�3M�f8sjN��F�L,=��ǔ��|��,�!�b���eʲ�`��/ck��x-.u������:���(A�J�&��1��s^�&ƽ\[1�}w�XP��Ÿ�����ι�nam�"mdz��.,�l%I��:;�=�579r��L�{�GQ�o�܎k���@��U+D�H������sK�u�?����=��g�N^�h4
�"���m츺cIEYmLM9jkFVF���ح�L�a�pqo\�zi'��[�`q*��ae�����W)��#�:
:�HA�Ӎy$�#y1��*�$��P1Su	��D.�8�����y���b�Lat`��*��d0<��p#C)�q�F-��:�!��}� �1"p �k
����]{�_Z'� ���Kq�rI����-L����+�,�
���Lo�;��2rE{lml�bXh����υf����`z&��Y'�	g���/��A茳���� ���qFp�s�s�IW���z�y��c�=�����:1��d^�����*���'�����D��Le�r�y^��f��b��Ses\��!Au>�8�V>|�}Q�4�8��-[߼ys"ѫP�"��� ��~��^��-���3O=���3k�0`�Z�c��3�^�m�G����b٣vR�7fr��ͽ��n�f���CG��quQ�c����8AHu�)��0�n]e5r�RI�b��z�B���oh���a���X:^�����y�di��G"v+����GD
I���6*w��se�"�*u�,p�.���(��|�v.N�-�M�X�g�,d:Vf����U��a�@.|]Z�����!�S Q'��&�&pf�S�9?т��/�J�1DQ��V�(u�����d5���~�sPuCȣD�<�.���{=]�Q� �V��ӌ�WQq���L�x�hh��s@����/{��7���g��p��q�) �~�T*�&��=;��=�H���q������Wz8�^u@�D߷�l�������K������޽�o������~>�S��Y��<]��@"��E]��Y�@���lf���^؎g��
b����&#���z\����n�ݐ.��Ւ\�i�VJ���9Mq��
YcX��˖�jy�#,_���.�#v�~�0�G�N���Վ��,M�{5���/#�1x�Z����(��2.��/#�^oP���}8vI��p;����tZ�cH1�DY�&�}9�dad�A�O+�7�S��;���9\r�� ؊���,��3�x��^<��&���&�4*������'��b3	�����PrGq��&���2�br����.��� ���Ԋn$�>#�g�lY�?m��RY�׫�dI�g�,����^x�m��6|�ؑ��җ�t�o��o�9�yE�*� �H$��Del�v�m��ܱ��<�o�%�jpp�/�.��P5t��/U��Ɏ�3��5�-t������{����8&����
�8AHt63-��!������`��;(9%K[�%���	��spax�G(�a�xK�d�rE ^%.�&���4���	��ժ9��00Sҋ
ݢ��1��:���u�,���5	=�U�AP�XX3����q�X����"��uu�b���S�O�aG���\��gw\�kiTp!��C�*�b �	�:Y�Sg�L8���N�iB��A�Pp�i7�ד���v9����HR��ޓ��BVQ�}�Tg��l%�(�Y0��<+B�e�����Y.�c�M���bH�r��2���l?���v���L���������q
�K���U!D�H�=k׮-����?�i��w~�̙�_H�l�����'��S��3A��[��� `��~�B�:�Z��ϲ^��̋��������s�ʒǖ5�Xy	'D�.�B�A1��� C�F�<Na�*V.�aժ
���0:���H�m����EM��T���)[:i�����:�
h�H�Lr�ss���G�q)�0j���~P_�klyb�c���z?ڢƇ񂞬]3�
v "��U�=v�V�t�(�Q��A��
��`�t�
����M^������K��S��� =�����m�*$�r�����L�0���T�����s�$p�d��Gx)����Az�i+"M����8�O�G4?�L<(%XK7�#A���p2����@1��˟y��?���]�0��m۶��|�W�E"���]�v������{����O��_��j��K/�fS�� w� �`כ-j�)EM>Bl�L$��b��\�NQ3O�$TLS���{��BV;�HN)��X�@�V4�lb�Vt-�U" X�܁uk�`��
�]�²�FF(��:�t ��(-�g�̫�v��@�uɂG%}|�J�H��#��P�O��c�7�8B�:��U�2Q�����X�3m	�]� ���s��"��UUg
�04��^w�nf9֦�H��c�nS*��C@ ��*��|u �á"/�v��K�aúA��lN�N���?Ԅ#ǚpvʅ�Y���S������>���9{������U�O��ŉ�\[\�:(y%7��������gA�׷-�fR�jY���^�N��h�ڨ[p�ɉ�߽��y�������ۻaÆ�D?B	 �D��Z�w������ͻ?t��w!�-��K�Y�hR�D%K�]�ٶ �Y�v?eci���2@��v4h:�֡�;�u��-v�"�3�v���U�m��ȍ�j�<U�i+�ފOei�ad8����0�W�p�*�XVeK��@�O�$3�`B�Gu����Ɠ�R/*	�3��&`��0�!�S�q����)�ͳ�U��N�I��%��²���&���&٧���PM>���U���n�����fm��{�-�J��M����T��O�S��9�E�d腀��ޣ��-�a�� W��G��p��;p�h/��`�K�Fp�pB*��C�+���=*�C���B%f2�r��׬LT��:R�c̵8�Ϥ�Y�9��X.�n�˚g�+�c�s��uc�	�;��� <��o�q{�j����Cm������G$D�H�]i߾}�;�����C�z��Gi����[��q�ƊH*w�0Y��;��.uSN辠Sm!����i_�#U�".�M���&)�j��H)t��'��������|� ֭���q�0�F5Q I�B/e4����]c�����M����[�(�O�)���2ڵ�'\�1�B@��8]����&�(�|��{��L:�22&�EՒ� �\��o��S;w2��-�]��RI�W�"��Q�MC�/�:�I.}� S�906Z��+`�ـÇ8~<���b8r�'N���b Bb
��4O��A���3 R�E��r�"�`O�a���}9���KY�-�!�v?���{���ҍ�hՑ�G�_�����B��w�u��7�x�$��~$@�D/�m۶U�����O>�[Ǐ�|ѭ�����L�7R��*�Y�x�u�uI�����9��SwK���c|Bp�b˾���c��3"+�dg4�z�4/�@�0>�����:\�`)~_�?G����"d�*O�;v��,KtݝL!����ֱ���|��/�7󸈌3�ef��X3���1d�����.��n�9�cT5sx���M����T��81Y�i� �f9�oE]C�jw��W���g&Y�$���k>F�?$t�̣�B�B��p��0:��}���9;�� G�%p��L�m��<>wy�
�}5��T���u9Mu�u�ʵ.��;����,wz��9W��#�O���7����U ��`Y�Exq���رc��d���W9rd����_��+��E"�yu�����_����7�篯V��W�kQ�5J�@
 �3�B���)Kc���-��`�Xi;��׃n�f��Nye�E�ץu�dw?�x�DY��
Sb���P�`t}X��
�n�úunA��@��@�ms��Ó��3�
�P��������gV���2V�"
�r��Uf~vz�r�+�(�� �+.��Pb��ku�W�/�ry�"�;/,�\��\��.0�����<��)��3��Q) eI����ȹ���?��\�:J�����zh;�1���c�)^q܁%#x?.��7���c1�{~�j��G�05A��#��p/H��N�?�w�Z�*��)F�kW*{�u�s�l-��\��T�(� r3�9R|"-���FϜ9��'����쳗�۷���#�n��"�I�"�hQ�}�ݍ[n���>��C�n���Y���J|�-L*��(���>��Ь>�4�ʙ���=��g�����*WC����AH�P���;��بk/������q}�-�al��M��)��Y���~1F9��vc��A���
��"�عi�~�%�mo�#�:Фz��@E��(q�i����u0�!�F.X�-$���U�ό>)+�U�J���M��>�����x�C�ff�lQTe��K�-�.[Ȕ+�XP2���R,&��h*�{ε��	�)��O�^E0ҨÊ�֬����;��:Ԅ������
�SY�@�ǲ�:W�\h���HY��ű�=[v����=���k�Sl"��2��5gnn��?�6M�L/I�g�����lٲ�͛7K\��"D�H�WT�����[������Ͽ�V�FQ�Ћ�^hd�XH�����&�|���h�&�A���,��JG�?Wn�n�.��rru"!Ρ��Q���E� �i�r��7���EU`�x�p���s����S���u� /�|�h�������&�$e�uu��O��s�q�j�LѦ�#+u�xQNn�>�Xe6Sl�鎩D����R*/db-s� F�(�c"�����A!*�8ʰ�C��B��A�噾����e+�m�tK� � ���':�?��i��u["�5�xOָ�_IF-���3{�]7e��2Ai���F���ʅ%+BX�&�K�%�_�A��6����5D�3��g>�<�D�,-�>~)��m=\�-��ϯ��X��3�ă���\q����{|���f���u�]��=�g�+.D�Ht�n��&�_��Տ?�п���|;�����y�
\��s�%�3
M&q�n?F2��n�~�(Fe�J���Tt:F��sl �)�U�*���`֭��͛R��B.X�C����Cl"���y��ʒG����c�� �ל��naIT�9��[�%z;]��\�p\��U*�ǎ��K�z9Sl 3v�5�A�s9"1�����U?���N �@�c�[�P��#�2ΤI�3h:0<���HA��.&�$��Ǎ���7������� ��?�F�=trS)G];�?V�Y)����HU/i7�\�zJ�\��e�Lip�ۃ� �j�~i�������g�q��*��`�JՋ��}tM�.��Z	3��r��b.�~�F�1)B��_S�Ie�g�>��D�`�̴i���F۝��O>�8�4����c�~���(zE%�(�����{����w��l_V����:���M)�AUBڸ�}��i�g�О�:q$��b�p������Q�Z�u���K�Ո�����0�E0�`�r�u�F�W��K�p�	l��Ei#%�[��bQ�>Y =�\BpH��b�R��Km	&3��a�暔����DF�$F�A�I��}1}�������Y�jhtx=��c�C$"%�d�E��<tV\�O�P)6�k�Sq�D�K*�C�o�,��%���jn.t �h���H��U*8U�2z\�'��ly��C�O�F!��=eE�ٮD��vrb�Y�~�Z�"�e��'�s�"к-<�6#$�s96V�e+F������N���p< ��xn���1��ך�$�څ�Y%��s���*����qoy!�YU��(���LeTs(D���sss���������`c8s������{���%�Y�JJ Q$�蓟��w���/��������*��$���!��(N�s��k^t��7OuL��n����#�"�)�8X���$��O�<(�ϴ�#�勬O���%\��+�!DmG�#���0>���� Woj�%k=X6>��|���^�T��]|��8�R����)9��=N<!�h2_g\������D�?s��q��v����)��)����d5L�e�'���r��g?H�!�ȱ��ZAYau,"er[�-�B���eh�9i��8��R��� �Fl�L�*,�x�YPǊ)>�,��Ù����Vr��*u�!~�:T#2�����4j[dA�b�'��d��4��O������>��aMs��j�G���=/-�4a�j�}X1������8=���X��y˵��^�s�CSG����$t�)��|�w���}N<5�^�J�/��q�� v�I�c���%3�_���ۙ�8��}�֪t�N�Cg&�~a�����z뭟Ɲ΂H�
I Q$��3�Y~�֭��ĉ_@^��H�4-�M�!����^~\e�J\1���7[��u��4ΐ5��������������q�a�L��e)��rn��J�j6���e����K�x�b�;���6��sP��nq�0T��~"mj�%j3W�9��1����QI�C��Љ���R�0�����r�maD0�9F/P�F���520rp�W����ʂ��/*x��FE�3]ew�:1�!���-7��R��@IY,�&��CT��()�LD=���'#��0��(6%5�e� ��00� ���.~wx]�O��!=+1Y{}�W� ���Sk�L��1pLR�qԳAY�Ɣ�^A��Po�FƆj�n� �XV�Vw`��8��i�m�Izx�5�/'���{�?~:���H�j|�T/��̔�u�,�-�� }ҿ
�g4�K��K&�&��~`˖-�m޼Yz7�^	 �D"������o����������N&K�qۙ�v̕�۰�5����
���g�?eI�V�\Er��\��e�A���SU�s��"�g��h�s��/y|<�u�p��!b���#�P,[�e��uɸU|�r��[6 ��A'Ť��������OE)tڔ9�ɹ1���Lbj���\��3��p���=q�:���]:��w��3ݩ%g���Z��k,�[_��w�-{�i�����n��ȍBc��C�V��;o�Q�q�B�&�����5r�Gx�Q��d�Ͻ�BX��z�q�{Pm�P���N�.h>2Y�yݤ�aW%<�n2�놞N�I����EP�����7���5,� `ǎ)���L����5�No�����Vh�<nH�< :�\� �>�c��:9�뉩,r_Lvf��n�cu�$.;&�~����n|�'>t��?��9"�+ D�Hw�uW��_�������<�/��Makzqk��-�j=/<;�ܟ�\8X���tl��1�4$�ucD�ѧ-G�b��`7cW�K-�p=?�`���5��ɛ��ի2� t8C�@�
gs�ƴ]�(6YȜ���-��,U�cr�s.0����b_�`'S�B�[��w`�"~ʹ�B�C��u���� ��/��3c]��<mALM�o�#�7�\Ւ���k�'_A��������>+܇Z�'����pr��]�s8�d)� ��9��U{C�2�].�u�AՆ��t��V�U��p�>�� Y�Cx'�� �QL`�������{P��,��zN�EYަd$WwJ�2@�B'���k��%K�t�,�~�'OL��\�|�4�PJ�:rg�XGU<R]W1�\)�t�����/�\�� ��@"�풦[��=�N�<y���v�x��w���w�{D��Y�"��\�߾뮷>��]u�\�V=z	Q�^Sz#�=eM��)Y T�N���q��L��b&�`���.��:B��z]�%�����<q1g��h�b�d+SW\�Z�+�.Y�/��e�k�j%���@��*�����1w`���T!�����lU�>G��Kũ�T%�P�I�J�2�j&i �$�D�af�$�h���q��q�&���v;V����4�
}�[�ܢ� %�xz�ݶwdU Knl+cAtM��F?�B�9~��xA���y�UIG�(��;�X�<�v�ER��
�sw*$�D\����5Sh��"@��"�Նp���*#ٯ��;a�Lɢ皎;��ٺK�@er�\u�avWYA����s�J�@M����a|d9��`v>s
v�o���y���>#5�V'f��K.���͜���N�߽X��~�F�E�����J��zF�u�`��s��gv�ᝍ�M�q��z�{����e� �H�:֮]���~��oy��G�pff�ma֩H/��H��|1Q ���\�y��Ѹ��ˎ�罖C3y`�S;:W�p��vvcea̻5�8��R�P��`x��/~�+/�MpɅ�XJ�4~�bjcW�����-T$9�5z����^��J�`(TP#��Q
mr!#v�R�Bz�'VJ��[��5��:C7-J�(���-�?��^�QI(��vP�lm�%y8�M�)�tL�"�K�!�1���:fҴ�SH��4��I2��*�3�fM�!�
�vPQqrT�Q[ςJ]3͔�0U�v,G���ʩ6)���|�oރ��j�4�1T�C��%]dW�-�LX=;\6(S��q.�=��G���R�����׿t"d�ή^�j����������wR��9;�ی��AHn~W M=ݎ�h�]�2��������|��o��r������?Lt\/�ԩSW<��C�W�W�=�e���&E�E/�E�שt!�|��ߝ:;u=��0�|Sj�����\U����L�C�H����\���q��lf��
���R�mL�P�J��d���V��yDN�j�H<!���!l�ă�߀ӥ>�Y��PЁ
��!�H%�O���U�)k����V�Lg�2�Q�Dr7:\�/�ȍL��T�F*��і?W��)~�ݎ9ՈT��&VOi�����4.�QVp����Յ�Ml!��jmS�#�?$�۵@�M��#��| �8C�D�f�zK�}A�TD�sO�q�5:�����{��`SU]�����S���x��c�àȖS���5tf�݁Z`p��)��0>cՀ-�TN	I_6�|��7Tn��Qe�5�Nnɹt?W��Y�cC�]���A\��=1�}����vB���P,�)�d�LŸ*{s�ϠcL�p����|	)��g�ӿ7SG��3��$�c����[���~�Ҩ���G7m��H�2H Q$z
_,���'��{�=��p����Gt��6�=Q�j�Z�5/7��!�J�p};)ņC�U��y�y�*֐�J�t�\���q�.�h	"�=�{�֭�å*��
.Y���-h�M�b���/W�<$ASGY8���5�5]Mv�:�l-���n%�i#^��nd��ⱅ�˗p�A��X�+0ׅ��ug�.�L��tn�-b/#�~�l=ʬq��C�n9�:S��0��f�v)�2<\�TY���r�� Y���x�*x�$vl	tT�)�-�N(\,�s�B�@�f�&�\�!���U�ᐲ�))�N��M2pH�Ӑp�?`�=�ss!��4��h�c���H�q=�����ĝ\��T��Y��6�U�
��#��M���@�F8�mh�<�h� x�v`�҄�;�p��4̵����*�#�'N7YH���֜��z��m�1��j.����]ˢ�9��z�x_��7>��O>ub��q�^�^	 �D�C}���]��o|�9tc�^_�/B���6�,D�t`<�� ʟ�V�p�s�[���qI�33I���&#�[Tu� �0z��	A���m�J�\�����z�V�/������K��y̙�T�/�ɱ��@�b�0�~é��0�z�NT(���t.*A�SE�]W���t�`�@Q'[����$�VG���P99���q�uɺ�nl�*f�<Y%S�|� ��8?��z�ʈvu�>DJJ8%9�:lM����ww	�\�zU#�ѹj�T�U�2D�1ױ�d���u?fU��4T�[��Ԙp��T�R��v[��:����5=sT��?��l��l�CTW1b�3���Z�1컁�AT'Ay�j����w3'��^�����`�Pc�Ò�#���ư�`f�.�n���?T���T�2��J�(q��7?h�+�~���~]�̺�6f�i]i���o�$��7�o߾w��?r��;�<�K��KS ��@�^g��;����w;�¯�Kg]���fS�кn,
��[��6Hi�sX�l�W�ʙ�1�0o��h˙��G��U��O�fm|�/��po��ux� V.�y�d%�9VQ��V`�+w��P�q��Ԙ�V@�E����I[���4��/�6?dA�\ݵE��t}B��9�	�C0�L�W�.[�T$���>8V��D[��~a���p��B-� 7����=r���p�S�8�k��08�>0'�,�����-}�E������>@Y��XEd��&���;G<�E��ȜV�mԶ��1e��E䐃�Ӯb����e
�SI7�`&��jۚ�+�ZBb �F�qg���"�ʍ�sAw��J�cA�⯸4�N�0�#h9Ӱn��_���h���=��>QBez�\\���?�dBq�>��w��gɗZG�V�~��eِh��*�N��z�v{́�~��{�=z��wK2�E?�E�ב(����]����>77�������kH��S��h.� �L�.g��FL���)�!\ ��� "����C	�b�He�mG�(BD2�3W�[��X���M����*p�R��|F�j糥('�!�S�T,��z�'���X��sE�C{!g�!'���1���:�O����yT�W��%I�wT�u\�B�EPnPNIu9���]�4^�� ǻ�����q�Ǥ��{9��sC��Ql#Y�dK�p?h?0��rv��-�3�s�ܦ���:�� U�IW��v��.\��S���WpU.���5W�hj�
WY.m�̴�X�5T�ڸ�y�"����� ZY��j.�"Ok6��� ��M��J."sf��=�[T��	GN^$ 3�ᝇ*t �֫Pp�:P�j#��{#8y�	YG0ԳM�9�/u���>�vR��LBIٽ\�v^,�X�[��yZ��K�$<q��߹�FG���{dÆ��O	 �D�Q��'?�ɋ�}zׯ"��Z�Fq쐫�\0��!���,f�>�]hf}�¥\v�Y�� �:g�K0����ɱr��$Z�N&�<��#X�$�M���WUa�FV.�D�)H�b�Y�T;�,��*�bj���d ��Ǎ=n���j1Ʊ*S��dG%(p��"IA�V�� M�0��$c2�ݷ�,s*)Ee�5'YVX�BO��2���e���v��lcO�����&3^��Z����(%g/�K����ZQ���T�O��g�r�i� ����R�gJt�|���ͮ)	��q9�G�c �Qm��,�x&�&c��d����I��9+�oC᪦��Wa��~ԩ*_�ieМ�`v>�!|&�@��5-���b+U�"c�Tu3�e���אv����9�[0:�?>�8C�X2ځǞ��/��ܼ��� Ǳ��9m+5h�Mƻ�3�
ɛ���{,��ᰟ�݆Cs��>��`��l;z�O<����V������,�>%�(�N�w���|�[�9���|�b�(�@дѣ�%"T�eh�u]�iO<��Ŋ`�-��J�]~�j[G5<�םY8�߸3P	T}�+�0׽e.�؃��i���3�ġ~sG  �:���ٯ\�P��oj�u0N!n�u�us�T�?f R1��6cVX�R$�N���v|���u��cJ�d�us�G��vt����{/;�}���*AR	�����'L�1�ƎWm�n�'��2ﴓ�g���O���j�=��+�$���d����I�c�Sr
'�@�w�TR� ׻tU/����W�3**��
��q$R�nS%ƴ���p��0�.zP٩*J�jT*�.[33��L�Wq��CxFC����JHQ�n�s�,jlO[q�u����\T2�Y�:00� � �Z���Ν<�	�zȹl��*�D���C����p����Z�5���i�/L��c�;��V�Y�/?t��/o��I����&/�H�}H Q$zh˖-�?��?�ā}��|�����@���K�`� ��=4��$�lbg+/��ζ����5��. �\�0��88_¾� �V\uy���֥02��2�0ц�k�d�u��L���9!�b�<e�Q.j�HA`�if��.�z��$\ߎX���{#+����L����~�m鸎��
Kg�u�K�v��]��D��%�(+'�@f��I�<����q�Q�N�i0	^�,��D�VO�+�;��#��በV�	�p>j�ʽ�d��O=��/v�|,�6%i�]��'JR�����S�e�3��T��{L��ʅ���4g�$Y{UQ��!��-sm�-��s]Ț&G�1[L��2C{:��J�paR�Af�)��r}.������"�,�3ܠd��:Q~q��ϑ�k@u�qC�n:�$c+)�o���pՃ�k�`�����O�����<>{�nWap�@��U\��-�94:_,b��E{?��E�WI��&��z�N��>�g�o/�۝�|�3�}��=-�D��*D��5�m۶���O���;��ߝN�r��^8w�m���<�n.���Cea�g���Iv!����V=�L���Tk�
�KOk�ZU�����5WU`����˼��S*��T�����Y� 8C��]���y9S�>*T�8����CLek�T���u�J����d�����LQm������虈<��-h�*	�-�xҸ��jY>�m�'P�2���^�̽Ʃ�ƒ�Ae쉰:r�q�O�^}2�,�	}!Kj������b/�|��`b|j~��D':�k��%����>��:HRMi��EVV�2&�rӺ�jͧ2|bU#�0�Q�r�I��Q����3�>������ٙ���3� .�V&������Ʈj��1�:k:	�3�0݌�=Cs�́���3�TTi��7�PUQ���'P��$���t�C�j��"�� �Ӏj#���#���$� ���Iα���B�~�h����2 �GwTV3��t?�D��V�����?353txϞ/�t�MGq��#�G�"�k\�>��G~��ǎ��V����S�ס3;�d�ei���H�B��2&)?��;��0����$�ė1�F!�U�y|�%����6�ϡ�r&3�]�N��V�U�9�J���)*s�+rB��@� ���6��q9�c(�4��{��v}S�'���n�ſ}�+�y�����w$:�]�W��K�0σ��@�C��w�Ep��8���Zeɓ�7��ZY����e�c�+��7$p�>����f.o�;�(�2�1���^�FRo*��/��H�=	�`J�]�B���tn+�ψ��8�U��������Q�V�;�~@l8���#�?qh�G�����X�"T/g�N�\��WE��6�*��:��\�<�R�>.`ަ����h���t�~������&W��&7>P}*Y�VE
���"�;�iqg�V�'!g����=�0פL�q�G�N|N�b�q��m�&�����=�V����@i�4����f���fK?N�TÔ����fff�>����?p3Ξ�軔 �H�����_�ō���u�%�R�T���P׊z���
�{Ue%K���#�j�7U�FZ�_vK��'T�Uk��T�|��l���.�W�*�i2��y�p��.��k�0>6��d�W@M3(C��X�d���E�8�!�t�>ʰ�8>�݋�tM+�)�t]<:O_�W��:6����K�:)����
�x,����6r��1���]���>ȉj�"�x^���g��t\��*#�ʒ��ڲ�Ǘ\�wx������9�ٜ��en'iF�ᡰnځ<�fL��\'K,B�x�aA����V�D���Tq ���P1jW���W9V�}�U��W�\�H�R��珯Ν����'n�~��w�ɢ�C59V�^�~�><��q��ql�
[���u��8�)��bG#��P%��3���mh���!1� �k���ҩ��N�8Ҳ�{�����%��ã��x
����^:Z��/�8�hTg��]p���^Y
ՁaC|����q<e� ��Tl�C��I�N˩�m�YI;:1��I�2���Lz�&��I	>�Q�.�Ms��J����i�-^X�םrG����J�"�kT[�l�~�?y�����=�B�Oʴ�8�T�r1�{)������tI!PL���Gw&) 3WEL����lT�Fq�K��Tf*p=��:�����
�����Y��(M��� ���q+9�R	U�fOg��e�ʧ�˒��P��N;��B
�N��r���i�UOg�r�a:a_�2�xF�׭���3��Lu���A�g��a#u�<�8I�v����ico����pdų����\P_q"��,�o6_�8��3^��nT��9B�c��(t��d��'�Ş�٘�,�p� ���=x�J�A�:G������w\t��_�p�����B��Eg?�����5����B?_Q�j��T\��Y[������\���x�)� �X�l���f����b�T%�p�F���� �:��)�]ϝ��#�\P�e�?P2*��JUj;[��7g�g��D!���/	,����x�\2��n����TZ	�>*��XYh)�����u���֧��\�;4�̿�r�mW� �/=����	t���B����󭹋v���<~�V|��J�"�kT�?����z��N�}c@�(r)�[������^´�)}�.hz�S�c��9]Wa��*CTl�-��F�N<�'6D��T�:��/r��MxæV�H�VI��Y���K��_U٘�W�=z�LA.e��(��$j�K��n�����C���
�)Uv�@/��-��r9*ק�	dJ}����rG��nr��*nUe�����ǝ�r6Ǟ�k�w6���k<ި_�k%����ޛIv]gb�޷�R[WWU�Ս�@c_��"rdR�u����1͉�-O(����p�
GL���P12eQ�D�"�QC����R @ M�XzA�[mY�����=�ܛ���$5$��x]Ȫ̗/_��~���}����)���D����b=�5��"�g��"�&ܘ����`	9�|��M�Z�dmx�a#{D#8�I�[I������֛΍���->���}��~�$��V�s�'�swu����l�6OgӾ���D��ޱ6I�9yY#��,���
�h0h����H�TV���5�DA�!�� �>J��(���uG���x��Y�Ƿ�e2%1�}�<�s8�(P�i3
t�1�+X�Z�F�|V��G)Ӊ�����i��9���l������k���s����;N��� _�aA�ʾ멓g����B�j.�G� �Q�5_�ԧj�~쑟o4�~F�j��R���뱎1�sBq`a��9{�!�R�l�����D8p����}>ft�4	����c;�-����}!�La�\���J�*�,f��dq�0d�Z�gy䓛"�1� �b�Ѐ�K�`������BR�JSV쀫��^���e$Yr��*���L�o�:}���T�JK��y&_��#۞��������W`�/�~ڌR�A�ޗ��Yk�>�	�|D�<�7Ŀ1˅@,�6�'%��²�>��
d�'�Ȉ��`)�X��S �`K�+�c��׿��z��љ��wd��{�x�foa_(Ŕ/�ȓ�+�W�$��M��
๊����mH�ڒM�����5�����Yj~�0a�Ou�Y�|�A���{����P;��S��,���nڋ��q����pq�'�:�fat�!/ni5%)i�ߏ�.����8_Btq���$��
�=��<� ��XY�+���Tz���3���g��ܡC��t�-��Y�2~h� ��2��@I�Ǿ���?{�7�i�ŃE�6\Nva�WK����ҕ�]/3�͛T��xTZ��}� Ag*�Q�k�Ir�����`���~��`Ǭ�[�Ep�M�o�C%�I(C�i������\E������$�ýiI�A#Q�[���/[�2
�!�0�$�f��D
�K`hOs�/vp']�����i�Z�f����4�[Zn8�v<F��N����ܴ�������S�����ߋ����o^��S��m�	�
�YF��L2;��9-��	KF�lۀU�E����+E2͂J�ݓ�m�*�x�+�^9�ځ�����O<�^����T�V��O��[�"68��X�����p�!9��H����<��\B@e{2R�	!��BR{������� �:~��u&�J{�ږ\N<�=��az�zwq:b�]Ӝ�)4[=3I����
̹�P�1 ;@mi�r����D�Z���,HMa A�����r���$���u@����v�C�^���z�9��Q(��%@,��k,�}���������;�P��<y�xT~I�y����;t���yd�J`Iϖ`Y��5��֜`���~?����HU�u[=���q���f��P�v�3�B�3 ����9��J��"H�u3�7Lm���j,C�ya �h5��Q��=Δa%��)��#��D���S�0�^"�8�y9�����?����M7�[�oAx��G{������@X���9� ��,h-��]��eZ�+]%tN|\�Ԗ���_V	��\�<��$"�b�h�v^��sg������Sߚ�p�������;)��ZB_�|��˼_:���ϒ���K��Y��BA�k�X���F��50�
&c�&���
����"�s%"'�/�+c7Mb:�����}��>��p�����zM8r��+����
A�eNS���j=�EEv�zB�x:-R��ډ���EC�.�<�q\9u���y�����'>�>�{��e��Q�2ʸ�ⳟ���g��ӿp����'i26R4�[*Y�a�I�����Z魱���2����/M�5*�i&�h���$R�a@�}�&)�F�p�N	�����a�VQԢ�!�UE&�<��X��YŔ��z����A?N��n(}�$��!�%exr�K���64�)`�<��.�\�i�6gDN����HϽx���$��u4�RX���Ju��w�ڸ��} o�0�96��7�`[�\���z5�dX#�*]��5D+@�S�<��(��X·`�}�Sj�� ��Ef�gYۃ#lVq�������ŕ�����ݟw�| ҹ;u�ެu�J$�De���+33�Rp�IO�H�v��c۷
�K�vYb&?����abZ@e�'�"�K�m*�T��B�4�Q�Y�,�9��\�6(�wS��:���`��=���p�����N� 1����@�~��}7�*����Q��0w}���67ڹl���v���ng�W^���?���߿��|��e\}Q�2ʸF�?�����¡?ҏ���S���s��s=I�>�$�������	������<K�6��(��Ä��D��mf�ިͬt*��&���1�i����1eԅ��!v��|ʴ�xq �W�ex��ْ��z(���TVF�Q�P0�V�p�3'�-��l�|���%l�yZ�t$c)94�M|�J��b��S�}kz�]�����b=��79^~��.��^�7�B	��	��^rb�|�I*۳�	K�p�K�b�
�|0��}������������:?4��6��ʲ����x���~��/���>�@(�w{��"A�<��q�1k't�d%��X̮l�)f���D��D*d������@{�����) ���@���%A��fN���G��	��b(z(ݔ-���	P�� �Ę��t��2�]f�71�א`���j=��˅u���{��u��N�5,5E��#���'�e4�28�n�{���=��[�l޼�$�Q�e��e�q��3�<3�����K����룑Hʐ8b
��L�? M�B��� o�bٙ5 %�\S�=j��g���A��sԪC�<�-!Aiff n�W���p8�%;3��1��U�p�r ilk�ң�|pm�5����Q [A��(s��{khG^�b(Ã�ɸ^��ځH1+I���e��f$�����
���^��d�k�S;��z�7G&����;0�7�+$�Ƈ�/�8�� �M���,����<d�f�m,Wkeh9C�� 5X�^ƺ�fvcƎ�)�@�����A��(�6������W^�������=y��^Z8���k��n�YG�YBԗ�O�L��Qo�"�lM��(�HZ�D��͛�V�h�!/��cΝ�����Bt`Q)d�m�E {P%k:�5����l���;�Dv!�ڐ�h�r��jBX�@��4��L,9F�=����I���j:��J���K����k�lk�Z%}I�^��2������|�_ݿ��|���Q�:Q�2ʸ����܇�?h�	�&ش��R��KL>���ɕ�1em�X`�3;�� �ۆ|��C��`�W�j��n�������>�*=*��
�T*>3n����ke���2K���阷��1���!-C�Vn����0#�sf '��u��n;��+����+�M+�D��m���S{���}yt�=�WDư�;�C�������wGYR�9�̤%s;7	�T*=>(���Nk3�kd]K)\�+��BF3�ޕ�*���c����O(>�ӇW�|mi�����ӿ�k�/
�j���P����0E'��n%
���	i�y��b�N�%��O�75k!��ԕ��e��*^�g��<��)�k��%���S���
��\sy� x�ؒ� ��e����������~�G�?z�6'+uIVp[��u[�mv�<Kej�9S�n����c�m�Ae�%@,��k �y�]���g������G�N�K���n q ��d�p�\�����\�˽�2�oXɷbC��cG��v8�z)�L(ػ���R������{DB� 3�E��XX��$bV�yڿ�4�VߐD���2I.�-�3�ZQ��=���j�&gj�-�?����h�(o㢊�<S��OF��xr��;�LF���8���2w]%P�Ȟ%x�)IKkqG�{���ږ��{�,�AC�C��Y�J���I�������8���WN�z����k�ӏ/�����JzD�ɰ4���f2�76�IK��HZb���z��,f��ߒ%)�g�G�k@�؆�}�~�y�Lf�E��5�Y�Y_�$�ځl� :]�Ng.$�駐�%��B�����s=�䭼�:sן�6��g9$��!��������{z������۾�䳿��O���>��>�Qƚ(be\������_}xqi�~3��#t5d 8;������^���R1�Ql�/�:�e�� Sg6KD�� ��K`㸆��W��=uع`�҇���<a�^��Av�t-���Sq��&�A3S����j/3�\����Č��ߙ����3&��ݐ2�X���o2э��#;��a�-��|�]�]��������͹�|�m�R&2�%[:�Gt�eF d7G���Hp��-AEYd'#4���SATڽ^��N����o{j��G�}����;��wLO�3Z�P�\`6O	���da�C��1Wt� �w��D(�Ǭ�9��HH�(�:R1nN2/��0�9KRAan�'&�����y�����#p�M��� �Z��}H�.C����bxH�fjν�͞s)r�Z��\,��顖iqB�T��L�0�O��Ϳ�رc�7��2�X%@,���8�N�٧�����O|(��-���a�����\PTط�q.;�'�]�P�6�:��g��J��n�~�(2�Yփ�zvΆpӞ ����Ơ�]�dD���A� V���B�\�b�Z�.f�94��&Fh �xd-���39I������,��(x��7��$��}]�u8u^�;������u�a�[��nWA�\<�=^>�������� :�f:�$�8���T:���$� *{�8�"nK��"�:��"��:������G��'^����/�|�W���z��~%�
���#eWd�dLdb1s��"��C�_J���$T2Ψo54��V7�Տ�O�M6�$O	���[�����T��@��@�فn��M$8��3Tʸ��^�Dweexx]:Ң���=M��u��������lu��r/������>�|�e�Q� �Q�U�<��?����� U$�`� �H��imO�چv��2p��D�AY� }�D�B�����`�@I�aff$ܸ�
�oaӔ�ȼ�v{�A�O1��f��2X²jU� OC�I���X���i�X�,8�N�Lۜq$}�l�K� �<��+K�����ƛ�~tr�C��ǅ��5~Wn\8�ھNsn�O���$^�� Y�H�R:�DN���/BR��e���*G^�a&R�g��Iyܜz�.���A�4%~�?���x�ؓ<�_��I��~#���#��P�)���a����|2i�#K��9K��E`��3A�=�Ov�T���|2� ��=�5�"���"�ڒ���� �,b�5��v�a�����=҅V�l�?��L㬷\EDq��E���&_��vˬ�4-�V��;����q���Ç�駟~A��O]��2��(be\�q�+_�>��c�>y����q����L"-���r�DЛٕ���g��b�a�Ō�����V8�{ �8��*��SShMV�={"���A�K�G1a�D�!��B/2 �>}|F}��^�	�=A �,�2�������S�� ��3�$]΄a��,xCSt�Љ�H�`�|0��k�S����7�?ځ�(N�~�������qsڃ�����T�%a�B�E��G�#�=|.�^6�>̘��<ִ�R����7�³�j�݃|<�����$���w, ������G��깓O�Js��G���ۀ�Z�	D31�����-�DP[��sC#��ˬ\�YX�IU��0�dι<%IeLBu44�%V4C<��Wk����(�k�x.O�+"c5�5h�c8|,�nl��<����*_W�k��8ֲ�b�p�����%�������s��Z
�9}��o��������C��6|e�(be\��Y�O~����ߵ��pC��+��Q(�1x=d0�H���lg&�	��9,� ؞*��]}���3���n�)`��#�e
�j2���D=�����>3�1��ڸ��3Ⱥ(Y���Iʄ���,gv
Y�IWV P`����DS��'�^�H�]�J$�Vz���b0r�ߎM��ѩ;>|�J���Q#�?>����|�U��Hn���>��l�ͩ�N��m��1�<�,!�FϺѰ���s�T��XV<�������֖3��X�S��b���\���t�쉙�_��~��sՙ��$tn�V��%$���y��˴�0� b�"����i1�`<���U������u���Hp�&L�6D��>eg�j��z��44��pn���"FxF�D��3:���y�  ����gp���{uK ���� t:�V��.=�j�9���:&��?�/=������˿|��hC�/�x�F	�(�*�'ND���3w�~��V�����LG�4���6� :�$�hcO5��2@��,�}M\>$}X��~@�i��I�@g�����jQ��xp���p���+�ž�"�09D����i������@ޞబ��2�
���S�W��|o3���fL=$�H�1�zH��<�@q�d����Ye���7���]�=6��w��-\m���*���=������ad���U�]������x �6�,j�^������n.a� 4"�V�,�c�D`HfA �Y5K�6�d� �M�ֳ@�|�K���ӧ?q��t�!��d���R�DNY;���f3hȰG�rh���z�C����6y{���D +��7�X�kFg)� 0׍U_4 R�GO���0;@|S������1x�
�q��6
ncF2@������a��#�Im֕��GVĝ�rQ|��/P{E�%�W�f������؟\�F��������s������7��9s拝N�����,�2��(be\e�Vjf���̹3��l�L�����kcI�U��E�ANrU�J9�f�����,�.B!kA}�3L$ț&0VװyJ��{�`ۖ &F���7R��p��(h��&~d�&
�]3h'��+��P0@����Ȓ�Ͷ��P��=�qo��Dqt�&OU�n�Zm�M���y�Sb��-�Jcᵻ�+��}I��	�L0+E�oa�mm5ís�}ϯ�A� ��9K�y"�H�H0p�A@O͞$%Tɓ�TO,�ę�?Jl���:Zx**��=�r�ߊ��ٓq=�@��$դ	���
�
�^B�?)*;���R��|�X@�L:�5E�
�q+!Y>�I�z2-��
ĳ�6��6�v�V�լ��B��hC+A��ЀĘd�PF3�5W �} ��yLIv����4ۆ�jO{�~E��� �P�H�+��v$���6���4o0�xߡC���z�����1 �h	߾Q�2ʸ��駟������ǎ}(�2�*ү��������E�Gp�MEb
f��	���k����-�|`=8�� ���&���.+Ȏ,�� v�0�_?R4��!)��}�h�M��g��f�Ųr+��������X'�Ԕ%��l!��%;�P�ӣ��Je�ے[��Hq5�+�G�ѽ�qj����7�\,����ٓ3K�#�^`	T�����q9V��t��8�t��'��"\���>DW�����B���qg��v��h78��c���ӿ�026�<���x�g�ty�h2D����û3�����wt��g��m��9ǋ�a�� p_��I�uQ���6�ubF܀� ��q`��-̷��}�+z#�m��>����K��;��}�
�Rs��E$v���Xz��`Ћ�V��"��I^uN�t�:湨�j���+��V��Hggg�̬�<�� �Q�U�f������/�����+��}����Hb����\��Q��y���ʥ�6N�DS�_
�b�2Ocu���*�{w6nD;��|3z�	8!@�$�Ao�bwb*�H�<�u�G~��P��fE]j��a"���tM��_CfK�y��#�+�_�o��Ϧ6�������̵�k�k/m��֮�{��m)ҥW�g3ʸ�4(�
���N�� M��/�A��+*�b&���o>wB��x�c�����Շ_}�����^�5P�L���ӥ��8e�9��#|�]�G�v�B�ͦ"�m�Hꩢ�u$dWE�:_K�H̪��by�'6���}��@���|���3�
��%�P�ɞ��8j$zV��7�Zp�$	��gRA�3'w�r��Xw�}��V$�9;M�d���n�w���kyꩧ�s����{��zr��O� �Q�U=��ȁ�p����]�Ϛ�K��r/x�ܥL�"��-Z�y�ir��.�H<;����
��j��7�̠�d0(���`�� fg=������������$m4o'=&�8#l3^R��	eS��J[�X=�Jt�cc!��i͒�,�8�8!db���v�T�|ϧ&f?�hu˃� �W{�;����_{����w(f��k�j�-aF���j�������řfI,�o�fYg��!�7��Ӏw�I���2���K��i�2ou�_0��;��h��0�Q�Fc�H;�%p��Z�����8�I[zijbְ2X���i3	�YDu�g�f�mؒY	p�4
��\����qzIͼ�BY�� 4�F�zK�5��u�C���%����x-�^�N?"�8�7���
W��?�Dm��A�{�{�w���ϙŗ���]� ��2���������������:��`3����]f�P��Ág��B���/�#���*M;ɍA����+6-��I��k�mk��8`vF�.��ؒu@��A~)�GA�˩Ya�/$�A}�ʖ��i�����PiP
NnQ�1'u�uC.Ǻ������}�p�?�n|�	�H4_<���8��+(��2$=䠂���m<$Of�O���f�p$�(�����I���K̹�c s˱@-��Sy<*T2
WH�{�M����}��c�����������_1�-�2q�~�$��R�A��ܣv
�8ii���9�h��W���9���aN"ܘ���݄<W�7�G=��v���[C����Gf��DU�Ɩ̈��o�	�Z����!������;�w?XO��x���א����PX���s��>v��(��2J�XFWI<��c���Go_Z\�-�Y$X�2�Y j��A)�:�X��S��9���� ��a���JW����|(���
�Ae)��0;[��w�az2�Hv@�m�	�]�a]Rlr˼W��l��Q�Ětz8�Qϛ�.$��}d���G%73 ۻ�����At������w���m�����r�X�;��ߘ�'u��<�l0jK�d
'�\-�@WQ�D)������ۚ=F�yw~l׭Hr�fy�<�i���

+�}B{��)j͖|�c�ݸE�$Բ��Q�."�?Z��2�,S�Z���RZʹ/М���{��,��259�S,
�S��i>ofc��@Ӝ�}h4{f!Dp��-��30ׁH�?�[G����`�SV����p��W�\�^ �jM� �����}��v��@����e\�Q�2ʸJ�СC[/�����&�[����@T��.� ��=p��D�. j'E�����]_#��8gK�@����'ع�۷0Z��{���+���qԀHA@Q%(k�`A�r(���#c΂��9�0б�찖 +3]Y�}�6u���q�;�-f�-p��}������;�~s��3�����9�Y?��V{l5k j료�{�L�%c;�k��44��.�44�R�5ȶ){L|XL#�&U�v_I���-f�������_9s�_�V��f�lDd+ .�)�'�]��Zò,�b��}�"0羵�4gn)��~�gY�Hz�	�*��c���EN��Ѝ;��`�q��,�R9悐:�>C�z�y�#Ú������z��eP)��'�\�����n�{f@���e�-��e�q���K�t�ٳg�V�!9�hn�Ǭ!J`���!I���4/zԲ 2����*�]�`8!�˓�ܕ��"��Ǣ�*��Ș۶����L�fyf�8�F}���DxHv�����X���(;�0s�%I͂ʹ}Xs2��i+�ì�
k9�U3;qp��M�r��c���㩝�_s�c����w���S	�SF2�8χ$�$`A���0�9��@3��P�&P����^��I����k�@sX+�$`c��dzef�L̟��R�Wz��N��}ׅ��t�>��2�hɇ�0�n�2Cמ4��l�e|�Ƒ��jH��\�Cy%ٷZ�h�gY����)�~.44V��L�G��8�tf=	�5b:݋Y�0D$j��v�L�O�W�@�?�L*aI�B��q��^�Q��
�������Њ5�v�=�_S ^QǱ�7/J�XFWA<������~mqqqk�g�$+,C���؉�9���|�T�uu��b���l��l2<�"��ZE�̴G��-3��;��)�@`���Շ�Y�G�fP�"n��^6$(�����߶��]����A	-Y��#0�#��?v�3S;���c��p��]���C����[��(����:��2�����G�3^�ϖ�*yY�����)N-�t���P	�g������ZfQ�vF�h�n��O	[&]8��'��Bǋ��k՝�#�3?���^��esn�� ����(x��_�O��� �Bc>#M�(�!�{���n�bx�wo`�g@y%�`�އ=�Gpq�|Ί��P�U�Y����1��J��5���r�{΅�~�eeg�f_,nN�S��$���,�m%@,��+<��������������vkJ�{~�u1xmV��K�*�9{h,-S�te[�}� a䲅��͠�R?5��&�l�����G�� �:|�(u`�,�c�d�d�jF�Ky�t餶�3���9����ܻ�z�p%�u�@�4"�jO�z�'뻟�o���&?�-���7���͌�#_;�ſxO�Y��IEsm�ƥ����$Po�P�1O�M�+�i�?��Lxs�G��,$�`"�S�y��Yn�X(C쩬�����䮻~o���?��NT�y���i_�����PF&a�9�0��)b�Yu�G�>\t*�T�5�5R���a'��%�����|s-�T=����*0w6�V���&G��Աȝ�9o2ϱ���cdVg�e�9E���3+i��i��=�pXl%�@�h����Qג�I�x[E	�(�
�/~�/Ɵ��3��nw�b9D�#���M�e]�e��Y�\Q�pmƱ8�H��z��4�^d]�<S��["�0�%�T�'F2�N��ܨ���G;2뤂Z�Z�	k��m?�c��,F�Yqg�Y��Q�LԆKͽ��_�}�:u�'7o��51�n{cܙ�Y�*DJeI</�~M3�ز�Y��	Pk,)3�/�["�$���c��Ɉ�>  ����&*Kf�^��L�v,��h��1{˿\:���������'���~��	�ˀ����kN�*��� d��N��d�����@��Q6���z�e�?$��1�j	"�eJ �nf6��Fpa��B[�F�3�\9;Y�>��1�CAցq�3��C9T5(��`�JѶŕ��^�.��x��t:�Fc��_y-e����e�q�Ǒ�O^w����k�������+>]�J" p�:����#��A�삁�ȼ �6s�ikg�M�I�9�e�z`�L�o�z�dʀ�̬+5�MTX����>e�h��fҩ��1��"�3X�3��f�<���Qߏ ��<�n�g��z|t򞿫m�b�YV����W�����JI��5��0�SL��,� {V)��bψȂY%�^���,�X2��Y�B��<DԵ�EDP����I���-{pĖ�������������ŋ�~,��]W�����ic�R�$�U赌D Z� Rs*�+*+��K��ԓ���[�ڢԐ�_H�عu7�p��
���@�%|�4]�T�Zb�߲�&{�R��N����Ş#�99���	n#�4�O����j��߁+�e���n� ��2��x��'���|�=�Vsg��,w�N>��=G�*���s�H�,ֺ)���M����ixb8�O�:y�2��z-��3!l5�pb���	y�����|M�Rh��^��C�8��p�m�W�U����n��f���[���!ѵ<��j�7>4���/�f\�k8N�����㯽;�4vD��a)�Ӕ��t�Px�QV��W��]l3��L^2` F�LrAg��CQh�*~n(9I�^E\zH-�a�u'�K5�Bk�������W��Е��ݏv�����K�s�,D���LR
ȈE��,1���C�������.R��}f�Mq/v�qri� |C�����캾�:p���S�W�D�G2�>�2�(ڍ�����|�X1X�`�@"��,�W-�y|ee��'N��:J�R7o�(be\����x���_Pi6%@*�g��p ��m�3Q�2(#�]6�#���� �^�f���(Dͺj�=s3�!LM���mu�8��Ek��YG� �[�P:�3��ʟ�
B�>pf;Ѹ��L�S��.�f"
�2P��j���o�֛���䖹��[���]���~�,��r�,�ݴܸ�Gf�e���@��b �#�
qr�(�����yAy�{�2쎣Ҩ��!j�2B-�,�!�E\�/9�l^Cd��5�s���7�7~�_�_�?�������>��A�D�l�<R9Ĭ,I4iE;��^��*#1��T&��4I@�y�����&�&�O>����#ؽ{N]�K&Y�=��tЇ��z�g$��3 �i�A`�6�Q W!'{��E����]���S¥���_z��z�!s]Ae�m��e�q�Ƒ#G������=s��>3��X΂� �x�%B�6���o���˘q�^(,�\�"��E�c:��+�G Q@֏�c	���0P ���@$ 2d.�䋌r3�1�Ϫ"t�A0�.(��2"hg~����`qYE:}����Ie�%p�d �
S������7z����Ӯ�g����߻�j�/�ZbQzO����1��!�����/|�&?l��\	�4"�_/��o�A�)�,X���
ޯx�{�FP�Y5H=�	 i�m��E>�A/��zփ]������4�^` O�`E��{���3�|{I��3�1�/W��5I�8p�=��7���=]�ޗ%�:�.�/��Pq�'��f?(�����{n@]g9��y��shQ~	��3Y4#��'�'Kf��T�ͺf�iر}\�-����Z���:·d,+n���iB�QD���8�WtNYK`+P\)9I�8Č�sY���n��[>��7�t���P��&J�XFWh<�䓛>�Εvk
�HP!���t���D��mղ>e 		��В�)y�֪�1H��K�IE�}s��H�A�Ɉ�*���C��� ���)�g4�L)�)x�ƀ�ȀM0�K�[���E[����͒��I�P�XS��J΀� 1���v��QX�h�eHp�`4�OΜ�M֗�����bv�A�]�G��񡟚5����c�3FB��`=�j��|*��4��Y��lj��9KrgT���k�@f��� I�-wi���w��������]j�M�b�I)s�e��5)���lF>�z鑩�s?w���#rK �8�e��(sH"�j��(@-�1��D"��s�sV5`�>�¾߁Ak�'-F-�J�����em��~����l����~�x�W�Z���ё���0w��`��@Ǖs���n���s��9P�uZM�a�K�t0��I����e^��)��Hh���Xp�6|�U49A�a�!�m8��Z�h�B�i���Іf7��5�����Zr+�9��u�QK]#�!$D�3B"p��zǃ>D皂�� #�DD��p��؃�a bd~�+��r?� �m%@,��+0<|��>�oi��u�^;$�c�2�)�,P`^ �НA�숧�I�� ��B��i��U`j�Fزc��$��74�g���oo�}���a#��	D!2�K�eDj�
LOE0Q�u@���J
Kbv`���|�.̂���,Y%0,~�PQ���IN�:|x�����G�'���l?���-+��8[�����RK�`��0��E�d�<�R�9juR'��JN�S���\�f`
A��jpt�m
�J1\�58X\�0����;���rmɞ���Ą<6rV��%`[,鍔�̕ҞJ�(�c�T3��W�66���+����ZU��oS���bu���~�b��c_SZ\ň-Ơ_U�̚��Ж8Ӻ&��B��{�n{�ғzt9�i%�^�+#G�3�\�o8;>�r%e�n����_�{HڣǓ~(n����҉�У$ѵXۀk�����z�|XY2����o�8��,��
�Sy�j����},E撂��9l����Es���8�>O�3$KM��p@3$e��Zu'_ST7pz����-�c^�Dt�f�(�m���Çx���?��'8_��Q�2ʸ��}a"ힽ��'7��JrH�T(��ɝ�!2%3�D=4ݡ>@�L iD�n����������hY҄�yo-�Ȗ�Y�"zq ���p�@�@�#��PY���Hv�c�{�������f� ��<c�Y���!x�
4{���%���3�5e�X���Z%i놯�����p�ʗ�t�m��FB!��*1.���9Ԟ��\�����T�U8������Z����`�G4��	���V��R���']ez;�(+�cߛ�s�fJ�C�Ϊ�;��<X�^'�� ��(��VLyU9R�A�����"A�u*tѡ�wj@�K�xy��y�?���ϒ��ޗ&{�ϥ^�E�?+.�?�h821�+� 1��_n���?�B�nno�}�w���	}�YW����w��;�g�_^2`����AE����]ѝ�\���o�|%:� ��
زm6�x~�m��Q3�f�Q�4�:�$�v���oz�!�I�8����h�W���,#m-y5G��Y.l4���M� �M��e�QsC����U9�x]��S�A��4Z�����op����k�v����[Y5�I�7�j�k��L%O]��Q�J�+���ѩS���w���������.\YHzb0��A!c}�̀��3�n��zq
yڃ\�������v�̖��V ���7f�8�^>i����>ͥ'��,%�1*�:Ǎ�XS���}J��}Ծ�Wr�[�3_9s"��m�Rsld���Rv���)�����#7�3��M�d�9��L��j���E��� F���:NKlZD����pϽZ���:��w�{"`s"P�j�h=�`�7;�]k�`]�Ϸ�3�u4�`=�����1d���p[
�E��ҫ1�@\���i[��R�k�;������(�LZ�(s��+� U�w��2���ᄁ���3M�߫�Ʒ��ſ��[�"��v��w����?���Ż@����E��1���~�$5S$���Q�]@�M�� �l0���H�� 3<E|��B�y�Ip���̹f��0��
l�&���6$����� ��^+��mFж��L��L�D��� �y6�i������j5lo�~�ĉ��k������� �Q��G�|a����_L��{�k���@�R��̀��IB+��8ʼ0����ݍT1�D�3�ԫ�B���)�00�-W��W����Z�FQ�us�y�.$�$���K�7d���P �?)e����1�~�L�yP�}�R�/����fr0�!mٌp��)c�O:T���9�lC��T����}#5�$�2r��f==�䣌���+��,(\]�� P��G�ޅE��`F)����y/t	`R�����p3�Fۓg�-����"qۋn�s��,�,��Q���'/^�b�:�Z�7g0�w��_�e�+e3��E˹eӺˀ� �]5�o��êe4�Ł-Ē/	��C�G�r��.�B�@����V���H	!c�7��R�~T��CcJ��[zi����<��c\�+ �l�u�����BޛLN�� AI^�(C�I�{�Ej��}dQ?�Ҽ�`��k,����>N����̥�D�X~H`Op&7D�sGv���J�z�_�k���f��·��XFv��(���v��Ŗ'�����[μg������������E^�2��(beؘ���r�����7*Yޞ�=�|1���p:pX^#6F!� �(����!�e]��M�=��B���d�Hb	��,����>�	⨁=IhF�MLP��~&lѭ��Z5�HTc�/��@5sXY����2�IF�M�z&�6���x,��Ă�ҡb� �P��\j@�c@d��^ȵ�cU�FC��le&�2����P&��kj ���!�Y�uV��Ě)[��Ҍ���V�/%Z��3�QLz��OE����-�lۚR����Һ�p��ٖA�;�N�e�6;t�ಾ��Cڏ0Ԙf�e�\o �c��W�V���~\�@�*G^nkŗ��J�9����AYC��AL�OŚ'�|�Sv�V�=UU"�NC�I�bsk9S�3���趟]z��T����~�������f!�^G�a`!w߀)���֧��G:NY_B������"؊�c+<��$DC����\���Y��Tfg�p�D������\{`>�`�S$?d�`1\��)ĵ =�a���첋���P+��w����t:��g�g�?�񏷠�k:J�XF6*I0����^حk��N�CK44�3<����-+��	i����a"J�PV�<����s�(Xl&6�f�t���N���ePr�%8X(�(��6]$"�	�.K|ࠧ`��K������a��2�Q�Ƭ�:V�-;���ݳ0�c�Fk,���({��T�f.�[�s'.@�|�k����0:9
��7���4�����R�[nA.���	���i����̶��@&�pd��`P�hA��G.'�g���(�w�V�eb�M{�Qd��B���V���}�����ZV�vgP1�H=k!{f;܈���x�K����K��pż9X��ax~���.jϹe����� �::'�B�R2}���=x���Յ������E�������~[e�P�u�d>s���������ovK��\x�WtO��$�ԶMp����K� ��taq.���Ce�J�(I��$^l�͋DF�uؼ`���4��IR�^�p0a*^# &俜_җX��~/���?�.��,�M��������y饗v��<e\�Q�2ʰ+I���nz	9N�(1ae>��Maքs�fst��^d|*.�J�No��UOm�̳�Μ�}�o��σ,j��8��+�fϨ�?)�'���X������,�]�������� ���,���؁�r�����
~��J�]�diN=�O���]�7$$=.��\�i����2;['��z\bV6��x�q�}"�پ��|��9��dD{��H� (��	���NXBǳ%`�l	�;7-P_]=]Z�.HC@�Y?�N�U(�%���-f��Ǭ�]�m��QOaf3~�-�P$}P���_���=�X�^�9�~�����4���es�m�X�V�냗�^Y�2F�"u�E�/:�v��d�:���_�w\��0H����+��}����uI�����{ea|�BZ�苜&1e͔π���.�K9�Mx�l� e]�'ѱ��u@�}��*?Df'3�����-?т~��5�ɀ�m0���/d�DGD)2�]�bџ��A��;�e��J����ĦM�*�z���)*�'%@,�'��u��������!��o�]����3y�����i�$�}�{}��!8�+6BU���=n�i�V;���B|��a�G��An�9�t	x��<�`9�@�$�0S�}���rM���12S����v.�?�O�C��C�G�
�)�� t�X�E� ��̘�	��
ЭbaνrN�r� �&��f ��@�>��GY�^�g������� ̑M��bC~
�������U�(;1�5��@��EyB6�V8�$�=����R�"�?$��<8�20�~��g15�k�ك�}�%/K݊� � Eo� �W��.�z>x��H�g<��p}^]o����}���(�'�/Y0~��e�w�
팃L#T��Cgw�+�����k�}�̞�>��T�W=�ɾ_���>��nO�,/��&&�׀�0l����ŋ�]�6���E�H�y�������rm��6$�r�̃����B�13ɪHs�`q9��w)��JJ&�0{�a ��n����!4�MQ��%<1 �P�!t�
��m�y�(�]��+Jܬm5p�pE�,�o��'y.�
� ��cŁ�(��jGq�����{ꩧ<�q�2����X���$������ssIG��$�Ʊ4�Vժ�Yi�ߗf]���y�Q��⋗܀4�F{�G|��-��k����2˺2�=int�o���D3fg�l�00P�:h��QO��ܻ}�w�q���ۆ%���s�$�̈́i���~�^��n����aɳ�}Q�uzˈM�� ��}��H����n@bT��;�t2X^l��ehΥ��S���J#�'���,��|Ν� 74n����U"0/@k~	��/A��C�j:}�K�ٞ,I٤�?
J&�8׀�P
�X ��+�0(H�E���FA�4\U�u��$ҷ�b��eٴ�];��D	+�C�Z!l"�e�T'��ź��G��#vY��eC�m"u�t�i����5�"�^��ᾶ�֗��|`��+��s\�~\��F�s�,����I�|���ǡ�ʊ�_�{!~�oaP����'�K���8��Z��xd��n���1	eSs��kQS��j��������1M�������m21�gwK S��l��M�>�=�A����
�%d��'����t��E��~DW�.��]9�e�}�,���^�Wo4�P�5%@,�G��ǏW�;6�����s�ر�.�����6���	sS�#�3�>�ݑ�=޸r�R�����ޖm[���:A�y��6�M��<"���'07�5U`nD>:|oH�Z`cMq��pT.DԭEe:�E<T�q۴V�(�y:YZ��+�w�����@���-3��Y�bťd�ʈ�Iec� �\(.3P;��7�@��:�c�
�H��		7ȣ���d����*j{"�/(t��� T'��P��@��B��P�F݃͘�F+�0�����f���`iq����=�*;�� �錥^ܲn�	�m�pn#L��2��ySF(�A�d֖h/-����̨��"�U���g�����V��. y>��z��7e����!�g��npy�hۂ�C �W� �چb���r�C����]aٴ�� 9`ˠ^�[��>T*�����5;�3�UB�}s���K�ռ Ok��{B<��,��	��~�����_m,��+嗢5�ǱE"1S$~7����ߜ��=�aŇn;��%�"
���h��ըL����(�Ct%�/b���a�lN�jB�Ӧ�8N�$�ې��$�"8t�K��X�.�[ƕ��sE�u��nb3��v���=z����_x����ӏ ������f�g>���:y��'N�|�ŋwu۝Q����t�8��J�Τ�eV*zzzZ��_�cyf*�����s�3����]v�rLK� �U8�0s�s,dZ/3-��q�=6����Q��՚�����e`�V2s�LA�[��S�Y���G���a����e�\>*'�3���Ҝ^=�b�!Q��	ܜ�Qz��"��!��h�!O%�]I˼?�m�0�˱fX�Q+���L4	Q# �{=Xn6��,�¨f>7������Y:�">a��J�����5��H Ìh�X��G��C��z�D�Pv�+��~buv�7६�+,^ p�`p��Rq+���s�V�������[+s�A\��O&O�Vm�$�X������f`��²�q2�ij�P�[77����������B������w�۟�n�⩿o�9�]��-��M�ؗi��r� ����:+�o�fR����<ѽ�1��rnGɰ��?WA����mU�<�#��,� ���X66�m���Lm :}C�����]�"N �GW��p�H�z�n��ҍ ���<j�^�2��(b��s�>�'r۷���:t�W��l�ݞ07�u�G!�İF���Ɠ�AVo<>{ڢ�h�ץ7su%��;�+����;�ʇp��P������F)��|Lt��=JQ�p��n��ì@�{=��+�i�&ۊ	+BXgA3��c�	�2N�����D;VdP z�u[��%ZA\�#�R��h|f0co"�HX)���;1�>��w�SwT�*�#{i	�� �ת �Й���͸� i? ����2s�k�e���BINĊ�.�N�lÓdZ|�{29B��ɪ�����9�*;��
ָlgt��v烴��^�
����X�����%��/�.�6��2�ו��_ b�z��ضZ��%����:�õ���a0���^��tγ {�:ɕ��y�mܧ��tMb;���HW�?�N�t��E{���|�Y�;�;���?�ZY��7OT��S,
^��e��u�<Lݶ�f`l�a�F)�=$pU�:�=o%Ky^3�U�6���+(6n^���B�X������qQ��I�`��D�	U8:0���D����Å������ ^�Q�2�G>������_���~&��7#;��W��2��f�&$�j��B�'����j�J~������ޯ��:ِ�ʍn��\��䔕X)����z�f&_	��qƃVT%��"�S'�E�n.������<"p�}2� 纼A��#�h[��40��/�mB���(�9���-1S�P��gNعdr/?���d&6��|�@{�c�����,)��nރ�t3[�aÆ	bA�i�1����,�I�&(Ӂ�Q�u�p�������,I�����B}��H���2x끡�w.�Q BN���Ѓ̕.H
�Z��}�]�J�#c_Cú�E�yt�dq��#3�/}�=��:��|�;3�f���^^/�Nk��k���.]���_p=��',�� V�ڹh��'��}�Cb�R�@�{�l�C���K���fg���.�y������<i�ZQ>\�ťr�_�j	S���ԇ�j(�!�y�i��)�ʓ+e-;�$02�æ-!LN4Z]y�o ��$���E�X��Ow��X�Y���z��>e�9�L�-��[�֞��~���|�+�>��1�qMF	˸$^}�ч�����c_�gN�~���Is�\r��@� 	��/; `f��3�����YD7���zt�ɭ�(z�tk������x���(:q��T��t�`_�0��dlb��K������ϴ�h��	��!������a=�y̗���pqP��r�y�~���'9 A.��A�bK�v�!��S���QF7Var��'ڰ�Ёn7%-��3`�t��87��'�f��ہP�P��uL�W�R��C��(�b[P��m���@ŀ�@t�����Eu��ɶ\̀�r�����n$U� e�+�so���l��0�&��[��0?ǝW����f��V��ǡӱ�X3����zO��/�H�W�^h�]�԰G�-��F ���M���j�Z&�]�C����ځ��R�s5��ҵ'�ja�^�Px�ݬ�����o����8���������^�;w<�ߦ�s�� H�#$�+���G�evZ)�4r��
��A�'��Yf=T�ʤ%N��U�İiS۷��܅�:(p=b�A�w��u{� {�w� �Z�I���W�q�Ҷ��<�t�YDs/�9y��=����#��P�5%@,cU �3������#?w��{��w\a� �W��9�^�g�Xz�>"��ִgA���
��@��Zp]e`s7��M��3Sd߹�B�C`�����Kj��8��3��@4`+�>:�=��J����Ce��q�O�ҁ4�\v�X�ѰV����j�4�p ]/!*�+<�eF=������b��8��2���i�1+��hrv���r ��:;~�N�x&�*�c����}0{�6r]�"&0�Y
���HY�B������lw��V�Ā#	�Zj�g =��c���V�^B�`{�N�l/'xC��C�-_Z��H;t�h�Լ�45���V��+��vvӹ�?�-k��n'����Xn� ��r��8��+�a��b�h�a^Z/Ӿ&����`��y�'��U��;`^X��/Sʦ��$P��"H�ɲ� j%��~�������ʓB��+����w?����^~�=�>��;��<W�t=	��M�r�.��4�z- 9Q�~E�צ��9&�KjE�{���D��Zݶ����`�ĕ�?sL6ʞ��22�	��V�'�Et���dq���>.�ժ���[̈́J�x�F	���?��O]������xј�3����؀�~�e�*fj�}e�`�
f�R�y�ْ����H�nn��r�?ohnl1a%��a	�I�a�Պ�� N��"���eya'��37b���u���Y�eYr{��o̡*+kꪮnv��-p%�2l؄!�� �?���kX��l�À���$�̖�Iu�!��2�U�5eU���;�io��q�>����efUw����n���=��'���+�7��*ak{�%[�J�~j�ĩ��(g�<>��[�(4@\:\�Z0��C�=��D��[�_O���(MM���ҚZ��Ƨ�KEJ׉A���lA�ɽ�o���L_�at�����]K{���o�	������q�O��Hk�� �lC����I�&>w-M�"�UL�:�I\T���4��1�z�l�1zX�s�=�U{"_��=�*����?��z�h��m�gJ.�-�jϨ�W���y��v-۷0�:z�,� � n0�h7o����v'u�����@�k��Cv�w}�ó����dɜ��ݬܷ��4������_�.;���j�2:�W�L��KϢTS�c��s������Oy����qv�Ͼo������f��O�L��8G+�;6kF�<n��~�����Q4Hvi�U��--9ޑfЬL	����^�?�-�����#8C�hج�#���<���9�َE�lD��|w�m��)�%9�Y���lt�������֙��#��l�u،+;6 q3�����_����������#�S�L���y8�8E/���rs~�h��U�����\G�Υvj�?"����e|Ձ~�t�:�Tu\�(�2lW�X[7}�Q����v���nW0�8��]��K1Z+)fz�E���7r�0��8U�U=��-nQ"��HS�9��b�^,^�)��P?f���^Û{/ë�_�P)79d#Hܵ����r�&�����t
�n� ������ϡXb�9��Wc��M�:�a^��8��w��7^�ۯ� )�lۂ��Xt���(�Vۥ��ßr����EҺ��=J�{�A1�_���p=���qn�?�9�_��H�����|�^����E9��t�C)l�G��u��h83�~����f�Fǯ�s 1���������;�ATg�[�����y
�E�*9;��'��;0��9'�L�d�aDiet�c* ��KxI��������#������d����zc���AՂ~ۣ��@^�&q��w�|1K�lw�H��	#��B�Z���G����jO� l�s=6 q3h��������o�޿���,�+1&L0��&vg� ��Âh�[T��T�7�rHFS8�+88�C���(!��8o�S�\ ���A�#j*FQC��MFȋ	�����{D{�4L�����q��4�t�A#��lhj1e�+�}1���W�|D����eʶ�����R�R���(�5\�lIF� (���H��]]�wH�n��Ib��a$�ˋ1�P�Xo�f,�/p�;��z	(ÁU�t�pO3�q����Ç3��<����U��4�a��ʭ?��p{^{��z���P��;'�;�N&Aku>��i�gݷu�h-H�)壍�W�Y��o���$B������{�(FZC}k����}��[��O�0����٣�����������\޶�"��.E�C�xb[<쪂�_�#�(M3;^��A�]�@�QE��)-���c_�B��=cQ�l�X��ۻ��'%|��ґ{�T�RwP����Ԗ�F��^h;qm�έ�L�����9�!�Y������ߧ��'/���;��6�ʍ@��!��������������4���z��x����Z����{����N'#�sp?���p��	8Ŋ�U�c���@[�Rq3�^*5�|CC���L/J}�X�&4r�?U�<p�Qi��m�u�s�p�uc�
EH���Tp$�,��?���(�r���|u�@+�r�=�����w����z�FR�ca\,���e9ly�,� ����Ut-�	�rb�Gaz�2Y�W ��~�]�|��|���-P*�MPn�C!���}���K��^�ۯ]�^��fI�4�%i0�L�@�����2� ;E�Z�TF�D����tl�	~����-qX�`���{�t�ȸ�m���N'��
��;0j��?���~��߻;?�E�ꗜ�+�1����=G�����+��
N��Ha{���t�����T���"�{�� p�R��[;p�s��H�uM����r�|����c���4%��fˠ�����x�8��nB7�y���FG��=z��6 �
�@�x�����w��_���y4ʶ�jԲ��n>�W^܅��lM��M�j��V�:8ڂځ����?�f!'/tgg&�[ԡ�����s*�h4��Ru�fϚ3kO?CL")}����(|(��#҇׶�b�6���ՙ�}D/]c�z�Y�����`��C�4���W���ϡ�!%���Bt��h�<C%�:.��&��x�(U�	u0��T���G|<��$�=����6�N�X��ȯM���-ػ�7^هO?��]JK] ��n��2����us e��Gn�ZP�yQ4��IK�G?�����Q�X�I�:@s1���421�ة@�<�������/깠��>���8\�E�m�����"lw����	z`�_�D:��a�F<��`���W'���7����U[/D��Ųp甀��f+�ǝ
��]:g�8��Ĺ��{���Q�^�BBD�Kꔄ��`�F$�mn\�!� %����{��u�L�	]�w;�C�&��r��?��H�9ԧE��뒮,HG;_�x���w��U݇͸rc7���Fw����Pʲ,"#�Ԑ��c�ى{���^C	�4&��ؚ�w�\A�S�I��AU8�9�	���)d���5�E�z�Ɓ��E�/%�6���N4�$pd�!�per�m����D���U��K�$��Ǟ��該�kZ�=���K�˦U�*��"�B��>^_��`�Q^BDy������E雜
Hpeu��TQ,f_�������dC��7�N�a�mع9����P��Z ?�`4�8`��:��t��jܺ� �^�9�P��\�����w?+��v\p�i.~�y��y�4�s"@0�/����3\4*N�.�r���s��?Mv�`�8�E�=�k����)Jn��;x�٨X�*X�e��T��jX�Uk9�$� ډ^����7�߉����]v�U�t<_�7:E�5�C�>���0d��� ���eqD?6������o~��'�}��?��_��
6�J�@�8::���%ۘ	(���Ho�)�<�����a����HI0�Z�8ӝA]8@P�9�r�C����q�{��1L/�Oj�]u�y 0L9���I���@.M��"l�0��xQ*<���5y��bUם��U�/��Vr-�|�ǐ��`wx|+�n��]���Y��)ih�W(���&��r~dXF�.�P��;������:~�Q�Ns4�ø���TW/�X��Q��,�b̷Ӎ���"�*6
����{�F �z�5`�'<VR�+ES�|\�g笫-:y2D�s��
S����u���K�0��`A�b��Il�yUn�s4~�?�����w�������M]����H��qT�g��}��f ��G%��"P)�`�	>G�I=�EjGj{-��Zõ�^����Ud~pY4m?�E�u�{��JU��M�D���B��1j��	GQ��~�뺺��w�}zz�=��#،+56 �k>܃�������/��~�%Gޥ�)��F��k� ����Tj����R,�4���Tu�0�مݽkPZn����IC�>���	��(�U��\2$
(vW�b[�Ɔ�i'�T��lդ��f0��`J�l���tBۤ��D�|C�"�zE���#�tפ�ß��_�*O��҉B3@m���={��.��������J/+�����"��M ��D*�D1�\�G�<��jyJQC�EG���������?\=m�l`c�A+���	\}كK��Op��m�1�I�?�yS�GQ�])�j�	C������Iy]�[�w�R��	�_���W�|����������q�fK|��8��N�����噁��͋#�n}X���4�_�Wc �t ���=[q���I��Ɛ�K.��N'�^b�S
��so?�i[�I:��( �s-��IYU��>�������� �+66 �k>�}���Ï�����M458���?$�X	�n��z�`P�+c���7��&�
�h������w}F�"T؂JW��ưA����t2��#�B;(ji�!c�Izd�zm��y5��{��ļ���4��-K�M�[Ņ����(�%�L ��
��3��$���.�ӻ�ϱok�Z��7��]�*/_-/���t̳��O�Nn��X�k�ۧsԮ�̤�8^W�t��9�cr�@��)2^���#d�"�h5\,�ц(Ԩ�#'���9oJD[|0��u4�=��^p~�X�-DT�v�J������uy^�������2�K.'�MA����h_����W�{)�W ;�wǒ���C�cB.tb�윘�R{������k���&n�Sxl���F����֕u��*�kC�2�L&�F�id�ƍ��j�Z����X���(r���{�!�~����Ѿ�0�L�������:[m�v �CW3WT|VhV2'mW<�R�L6�k.�ʒbFJw!�m��a��=�����o���{߰������f\���_�X,�w�\��"��9!;2
,:�AU��K���!�թb,��`��5�߻N�4�������6|z��wC51V���.zhZ���Z���ǿ�������lz�r.	W�֖*vc��s>����#��y�$�m9e�8 +L��D���?1��:��Oq����0��X�[���-I�x�&�k��i�tb�$KE.�ʩw�BƶE��ME��N�u�PAj��Ů�-�j��ӰqHQ=o|ّ�g�x�[�y)�ˀןj���O�~88"�BZ��[�J��w��1E�r����ڧ�J��_��Ͼg����.��wQ�J��D��~Ϋ���=��t�6��~��DEg�ލ��P�Q�˞�*J+��M�˚�uα��������/����z���J���%�&�_MN'�X�b7�b�E+�FE���zP�������>�"��WK��	��f�=���Q>r�,9�"��Ά
m�����p��H#)˺�h�]g+�*U2;;{��_�����W��}��͸2c����޽�g��JY���b����BbR�G�C-�EQQj4�^��H`
���t�ְ��*P 6b �r
hg0b���Ձ�_hg����K>�(`�Gغ��Cl�(�Z���V�-���ld��R>:f����=�zn}�<J�i��	�SJ�'�8�k�b�����1]�P�ߗ�_w4��I�����|�H@���`֯��8d�p��$0�,D�E�"h!`1��fAo �U��g�R9��H��"k�,�岗�a��2�zr��� sx�>:�����wpu=Z��WD��"����Üa����x���#�����/�����;I��H� ��8؇���4nu**i���'�m��%�A�l�ҍѦ*�{>u�@_���6h�H� Ul�)��C�2���m��&snblTl32��(~��zq��L��s�H�����ᨡ�.p�(0�����b�`R�g�.V2��|;L�|D�kו�~��M��Q����2xpj��%n��A�q�-�?trCGFl,�?�KO���[l.�����ŷBK�Q��|��O�ppp����x�� ~��iUm>��j�T9��4�H��~U��C�9u@ �P�Q�ӡ�@�"I֦a�3r�LĆ�$��{5Dmu��ru�B�bg�tk��oӂC)N���G���X�ʉ�m"���/fO99���-3�+��l�\�z���"�qӦ1 �P����p���]�#+��)QA��Qaes�g��ک���n�4��^Wm쁠�>j��R�F`\��>ȏ�U�K�/#�v�h!/ק8��������eR�?������U���`��߻�1�]�^#���Bg趤�����*2��kw?}�o����U*��B��P�!|Hސ1r��z~-�,������H�Dq��2��d)oʼ7��T�\B����2���l��%��ӴX��s���G��-��9Du��S8�b<g7��N��(�cSC�^��e���-��J�Q���sᶍ�6NYс�^vF�6*8���hwE�&T��phS�T��4������S�>�͸2c��������lv�����L���PE�0($���)���췞�@��D���nqQrn�H!�H[�d�Vę�z�R�S���N�yf���Q��6���C<^�/(t��{�q���:�] ��g�y6)�� �	ʳ�F���m��%%P�� 
���yc��
nܾ1D��ut<�y�����x\�I@�����YIs�\��0��,G�T�>mlZ��(̲:�O�$��L�oFB�a�GHH���eB������]w����:�!�����E�]����%�yLU�E@i���6��h�r��E<�^��Ǔ��*��W�ӁOW��S}�L����ʝwb�և;����8�Bl�E�V�ڝ�O�a�s���9���E�Xq6=?���`QԲ"0�:�1�L�.K^��s@Яl�8_
*,�s�`Q䰘%P5$R�^H�A�|\���hʍ�5�D�pT�K��LH� u��T���A%D�*�tv�Sr/J����u�p��p��dY.����،+56 ��=��G'�E�/�%�����*�
*���sj�nJ��3$-)R��a�äv��"�/�FH�o�+X.��M�q�pY����s�۴��T�@���!F~v|��b&��qy-���	 J�����w�L@�vYR�	�/V��c�Y�(K�N�bJ��ga'J���s
�ķB}4����H?�U�3~p��$ZZEh��Z���4���)?ق�
fZt��'Z��p�D}AZ���5]�� �ȓjP�-�p�D G�đ�s��@߳p�[�0B��"�?)��n�ֽ�>�z�w��/}��`�,�!�w�Xd���F�Vs�r���wJ���i�tc��N�@��񚧦�}��g�ﳡJ-��Э��i�㧍�t�tA��J�Ym��m%��1[B�׵Ϝ�N*���' �YY嶓:kx��:$�Y�z��q�E%ܸ��dZC��1�}�]�9����!������QD�����b@��n����J~h3�}l ��x���;z�8�I�R�+�' �JV2nX����XQG ��qTAS�Pg�(b5���&��G9�\Ɖ�6k�IĪg� ���p��^*Y�mDRA^!G����C����c5 y�򺫺 ��!	L�}3TP3�r���AeD����h*.��-U�~����zب�Ds�&�*����XP����2����K�iN�� ��'��Tx��X��T;�R�)��r��"��p��Om��EQD��m��>���0��:詿z���q��]�����ǥ�/�~QE�X�P�����ߺut�yQ��&����B�%Ix�!�ץI#pA�'�a��R�D=�����;�#��e^�՛��hԶ����Y�FR�uu�T��1���g*���k�sF�r�S��g��avjܫ�i��\qt�Z�����0�;�^�p6���/�p��GT�FD��MO�T���
�#�C�f��֤�l��#���SU�{��ǻ��H�|n�6��� ~�G�L���t<Z�2�~Gu�����Q��>'K�̫��D_�l@2�L��'1���~1�BÄ����l�VuИ#�(�dU��id, A^ ����^M?�sN��?=�3��=&�3)XiE�q��ư��. Tp)"V��̍���t`��Z[�z�I��]j����/���/��("q�r�{(	�j�ڇ��뉟��Hz$�	�	����\�����D�M� �JW���r���sF;��}�`�w.9�uR�<�G�¨��x��E�;���4�
_S�a�V��.���}���o{A*X�}��N��p�b�'R5��0a�|�ِ�s������2�be�:��A���9p��Ӱ\9֥�e�������S�D��g�oq��!<g(�����$�ɤ����ys؊�!��PFF��������ZXX��-r���Y�vx#���?�|mP ����-ؙྖ���$+Iс�}��%)�F�Ȉ��75�V8��a�v����e����m�XDUU�_������_K،+16 �k6,[����������n]��ſ𫿴���-j8:����!4ȞN�0�s9�wk:%���
YT�R+�&j ���o~v�*tv��HE�ȹ���]�s���$�P��}� 
�`E3����f��{W�} $�LSL9I�]=#�]J�{�uC��t��Pl�Z�S�
��6"�,FP���"(��wh�8J s�#]#��ۂ)6�ࣇ��2y�@��"��(� �Z��LO��3�K�=7	(��}�ӧ�q���y�DWi�R���%E��A�� �R{����!��N��hĎ)~"jci=�(}��lVa@;�3�r5�% �����6�w���>M~1+�i+8x�0^� ڹ�<��=d@�LQ�;^��U<�S�/��= ���i��ȝD�L���N]ʰ;G\����)��(̎�<[����%6D�q@N�}�l��GM(��\5tG8w5J�ݨܳ0'wǚ�T�w��5�Ɇ�U˂ ������t�c��Qy;��u!:��LMӳŅs|��i�M75���A!�a�� �⚨ ���A,;������%eu1��,��������f�6 �D�3�aDI�?���=��ma
p���G�&'PW�
��w�� ud�H�Y�a�WX#���kM�Q��eQ��G�j*�:��z�yE�<ϑ��}:?ۇ��Rcs1��>�)��f������ݗu�wT�n�f'i��߹u��V>ޅ�e���-9��ڭk�Wn�45�a��.@�IҦh�S�`*q6�5;���6	, �8����{��8�Lq�|�8Eh`��î�e(���-��	{��4���K=L}$��h�Ac��a�	�(�V"8�QP�Z�C�|�&L�0������/:�^��}Be��i=p���q��e�TH6O(fI�!NT���AJ�J����`p0� Єƽ���]���<A�%�>����:�<�x6�壈�c.���!5 �u�'�~��H�{��M�J I�R��_t#�R���#�"q$�2܇�:�[�HK�)��լ��D�	�Դ�
�ڛ.������>�w�N��ze��НU��Z���Ӎ|iVD��%��g�	~����g2��D�OW�Vn�ȟc:� �?W����4�=Ȳ�H{���r(����?b�\7�bэ�h�NS���[DΡ�s�rȁ;C�y`�p��yY���vL�U�����x{�)r�N�;��^��ĸ�UG^]1K�
g�͍�*���=����>�<�͸2c��{���Σ;�Ï��O~�ů�����y���]�ϧ��qY,��陳��`u�����d/�o�[�����q��y��)�˙�O̗%���*(�;ԋ��t�lsC�h��:;;�����*���r_tL���@�e�\ð�^�B�����)r "����:��n"�@ZYi��g��;�H�*�S��sf�T;��dJ��>*� Sc�StF��LN5O)�����a!x�n
uZ�O�g���N�?���*�����= �y�}&���|���=�'���������"�K��)���'�?x��5qN�<
%�{L���GGUniC����~�ם#�vmX�r��Y!!��Q�������a�,=�X��SĖ��ܾ��3JY�Qf���k�� np�)�FVrF���Ϣ8f��WyY)�2�1�򷽶,���`�a��i6M���I@P8� QĩKȢ$i{{;������jk�_����.�B<Ĳnmc(&�#�C�t��5�&m!a~z|r�Q}2���͕�xE�{x�?��o�����]��o8`7��I*0�$�mI���7Y8�u��
4,�9NF��f1E�����r� `��{hx�v�@)	4�˲�I�R%1F�8"���1D�g�Q>�����0�z����b�Шi_��CNaEsg蚞�ci�J`�}Q>z��O,�9�pU���޾�DzC��q3�q����(��#�w���E��#�
�
���u,��Y��W6��텑��z�����y�cݾ�z覅$���&֪O�3��A�P�����ծH��at�X����/J����ۡTM�����;�8
��s��j���ߠ��;8p���g�@p&A)��׾	#ľ�y��4�(�y�j|0�VB�����F��K��G*�bj�j�v������((ɉ��R�d��5�V\��XC�ݮo�I\j�I�I�3g*$ |kڷ���K�4�.)��i�G�
��eX6�����fg�N��ǟ�f\���Wt�������7�����h�8�X����h˧��px�<|���9۟���5�a���99s�G:cS���O&EM�9`�@bT.�7��ҁ�&C@��/�� ORj۔�	$0��S�'�A���cD�q�/�4��'��|'��@��(��60������_ۄ���I�ځMM� .x��ZyI���t�aM��с���r�W��q�6u��f�E`|d�N�-���v߭��V`V'a�Z��:��pY��� 	^��;�< '�']�E����Fe���Y���z�A����lh����e0Uw\��[[R�Y����@py��$m�<��sIEl�w�Ttb|�[��^ n�h�Cȅ 1tH ��}x^T�`�n%rʅ�a��n����jW�ܫt�8�G�+F�B_y5ܷP��v��^1*4tm+�_rHũ�홹�Ϯ�Cc��R��9�H�Q�c�H/)��+���~C�[�(O`{��е�����Sw��]F%���u
30��,��%��Jq��r�?;^��M%��xE���\�{�o�lM'I4�����8::�{�C2��b����c8>����=w�A��D�d����)�#H����d�����	���HKL_,E\����e�%ZZ�-�炨g��*c�(��c�钿q_��Wz7ۦ�X����h�k��e�|7��x@��Uy �����	ދ�jX�<z�6-�{#�l1Z��qO���6b�~�XR��Yr��U���L��W5z��g\�e��O�U����[�i�O�|�����q�/�~�����6U�Nt�,��۰a�Ff��e$��8C�����G��t-�����^m#e �� ���ĵ�y��;pr^@��"i;7-gN��en"J�׍�J׽�����1�Խ�^^�����PpM�@�*�WS�""4َ�_L�n���wPRb<��t}]�\4Д	�#.�a`�	V�Tw��D=đs���O!I5��4=��Hc���M��_��Є4鮂�L
Z���Wt���NO������R݌���Wt,��n8��4�r4h��;9:��� O��:`��&͒H��ε�0�ڃ�֔�U��M@�.vƒ���h�$L��ƢN"��I*.9͌Ut�M�)��y�<:�E�X�9Rz�!-���e��:ml�ug�)�����	�P`W�$��68Y7d�%}L, �_"N�P4�D�Ӵ^���)�� ��ibU����+�SwnS�/��b�S�u[�a�KF ��C���oL�I\��׻~{Oچ�J]�D�.��i�eۿ����y�`]�����G�I&Y�}�˚�Fo|��F�)�(�5�Ђ�h���X��8�P���%�iu�M+�:�����:}j��⍯Tf�1���x����<�:~�n:��0J����jl0P�0=����#c�KT���R��0���jo-/M��mW�s4.b��4[eS��������r�<�]�ԛY��#L/�f֐5���8���- #1DyvI��,`����N��>lwP��*�S��{<�=��	r}$#C�ǘo����J��[K���i�:S�G����w�}���
��܌@���"��?������V��a��b0����J�h4��Y2�)6�}C
NA�W䚊�]���6���a����g(�߂�k뻗4��G���%�DN��lt��ڈ��Ġ�i��w���MJa��Hע?�'��9U���$#� x"?n'�h���r0�ɣ���ĝ���V¢����ؽR�:�Z�� (z�yW>���.��u�W��q&׍�>x�u���+?�˸���L��P���G�p9�η�����3^��=ؚdL���Y̸��xC�[���	<�!ÎB���R�l�B�>j)�����y����?<t�a֞*�E�$��~�GPW/����e+�/)O5p``�)^�Bu��˿�D`��Fa#/���i[��Σ�޼��d'�\��؛�y�|=�9�$yS%����F�(��Nɓ�Jw<����1����g%Y���6P��mT��ِ��L��4I����'w�%IEi����@�"c��s�N�(��C;�RVj4<Ky�̯P�4�H VO&[�/�IŽ�(]�,��|D�h��*��wQ&!J�[�Cf"��x�I����AcT�l�$�Hch��S]g��cH)\��t����9���C����&O�����(�&z`\6Ҝ$6���I߯�xG��92��uB\L��Apí�b:1�ޖ��}��'�l
��-���<�r��74�4a
gG5Q�	'�Ag�t ����dt�	���C]q�L���Z}��X��e��F/�B�4�j9�p��G�z�<�R�3�c/W���g1�l�sE��-�f�Q]���C����s��-M�P8��F���0r��xA���
�7G#��7)>� �#~���C]�_$Ql��i��k]TP�h�vY��48��~��?�t,FS�E4�e"�RX�6��2Y'��Gm��3~���OIܹ�����%�)ny9/��o�r@׺�k빝t�l�Up4X�lXk����X�,sTbO��9�%��N�������eU(W�b�K�T{=��E�wC����""�>#ЍUW�,�֑dm$Ō�THۑ�b��@����B��8���l�Otl ��d�6����X�3�XC��U�h@�O]�;��e#�F�s�)l��|�#
Q-iL!+(1��QbD#c�[A�!jH�:m� K��`�4��1�O,�R���C�<Qp]
+�  &�փ�(�9���Є��"��[Z_���z���1�b�q��R��՚ͱ�;?�- OӜ*�1u��,�	�;g�kM�i��p�踤�o1�ٍ~��YRʗ����]�w%�#��u��Z�&Y���AI u;1���a�>��:'�/ �T�f�`QMaY��#B��:`)w�X��3^S���b���=�5L��'���F�O'2Ww8�6��uɜ:e$�6�������\��}���8��
�7��1����x�/����Vh3�όUE4�0��M�Q�:�}��_w�0�rv���ق��\&��b�{h����(�1|��
]R�r^�;,�J���$2�_��)Ռ���v=��.E:�����ҡ�ځ4爧���֞�t��ԅ5�]hc;�Zm~^Ꙗ�)l(��|�L6�+26 �
[�YS7���Rm9b��Έ�I#z��S�_��I8��#�?ܚ��ژx�e	g�R7�D����5z���-0��,��Xb��R�*���� "W=
��N���t��>� �C8��yɑԔ�Vc���*B�W��L��Y3�P��+*�˝8��2%��� [j�y�?'ԕ��s8;�����K宏����MX5����F9KM�|�Ƹ	E+�G�e� ���bx�Δ�U.��ɠH�y�l�ˮۗ����+��Hz������[��7+]|��~^#Z�	T�TU�~���-�Խ��)d;n{��;K.<�sA�@|N�m�9�igP���Xރ��sP
HFL���cg���1r�I�����xL��·j)�gv�8���@c���i,Ŵlm����7aׁܭ�8L�������'�s���;�"j:[����sV�J���=��ӻP���M�Z�ܝ�i#�t|�f��Ck����N�5(��Ji)�'���۹���8hp�� 3�ؓ9���`:� u�9�t��*��oHȿ�&�wL�G�%�*�@��(I�����\�Ei�Ng36�+26 �
5��1�	��FwᇝR�[����{bgdR�N&Eį�DS�I����R�0�nn��o�}B�SM6rj4��ӽ1�Ci�3B�k�;����w[#��!����^�w�t�8Z��E[����0݇�5��Q����bd5����I# ����-ĒT�$ �n�*Hp��S�Q��S���J����3>��N�_�q8|��.�~8i�wz�Y�(\�_��F�`Ő�;0~UWH�pN����7�3�&��uh�m0��h��1
��9����32���9�{����eu��}h�O`���d�A1�,�$��6����vNii	���=� v������=�ʧ�)|�W���y� �w���L�T��5�V>j��[����s�5ĚtN#�[L�{e�Q��d���|ѽG07��é�NH�O�@�*O��'��5k& C%�̄-�49���!�^4�}q	rVT 	�
T��5L���%OC�N�O��2\��\ɾP*9M�*�p��"�+�ƌu�$_s+tu� ^���D��qL�7�)�� �<j�G����,���e	��9��q���5FPX{v�p������Կ�R�9F�^4��WI�q����0Ң]e �yq=�� P����;�l�F�ԟ��IJw)�"����3z�5�ʪ���i.�q�sCu�1S�5E�܄��H<�r�e���3��g�	��Z�woAD )$#���IBU�Ľ"���[��-1;�v|�c]$���?��+?��)F %�d�?n�G���܇�����2u����i����-��U=r���oC���~���>��ϒ����{u������0�9v 3��wbv�.��#8�}��%�]O')�Q�\���m�}�w2�2)�"o-V��a�2���:i$!eYH��G�F��u��t��ō�<RZX�^����������ge�(���+����0�&1�2!}I��[��La~"	^Y�r���|D�#=h��H�帯^�ٜ�E��ڶZ�t�������9E���穆��ĸ��Uc���Y>n���]6�i���5>U��O�#@ė�A�2��VY�-�٦��U�xGa���FZ;�#~�2X,��dت)qvL*�v��b���E^��f�E�'�U
/q@��
�
��X�
e��K+�CPX��#L���G|՞\�d�p}mjFu�Tx�Qg<M ����|X[��+$�t���4�Ѳh1F �!ZC)��1j�����M��/��2Lw�H,�ejx�����7a�6�@� U�|�|��j|቟[�*�S�@���W~��9���}��}`��]G����8�Lc`�)�(��f,�2����6#�׾��_u������l;�)���͘#AƂ� ��2xF��j۽���f��aہ����{������&���&h���y ��'�ΆE*����3�:�x�p٪u�1}����5�u�Нcȑ6v��FD�=�v^q�g,�Cp��Jr������!�ǔz.+�tjz�cy��sN��J��?�|lJ�Xw�%���E�tF3r�mt����*&�D<m����0#�P#N,_�X��cwF��v�Q�ψk�;@���V!��������������{z��f<Wc��ht��U�=15�ܹ�i��C��A3x�hX9�qze,W�"��^��8c�(*X��Oȇ!n��}7a���.J�x�Һ~�Q���������a{�������� ������Mi�D����Pf�[!���L�|I�rʞ�k;��X���t.p��,�`Eٌ+��@�t�p���C�&�����I'��&�/ׄ�&끩��B`���X���+�g����g.XGSx�r�}vYb�Y�Y9��2��7JUpc��	e�A��#�ܖ�GnC����>��o>����9o�s��H�9�JD]E��Q ���ܜz�s�q�nQ�_@bnB��/N�P�_�y�1��H"�����*��%)�l
���c�SF�B���׫[
�K(?��v��kXzK���T�VUC��n�}�g�"���r�	;st�|��������d>1�j�k��g����4-C�p�J�@lE�) �e�*;䰚����~#��@�/ܻ�),�9��$"�>�vaw)X����V�o�`��!��!U͔�#�g��GJތ��xGӨ�4���0�;7َr��9$��a�=���T��h"���2�W�v2c���K<`��*&c�)���J:�6�p��Ζ�:C�̰j.����DL�Gݒ��(�|7lۗ&)H��#*��4S���m�"9*H9%���"l����G�W���L�o8=d��Dˬ�]g��ΊR�\x�ݲJ�QS5z/^A1���]���.�
�����KGP�z��D7�ϧ�o���g��n���g
Iv�������9w^!���{~u�5[8'�$:�!�\�x�R�vpDi�wjHa�9")��	��(��9qa���$W�ӳ%�,���q��1�������!��ofy�|��j��(�|�-�1���r+,@����!(^�0;������%�/�[O�r�ޝ�d;�b,�c.`��5�dI��ގDT���F�T�[/kC���H �Ȋ�9;Ά����c9n"�rbu�5J��� �+����	��(a�%��7`Wle�r���gpB�}�=�ÿE?��Xbݳ��zlRWhl ��|>��:����F#7�K��/gx���8'��+(���	�����l�tD�	I��uU������G$FiOq���c~�84B�5J�*�B��D��$�n�n'ҍE�X�3��'/���tҁ$anK�o��q��w��vǌ�p��xM:�}k�q✔r;2�� 3��I'����S��w�0,ϧ�	x�~0�����"K�ph�)gL?5���~��t�%v�P����,%�Q[ߦ�Gu��b�<� �-�V�Ѕ�>��:y4�χ\�u��� s8W�7,,�'��5v�vz����ৼ���m1�.�:o�O�d�Y�O�kY���v����3!�4E�SM����/0����(|#rR�#����Vʠ$��i�sr얅u�1н�\�������J! �����G���a�YBg(���t�"2aqr���`�t��B���#mO�E�(-N Ð)�|�J$�/��B��8��@6����jJ���$���Xg�L��+�($%<�U�g�����)��Q'��3_aA��ci�n�g�Eg�^La��(ʬ`�&�pD�^�UKe :�H�ԋ�NS�#S���r���(x�����a��_��  ��IDATC[e���b^�ʠ������e�=tM��2�UάaI�ts!�o(E3h����S�9W\D�֓8`�)vJj`����R�'�?[�"��"���tt:RT�D#��¾ ����FXl�Ե��͛77 �@�b�MT�?�A���yw����{N�R���i,��iz�1��,�����1����y�Q6�xEһBt�ed(Q��ځ^oG���ta�P�3ѝ��*e{뱁��0����d�h���#Î)(���e]�Ň�� ��@O=�P�EDu��1�WTJt����'��ca��֔nb���&"���s2��y���8`��x���\�t�J���⺔�p]}p+<���!@T���{����$�e������M�ۀj��C���t�J`�8`�<���#(@4�!�}H`��iV;g���qF���=Ra���8�9}���PB1��m�qe=Qן=E5�&q><��jܡp޹me�9��kA?c#��-�v�9��nR8yp
w>z�>9���o��mPB�@�X�A}�Y�3'y��#�t���"�t�>X�q�Rגc�̪�_~��ȸ}hгľ��f�R�"�6>����&ir��4���t�����EK]v�	���"�X~�&��5��;>f���ThȎ����s�k:��v�}c�7DeYf'''�+26 �ꍨiʱ��4�ݛ>2�;4�U�Pz	y��"mL?W�oy<�؉�v�&)+ߛY��o��#p��}1D�X�D���u�N�'�˺�+�	��)�u�-dܡ����ѭ��
� � wHP�+�UP�?����Q��ŃVN�1 �*J���<i�P[b�����<@�uQ�/�����u<A��?W��ׁ�>�r�q��~�i# H���v�h�*�9��D�J��ƠrrF�F���0Ø�vXP�9��O�
�wGPg`ʂ�����F�����Tm9̒Q:Vy������k�<؅�́ �:H1����"��=?���\_�߱Hl�dq/���I=��6`ŬaX���������<^��Wu��m�pc��{~N���K9��m��ܦ��ƿ��L��jޏ���ȩ9�ƴ>�.tі�k��_a�*�1#��DY��ǳA^{ex~�>�QD>;i��H'�4���hZ�9�v3�V�[WT%���	�7���gUU������O>ٔ2_���Wl��Nf/9�v*^���*0H�Tk�+vѠ P
bU:p�/�����D4� 04��ʦ��Z9�w;�8$:�,�D�!���gۍ%�P��E��Fu@T�+�%b��Q��t���j��E��b-
����������ǘ���o����#/��';Ju��ڿ"���������Ӂ���4׭���yp��D��{M����T����h�N��f6�CPW�0iR��i�5\�	F�c4����P.gT�Q��c�8 	;��uN�9;��}��R :�e������<_%MQ��]Π�a�i��U������"��
��4��=��ߒ/uǂ�b�<��G�<)a�x��2�lad�}���d`y����d7����I�I���k�v.A
�(2��;Љ]��	F3]7L���R�Y��&���(�����7H��)RDG��^-�4�����}5>�}��(�[i�V/�Q��1��/���f]����f�����@�f\���Wh�4������������$�{�:r`�$c���)}�b�	��;#�B���=_P��$�W���Vĸ}��m�ZV��������>�&��X��@�#�ve���|wqCqX��r�����t��µ,5©��&Qh#"P�B�o�}�b�{d��ķ@�D۴zc��p>;�js��`�QD T�?#cYk��d�h%�w�нhb?��m��vO2��u���K@-E)چ7����z`���E�F�����c:UM��9�F3 DQhꇎիK%`l�e��y#LWK�ධ�꒺n �C;�=�eS�MY� Nv�~�8g)��Y����GP$��sԌ�Ti��wκ����g���=`cz��Wi)��f(�/aqR@�D���cS��@e!O�����5r�G5,��U-!�X���*HC�^D���|��/�ݹI��q�e���B�(��I�������?�\������#e�W?Y��Y���j5#����ｄ���֋�X_�fUϾu63L�sZZY�pY��h�0�-��֦�J�"z`s[��s�4���}���7�ߟ)2���<6 �
������;���_����_z�[?7�3�-Ws��q��D��G��.���tD��� ��-/Ê����:��BTTѶ���%U<M�� ��s�(�K��u���(� ���뎋�D$��U�G��6$]68J�X��28��+V����0�,Nں{��j�)��"�'梨��MU"����Ǫ�������ks�����/�N{鿇ߥ��4��/[��%��	�Ӵt'�"D(�^a�2��c�p�Z�_Dp,F0>��ُ�F]���uv��A'���`�rS*��.��߰����Y:D��G�J�0kH�^^}�=����A�|6�CG��(fG���;�b� �C��y3�6(�5Q �1��Y���%�yY�f*ُ��'ro�[a�
J�^�c���Ni��Pe�~8����{7��On���n�&'�K�>����G����ӣ�_P�Q
�iհ]���b|!� ����?z�s���1m��q��s�f���|C��l�|_�q�,����{�����;�1܌�ٱ�Wd�S�O��߻����EY�|�Pi��>�J��62�Q'����QB@��hKEU�q�b�MBMD�.��61�P�!�Z�@.��,Ajً��ce����I�"��J�>o��0��i�{�6�&��h��K{�_����-t|�.mμQ��	���՚(�s2.�OmD�;�яV�^�"��i_H�ǺTs�d��m��O��k;Љ�to�˟�����9�ۄtρU���`'��5ek<�� &���)*+��S��S��*�oȝZ���A=r��حaDE'X�Bܬ��!��0���k��	](��a	����-˿@ �����@�<i�?���K�������� ب��%ZO���I�d�W9ƧYS�	��ݹE�!�P�������ā��9��e��<_�q"hCШ}�9n�����K�9�� N���d��������7x����#զm�6��(��p�ݩ��SJ!kꫬ��I��Ưߨ��r{��q*��<�D�*�[t\}�r��m5����:�R�|�퇒�v�O��e>��?�O<6 ���KO�(�Uy>rޜ*��yD$x4>��=J'Ъ��LT���q�cǂ�*)�fW/o�Ip�3&�0�R���y18BN�C�5���I��)= O�! fd�T� C>�������F�U����8�<����c1�!{�-��]�qQd�I��%ey��qw�'�!�� �O�w�r�}�]"�6�m5����B� /�+�h�9�f���R�!�P�.H[�3*6���iMڇX�-�eTL2N(���ְ�7z@����I�@uD�V�;��8:��H�<_�p��K���{T��~�>|VIG������9�����Q�ݕ��^�<�jd�:���S+P�R���8FؐP��i��%�l�J�U�E+V�'�����o����{7��_���8`x�H��o������tgym�U�n��!U,�5th�m�uw�Ϗt�����,���ׁʖ!Yz�ؖ`�a�u��p����6�"�{����0D_��Wg�o��z����ՃG5F���z�����p�Z�VĚ��y�.�؟S���vަ��p6��Ҩ�
��a
��L��t 襋�J��@C�ׂض���[��'��RX��2�wk�z�EFW[`�S�M�=�Z���i"IAkE}�%Ҋ�&� lm����LG�ĽQf�y��O8# �ڢ�>�F�ȟv��a���|�,B=���>��������
�K[��_�t	��#���{��!K@!���\+m�/��(}��(�ŧ�Sw��=w�`Q��8���
���=��^ζa���sS."���P�+����� �l���q���#�ȳ����G�|����cK|FE=�5�Dc ���C�i�*�H��;8J���jR�-Q��8MQ�s1�� YY����}o�+�r@���v'��N���g���<"8����HAꜯQ�3_�_��$��S�Ll��^�4n��T4~?�����/~�{�/��Mn�~x�}��؝�lgZZ�4����cr�IÐ
�.4Ü�� �\t�°��~zP؄��nR�g@z��uӦ��=tЮ�� �����N���!H�$.������xn� ^�1��i����ܞ���S��q�2��� )MItwub��'Ec�M[_��Z�B���[, �x����}k#{0���u��u�G@`-�^�いtE�A���N��C�~�D��	���L`�Q�/0��p����R���s���'v�~"G)���<{AZ.m�nx���'A�*�Ǎ'�h�Om� 1�e����vg�l �)�����P�>�x���UM|ATa)��z�A��MݽX��c�'u�d��{V�o[�Pw��/S#(E��t������>f.YA�'f���D�4�� ��4�R��/.������ωm��g�#^,�
�iӭ�&-��GE��	��L�Gi��[v?�|�{.h�E/g���B��<�����x{���wn�����������kw�忾Tk�𨶌s:���|W&��i�]���y���G]����tErC�J�Yu��E�ÌK�� C	*�TX���Lm���� ī3ԏ?�h��?�����as���Y�;) ��g�qv�[	=�>2�ZaT\.�*��}��nŔ���NkQA�}�ɏG�b����X�9�N���� U�G����V�!Hg��� /\oC:�X�YSW��v��!g���|��|�|��������`sCl}�)��F�m7��Rw��6$?"DtهN�� jϲk�a @�~��݃���A$��'�6����p{}.���f]?�|�v�a$�D����0�����kL�,qx"�̊�p��O�}p�1v?�NK��	��4���Şu�I4&�ý��s�2�%E1l\����X�q�2�'p����>L��=����b�L�� ��x�6���CǑ�ݢ���fqk�;/�V���
���2NX�Y�Ɠ����{6`	y��t'��/�@U/���!,0[�#��@	C��$���x?��'���{�k���J*�ҩMv_�7�������}��k�o�蕽_8����0�Q��+�D�(�M�����`��J#>�к��� ��碿
쌷˨�F�؉!8��D�H` q�+�9H/KRl݌+16 ����G5?��å��eQm��Ua%3� P2�����9�����*��⩢m�*;�猣6���� -��g���*�Ž��ֻ�RDm�H�����Xv@_q�j-�O�b6k$�M�LiRcV	�Y<���w��`����)5.��n;PJ}m�3��׬��8!�X�_�B�m��`�K�}�Y�����$�T��l��_�+���Cp�n[��W�O�@־�~l��\J������'��8:�J�-��@�uNJw�:@��#X,g�pbǖ�{@���8JM�Ӊ���;Ư�C)�[v��ó{�8�1��!d�(�K��#�^'W#\ʮ���Q}��*�ox"��v[�k��HnK��{�:��<��`����_T���c�O��Stw�q���ݚR��h�B9���H���Ii���/����폾�/��5=R���4�^Xg?;I��*V�@��p�Mi7�v�A\9A�v�� ��P�u�ϯ���3 �wC0(�Y:h���=Uggg�l6�6=���� �+2��[��[�TU�{?���i�f���Е%�A���,#��r/u��W�mԥC[�\��_���z����=j���x�
F("@���v�3f��4c��![�f	���/�hUI,@0H�(�QK� wQ�@�TdS7��uP�f��|��h�3�A!{�(�QW����P/�nK �WŶ禍R��!W�I�h'�˃E�h���Ee���u��>�P��M���Hp���ߔIٞs.D
I6�W��um��#D&���ٞf5��_��g?�j6����5@m��"���+c�O�o�G�8k�4��D�ǯ�N!0qΑ����Ϡ�}�|[��/����AǞ��+�4������er���ޭ탛.r؝/ (}���SWr1m�	[gq��C�oܗ8�a��L~��N$�U�܊n�;��v�� ����%�On(ZY�ʝ����m�|������L�-��`����k�߬��������i����B�f�o�j��0<|·�3�
@��ѕ
��Ɏu�R��ΆY�aEQl���x��o��oL&�ߵ*������b���)�eU���	�`z�|�$j���=��
�Hu�i�@�'���H*&���3l�$��-T�{Yg e9|Q%��������<r�2�������^��K)[�2�Z.���c���R7����֞�S���y�਩͟%���@q�_��n���P�Lu�9�@��|��	��.3`=�������y�_�}Z�9t`1�'-\b���w"b��`��P�����W�|���p�y�x��"�l��ti�w/�	8Y�BEE@ 
#�T)��X��;�G~'�뇰5�c�I��V�@S�T��&+�j|Z���m�jux_�����U�j���Nދ��E�<��=H��F1L��-;ק�QłE�Q��A��u��@CE;�2!�\�B�F��OF�n³�����jF���P��jt�������w���mh���mC��:�����Pt���K���b��[���a3~�� ^��ܘ�?��ާ�~�����3�װ�	J� ��,V�j���hd�U��:���1ȱXߛ�Ů=hT}@B˙Z��g؆ Q��b�ցBYN&��+����B�ۮ�s]�1��(7����������k�7��,b�F������hZ�	*��_s@n{������������5#hc؎>73���Gk΋ v�խ

��߶���������q��C�>C=~��%�g��c8��.�l�4�e�����Mʈ9��|�c���[�uHU���+�����G�ރj�1���َ	F6w�+�k�b(��^tY�6�9$^`w|J����U�`�5N�V��`��|M�P��c�\�ـ��q�Q��H �"�I�vϖ;�e����,o�-Gau����|������~qO���u�mKE�%�V�l�Z��)|qBB����_ml��E�a�ćQE����uԜ>�Qy�4j�Jr](�D���L&��hT��e��� �+6nݺU���â��gK�򲤗�m�2� Hc�W���f�-�r(ʥOoV6�b �/qC�'!���>�Y�	��=7E���S!@$�����haY\���$mI[Ai(C�)������*��,�ȼW�9b�$�I�������<?��ח0?̪.u%1�5�.6-q7.`vv㬄,-�h���~��� �w���Xoٓg�O>�"$Eq?�Xk��Hq��*V���b%��a.-����'9�_�`��;>��h�H�d7�!l�Ş��%C�f����M�5�)v���m�b������=8~����m?���)d�;���[*0#).f�B5�=P�}%�_���=��	�z���n{�\|M���6��5GF�+��v��G�	�BQ3�T'] j��(������Ƃ;���8넣��]�$n�cwQ&���S�?{o�kە܇�Z{:Ý�D6��T�bK��nY�:�Ղ�A�_� �� @��| ��p8@I4�"�n�-K�вe�[=���#�t�{�=���U���>w �k���O��sϰ�]뷪~�+���'�b�6�23�A�_.��8�o$n�E72�@�r�`�b[$��� (�	�O��ߓ���U�U��t�;p��Xwrb��DiiW��}�ɓu���y���5}��W���Y��mk����⊅O��ұ_��`�lS)���Z�l�)�`���|>e�8g`7�,UP��!�!ҝe�M�^(ht��)�O���ZP��I�q���ۮ�D���Ĕ� �V� +VZ�$���j�)�X�׼@p*����<�6[�q�I�^�D�!��2��\{
"���M������vb
I��Q�,�m�'�5:\��C^�P�r��m ��v��-�S]�<�9"�2p��9!Z�Ϥ3�f��Ԇh%��p�<�������\�r�z�>�(d���`�!��p��*`����n�nQ�+M�����«�a.�[�<���/�p��
�.L���U����'~~�2 �Әs�'�F�յ�'��H�N?�!�ل����=���vA����s:<��po��)����T�#)�X6<��k�/C�EI)�<;� 2�ptz�=:9�U˷h<:���1%�v1	
��.\���]_Bm[H�"��3���W�&��̴�;3ʸ�%ka����1FR�I��}�����K���R���z�^�9֘�6r��M��lp'��;��h���q#9�0�M��޸�~� ��?I��]� ���<�3�Hk_J�� �p�nk���4�}g^�,H"�^"ɹ����G�՗��t���h���X���!LZ5�*��ƈ�p^��hbQ_&�]����hZ�^.��J  ׷vp1T��&ϳ��~JO�>��kkk����̿�;�Q�$�j	�&��d��d08�L�+
�(O�U(U$6EH����
*?�6u�ORx��d�Ĩ\�٠�'%3�~�l"I�����H���"��izCg��
ZS6a��D���C8�]ղ��Z��%�BY�m�d_���I<Q����f�� ���%�F�+b�ؖ��\:I;e��9��@�n&@�k�Q[���w��Ͱ��4j�����S�X�8�B���'O�=|��^��z=ʧ�}��6���T��r\�6!�e��F|��ո��^ޣ�|�WJwh8�h8�T�`�$[J
?i�ȃ�lv�>�.ͧoRS>d�uFwnoP��}��q
��p^����>�׺kel�s�>n���&0"��~_iA
&m�L�=�4��'��N5���	֠�϶�zQ�ȚEeI�{6o2�<�3?eH3�࣡A�ǹjlQ[�P��?e�����xAɍ�Ez�+۷��郰da��ȗYF����QW�~1p�H��f�'�T
�|=T�<#x�,)p�C�4$���-�"��X>���F��M ��t�A���~���� N����r�k���5@|-�Ғ��b:�:�y-"h���!��&i9$����T��a�De%o�5"i�:�����pp^S?���#��X!���P�Jžx+ݭ�2.F`.���2�t�.I�;>�7vHmlx�P�D '�6<3F;4k�K��?S6��@���U��$�C���r����#]ÃW���+r�t8�@oD�/��1�րPi���&yo�ol�m��>� �s߁��2�ǒ/}�M?m���6�vRя�ڶ�������#ڻ�%�������}z������6mnސ�)&��8�eE&��J��-Nx����D�7jmh4�9�n��!�H!
�ۛ$TS�a�ň�S��G
�W&�}� )�%�hZY9:8����H�_��;�)��gMr�{dw�>�y�/��o�wn=v"��1�Hm�ʤr�,/-�kr��Y8����+���pa��4�Ű�u�Yy#QRL�%�+9zY��֐K�w�{ -����$�'|�e���O��T��ZOQWQ��]� Ek������.�O/_E�!@ �M��ۿ�󼢵=��Ϡe�p� ��������*����D�����sF���4�Lhk4��XHXI���F��D��s*�.V�Ay?��:T3Jd��R~�N/��JU�}�/Z���wH���y�]�����L��@T�D^W�+D{TjV
m }pΌ� �+�R0k������)����nt9�z��(�|��R፴]&@�U!�����	���X�>�K�e&�ɼ]��nY���yQ��4T{��4i#9�Gͮ���\��@e�Vy�O�m�"�a5�fZP�R,<O2D�oD;7�4|�T�xFu��M����d����j@o�5��ͨ�y���{~H��!�դ�M
�m�mK�#@� 4ܕ��������1"��4K�%��ٯ̗���j:�g�V7�7�}gӯ�v���s�~e��g�����=�[����}XR�iU���L�5��h��vvI$���T���["�q��q��e���O%�\.u2�Jw��K��5�U�W]߲=AJ,�~�^n�N�~nu�[.�:�c��~�m�A+��ɰ���ST*�ϺkIO�YA�����#�
r���|.��
Bک��A�h�\#j	�Vǐ�_ƳLp� 8��͏Jr�ҸK��	 _�uH@���� ���)Q:iS���*� 1r��#x�oh���.�Dj]��T��^�a"�5���lЪ�9�qv4=X�s�����"��!a~fU3H���ԕeN�Y�|�D�E�J �\*��F���l��h���KҤF�8ƷE���Ք`��K?oq��#G�],>�x��D����U��O��sĖ'���Å�n��ZTP�c)b�6��vJ�f.��糚N'<�[NH�#=r�Ai��2��3�@"@b[@���(*�����k\S��}:�X%��ۭ�M���O���D2 .]؂�z�O��6�bw�㿻q�����o~*���3ߧ�����$��r��&M�A������Tx�(bs����W�$]t�����L� �$�Q.bUi�+k� ب��:�����9\i�p���n�C��f���^UU������|m���3h{{{��ͭ�o���=��q����M�����rH%�@~G ���a6��T�X�X˜���A�]~ �=I����<D�$:�(� �x��ko%;�:�N,�Z5r�T{1��ΐ�H�nǪ�V�<�䔚2��9���ޠ/x��|�ԡ FRp��J�h��H��
���Lp��6�d��)M�<���h2-y@Gc��<`oP�	���o:����mm%"�T>�C�4�>6½��$i��:aO=|ڂ��Z��X��X,*{u��C�Y�
wW����Dd���F^А�"�	�8[��Z��+�T���UP(�Ted��I �r�	o��m[X��m���Y��%��B�zD��k���9�qR'�?��O���^�ܗ?�w>q�aG/3[�n���U���b �:����	�?�i{9�&єr?��T9��p�@�iw/�D����F*O�'ݜ\��"�&T����'),��`�ї�gǏ�`0(�Ӵ#\۵�5@|-���x4:����ɔ�����m��������B��vs���ѫ��bJ�2��x >/3vb�%�>�H��!:&�<��%�
��ye0j�F�̙F�&�JSu�& ʖ+U0FY�����u����5]��l;�~.�3u�&3�"� I "�-q]�wš����E��(��@V#O7�ȷ(�2�@��gT1bG�a�64 �Nz�#Ϭt����|L���2 u�ܭ�����!�^taP~��8E��*7t>��}G���~��K�I�=�`�*��z�\f'7�|�� �P#ׯ;������%�- 
��%2�m�1��:\�6���RݺTQ����\S͵Q1Ţ� ���6��z-Ŷ{���� ��pd�n,���b�kN �h��P���߬��y��?^����^��╟�oO�Z�X�M��d���T��dEb��L���"4�p��}�(�_��.^&�n�J��3H�5J�qP��.Q�^�F�x��mQߵ+=O���ڠJ��x}�P-$��0@������ >����1��h:�NONN�����vnޢ�_�I{�����T-��ᡐ�糉V3.�TA��s7�T� R��$B�ܽT�rI���XMQ��Ӆ�dZ̵U���hƴ==c���XL#�}�pY���m�(�X���̀�.m���B�5�-�I�&�TF9/��Q��H,�ڤ8���8����F:��|*66T�bk�=�v�c8$��)�mn�4X~�JW�F�%ykl�y9�P���2��4!?x[-�j;~ؑ����gth�k�Kk��Ӈ�
B�R0��WW/eЖ
�4T�{�oH\\�f5Vi���0PD�z2K��v���D��Mno���O��Ox�� �����p�eqA�����ޝ��|j�����um�!;3��_�p�����_8MCg2������*�QQ!��#F�LL̛�<���*Z,K�Q�hQ�V���H6���Pö� ��d�?���ב��<���,��c�[�g��ܹ3/��Q�������tl�|@/��Iz�㟦;/�$ځ���4�Ym���A����#�F�`�H5��6���#�}s[�MՔ<3����R��ז��#��T%VF�!��h;? QT6C�\�!����;�'��,�mƿ�߳�IǙ,I�R����V�e$t@����/b��#�HL����C��Hd�r!�ǭ�H-�jd�޾Z1A��wD�����#m����ID��2�0R��r���kM��)��S>��6��bʃ<�W%��$ i߂�6�"���=������j ��	�2���\�.�^٫"��e]mW��M���=1P|Ϟ�L����<�L��=�%�;��b�6�ɇ�wc����(��Y�0���SNZE��De��}��+��oT0�m�=�d��l_rN�h
0�h�RDV'�"�����g��$��6���8��m���n����&��	+|[�>,�B����D_u0ʤ��5�*�a"�C'&�'��'�g�%���X��4<+���:�C()�ym|W iG��i�F1F�;��1����ʰ�IHe+�,��d�>�u�ֵK�����5@|\����#>O���g{�I1��)��d:�l9pWWjjy:�:#�T*;�L&e<���Q��4�W5��ZR��;���3��Yl�&Jt�@�,aG���/d�-�S�k�ۈ����k�v�¬��C�|� ҬjwY��&��o?��t!�9���%�#���(��s!R�[�V V2�+�^^�y{�\ ��$
L���j���2'��Y��e��攌K�!��a� ֫�.��)$�4��v?�`�����=8<'��ò�[y����W����m#Il��#����	�^���چF�]�@|�p/�����#g�gVh>t6�I߬z���)F������|�}Y!#���L�[�{=E�_&sK�^�!����%��j� ��":�Q�x�HZ�R�д��*N��{M|Ϯ�ˆ6��
��1�KA�6
ɀ�����`��ψ��3j�7w�|���ʳ���?x>qsQCu�� ���,����|������7��>�3�������0�4 DT1/�RRSHCM'�����#ƈT�+*�)-�����h��ruI˲f����b���>�M#�����j�S��f�Y��N�E��U�G�r[b�x;-,���B+1<D�Z��:ju��5�Q�T�Ę���GN��<��@袅V�6@Jh`+YvS��a=�c��B�e�<�&�E;Qr�q�|���� *~Ͼ��	]?{r�cV���\��k�.������~�&<���#HjD����V��)	��޿1�����潸�W�}p����u�r{���˴��\�}�k���y2/���_IZ�p�9�vFϗQrOY��l�g*�}���($��V!�/
�s�U4_TTչLdc�~[�����&�R�BԂ?+`R[~��J&�K��c;T����Ά�	�1���[����5@|Fl�Q�{���o�������f4���85�ݝ%�ђo�e��U�,����}tt�_���r�/K ;C*���퍩��h�9h)��eYK�^'�BR�K���iI�'K:�͠��n
B��9\rJ��(�f�j$�Cb�}M.j_�!�}Fo���s�I���q&Mm0FJ

��ǭ����i��LM�{9�6��hT��t��N�{�"��w]1,%}�!U��[����	��	�t��s8w��'i�i��iю��ڞ�VA��q)?��ak�C�c�'~�]���'.�F����2���(��q�
�P�k��s=�_�,�HXx�{	�C��?�� �q9ɖ����,��P�p�TA�+�E�p�+
��s�,����M�����ST/:=Y�r�EY���>Mx�e �*�/ٓ4��4Qʈ�֧0 C}4R������ױ�<�rssc��+����=#��Ϩ���ǥ������?]�{���'߽����Į��߰0ts���w�<�K� %_-��:�0xYB7�A���N��|��y8��%;�|{w��O!bܙ]�
#�X:�hE��J�`�ʎ0͊W�, ��E�(b�¡�����Q�M�}�)V&��M�_��il�8h��b��T���>V[�����|VH�	��Ά��$eV{>��$r�Db"U�9H�$���F�B��. ࢆY�^��x�+�I#�?8��kemD{Uw�I��S�]��rs%�֩@r�#j����zM���j�É��qY��;�_o���^����Diq��X!u���=�7�-�26�5@l���t��S�/6P�[7ڻz�I(�s�	�ҶST1��hPXz�7�p��B��:�	&��d.f:�L��<�6�?
��q�T���p��EJ�Dh��("~���hC0,�c_��4����=[��a3��o���~0��OO'����^_������EB#S�;�f`D�pEZ�%+��\�������t�hA��n�E�{7��ecc�/s9�0V`EWj����n�o�Jg����YQ�����g�NJ���}�;p������햶�ɚz&I9�K��)E�nC�ie�A"��z$�*O�mN�#&���#�^Dn%R�~��Nf"<�p�ؙK��0@z�a{���E�����8I�/�����Z����Gc�h�E�h�t�5�\ �͎�Sėec]�!��w��\a?`^��5��r���^[I���kBP�|�O������Ɣ#߁^"�=p�����F�Y"��	�櫒\Q"�1	?�@#��"D����'*�x�m��P �������ʵ�[��OD�- D�z|=��i�q�e��(�=9�em��� �#n��xv����˴i��aGS�3*�'Td<;d`R���W���'�`��9~@f-���t6�T�c�\&Unh�4��*MQ��-�����D c)��Ym�z�%u������H��� $�5�ϘU� ��ޯL�^����J۪Վ�����=� �>�(@dT������*����Jlt(�9�<�����m��z�)iTT�j%��U���E�)~�K$�>>���*O��ˣ\��=�u��Oc+4���K��W-�C�z�אb�0F��)�^�.Ld\��&0qzc�m7��<�	������B�ӂ�fL��[���#�x�`��k�.g������ܗ&����I�
dyʓ[4�1�RBu0���d.�1m�'Z��-��d"�2������_H�Ԡ���m؏�G���<�{��DVF8�\��x&�U�8֣�`4�c� ��5@���x|c���sv|2s[�yA[�c��l�ps��4*yH���P#v��Z�k�B\*�+x@��.˅�:����\L��EIS0@L�S%:gZqS���Y��t�Ob�r�-a�\ͶEQ;t���<u�n$�2��G��� �	I�\CII��P�ngB���a�q`�.�/aЖd�j%=]�wdoc�	@��4��P�2����Ҋ*g*A�� �@����`b��y�RI���U�}����9�}���=F&�M��S����)'�P^�ꄬ�>�u�.�ҹ�,��V�+�ǥ�4E�c�>Y�`[w�A�g����[Myz>���o5��O2� �KI��P*>�n��F۷[����ON�t��Qc2�6R���%��BOg�s���D��U�m�ԇ�	5_<e�)e�Y���G~b���y^<��k�K����5@���b�0������mn��( �F�� 0h<�`"��g�5*�ٙ,˥T( XC�i��N��$�x����ޠr���&�����x�#��:k�(��7hl�,�*���:�tթi:$k[�!:	�'y�"��M��0��m����Q���`������(8�D�'3j�tWK52���k-|���d�K%�(z���vV�D�%X���kDh�0�k�g%���V���3IA2��$�����/QL�c��\Wp����Wa^��ҍZC2�r?a�hx#|���A-D�t��Gn�k�J��W�k&���*n����������F'���vV�r�^^���X�&�vt���~ث�A������齟��ݏXH��9�]�$������Ő!Z�� ���(�Z���'¸���p��a��k�dq
#�wA����8A�7����Z�,�|'%�;�|�>�߃3������OsG��!_���d7��>
�ㄯ��HV��DwvӅ�������H�Av�7	2'���.�hnp�qt�J4FQ��֝OOY:`_>TKZ��������LpL�~,|�p0X�b������� ~čox�û��MfK���*����v�6Z%�\�����Hj�X�gF�K�����f�mmhJ���F�	��g���P<�W�Q�.5�͚�ɲP��U~A�l{��U\7��)	)l���2�3ڐI��EJƸ��"���3��>G��&��V�N'�-ic����4 B�C��j
�z �'s�j0R7� ��£�����yD�N�д�r&DYðl�Ãb;�C&�?[�����"ưZ�g�B�B���>�����Q�k�6.�9�ƻ�{�%��A1����	���J��)��j�.��Q�u��vzz:���K�Y�p�;�:q/��U�
�SR�}��PI�[ȄR���0��<g�<䉰e���c�$�7=�d�K�VTE"�T4�yU��m�cbщ<$���Y�%��<�À�3H��/>�KZ�3ck��7v �`c<M�1�R@"mu9%?�I�������e"�B���3��@�S��T���h�b1c'�ݮ3�@�؄{ q�N$�B�) �:�e��Z].�u��L�w�{A�61�+�Q�+�5�e ���Nz���|kt����wy.�ߩy����]��}���hZ:J{q�1��D�~S��ohW�V k����Ç�i�?Θ���ժ��[�{l�c�ԑQ0al��D@S�A���9�Fnh/%��?���$��O�cW�z�tvu�{���}��P�z���uÑKWS���	P8�焟��Z�}2"�����n����R9�3h�d���z�D|��Hz�}�}*R̉uh
��}QU��w����|H�2@�M:::��	�ܹd�mƤNe$�������[>���AE�O�(Tk�(8Ԩc�}�I����y����?��ϖ��g�� �#n�f]�w�'�ᰪE��oxW�#[�C�F��$�"R�ehDR+��L�7�� ���i��C,+:lu���J��Ry�t��YBA�UӮ��]�N'����Hc��G��mД
K ������������)�#-�e�d]��q�0��T�F�\���ަ�9R:&DP�DE�Gx��1���*��J��q%i%��
��Z�`�zխV#�Q��S��D���k;����:h$`4<���δ����MH��9��T
(>�~؂������ @b����soC��r�]H�K�-�w;Qr][���tr�����O& v���`ꭐ �뾑l�(��	�N�$��[Ꮵ�%y��7�ݠ��NN1�w"V���#�������?kbZ��#%'fp�����w�P|?}.�p��`��{7��~�O�{��W�}��![ď�C7���T�R�tS�E9�*X $K�D� :|F�n|BK�U�Q<
��؂):�6 H�	��qI �Eђ��H%���܂	���c�3�"���|`=�L�lYbp�y�%BZ�p�g�� �,is|B�h� �KZ���&�hV�[��=m&!�:��H�r�;K��l�`��"��
�"zi�:p��Z��IC*8$�!��m_!"��[�e��&���=�^�K/-�%rH� �BP��>rM�׉TI��?��R�e�I�ۥ���|z������'�?֧9\��.P
B�@?OV����MRTF�ᡭ��O�ʩ�V4��?c���6i���j��R��ʓ"a�X+GD[(�ĩ�����VI���H�)h$jZb���μ��5�imm��ĺ�h;ч&=�);��,N_7��`0�c/���O�~�\ݚhm?���q���t��x�Ρ�CK��'���q�C��T��P񫼚m�L*^��z��
�
ҶI��
��^�e^���[�����#�F�
Ҭ�y��ә.��!�u�����m�ЀwSd���X�mT�̄Ԯ5��%]$�U42�
��4m�6QWA��;z%���#�L&�7B"��m�Gl��)h��Kw/ܘ0�F���S����c�<;���	��8>Ԩ�p.$�iM���x��\�p�� �w�G$��؇9�:ݜ�(a���K'F���]�I��� ����
F��w����S;Z"�����{�dՆ�a�(X���&)�P=�
�;��O�~s����%9-�9=|8���B�g-�Ɲv��Yߞv�ܤ�j(���y��22GQ$;B�l���U��+˅���=y啗_�s�'��g�� �#n[[[����$˓f��~'V����3h���R�������T&������e�ߗ�v��w�3Q�d��`V�X4����[7�nv�Ö{���=ᾘ�u`*��E$b%r������'mD+�h���9�z�5��;�	mm/h8�jf��
W/yD�
�� j,��T�2p�������:��m�
����)
��`t�6�:?�|�PN��>�۠�ؑ����¼׃��k	�Q`X�k�I8�����;��r�J���š�J���]� ГZ���l��6��g�{�)�����#!$�촡�1]S;���	_����0�)Ps����$��0N�a6dW3���	>W�RyB�p%���:�Z�J����LHD��>Y
��䵟�qA�:Z_��j,��
aQ3�u��jgw���~��o|�_��ڞ)[ď�4���0ϳF;�$r���k�F���r�-����9���f���}���N��)R��n���;�B��x4��v酗^�g���rm$Q���T�c�q?��+�����AF��Z�oT_��1M�#�Y*��ny_��J�Q�izE���gJN�6��]�.��0 v:���;vI��E:����FG�w�,���P���U�!z����lSȮ��I�::��&GX��æ�N��Z8cñ�v��r�����Y΅����P�~<]6�6�z}�����(i��>��g��b�;i��Rt��_Q:��J%<?I,�tT�����>�e��B�1�nA�v���ےlnCf#��Ő.��9�ܕ�]a�%�S� q>����f����㚤YKّLM̮PGS�ɲ�~L�8FNa,J���(����B|6˛{{�{��O�e�(��g�� �#n����_��_�g��u����,�8#G'S*�*rU�o�>\R��,�b��|FKRY1�y���� �����6;) 9>>�|PвR"4�X���`K�sD��V�/��ŭ#/Qb'��ݎˬ�Z{FI��������UЍ͂An.�˲�#�
m�\�L>ȴ�6`�4 bC�)÷]���@!�p�`)�&�Ԇu��-i%k*���r/�PX���D�*AW�|�k�Q�<p��*!��qUЮ��P��� ��i#�o����@�86�q���P�őtT���8�hd�_�M]�]{�*������e]�>T�����F�S��~����`�����k�QvL�����xgr���X��
�g��� �b 8�u>�4�ZD��I���@���������YF���N
z�?�����K���&������T�j�n���6T�cK��V.G25�^x��ಟN�$�9��{��7n�ܿy�3Z�3gk��6�q�������7}�H���20|��e^S> ���c @��������R�YB�h.����wޡ�|���a�K�2��Y!`�<�@��V�B+Q@9�>�*'Q��@F�u�0�����zJņ�ͭOЏ���]�z���c�?F;B����Y����#�]�
MAwQOZ����������~�=r�b�P��>�WR2���خ0,`��S���,����')	�[LH�k�K,<��o
ʁբ��|&�`��	X��rDB4XzL{Ն��UI�k��C�^7���&�W.(0�Y�4I��m�x�Zv찓w^u���0��E
@X�\l���_�nJya��D�v�:��e�ѝ
�/#��9ߛ[�z��D�k����I����=+1q��9qr���2 � ��7��ٿ c�r0���c���Ϡ���������E6c�g�Y(����)U�Bf�.�ٰ4n/��\V䴬J�D3�?MY�;�٤����c�4�TtՆH�`����b$1FaQ;ZL�F���yѹ��Q`��_Y�):<�aG��Ռ�K�G#�%�9�P�+�A�Ӊ�(���|�v;����P�aƻ0�y�W*Q�����w#���~��iB��������qnH;���z��%�� �FDӡ9雰��U�<�h�^��ɔә �1���Ɛ��1��kW��HC���`b��ڮ�����Um�J ]��>N����m2�L��5��N�G�p��1_�隙��W�{����9z����K���0I�lDY	�ɚ�D CH\e�JLh�؅	�R��4�l�٩�7��/�(NA�i���Am\�E|��A�P�j9αE��|��C�F�J�����
�{.�v��=����;k{���k�;w�7o�x���{4���j�=D�,Q
�׈J!���P��Ȩ�_���Tʱ����D ZEe*c��z5L�:�z}�V����KV�`��9�ե�N�$�km_c'=���mRw-]M$�i5�b��^��%gL��	io����u��FS�^+U�M�ZDY�D�a_v�ݺ�%�.�س�o�]ZE��c`*�J�����4@�Ʌ�b���d �v����X,������?8���)MON%]�5��&�y�yڽ�G�F�¾�
Q-�=�=�A�	B���^7f�j���!y��0!I
��䴘��l�uD����?��r��oevɷ�gX�\N�%5���YJ�Z��S��R}؊}�R�a�#��f������{<GGd1�.�֯L��{�7�t��>�#fU�w��! $|^�`V��e�Ϩ"��/��)�imϜ����W^�n����;7n|�9<�T�������A�U��1�WH_��N��"լ�Di�4u(�v~ ���now]T���&��g�ED���Ү����}v>M��b� }�Ь���o4"�	��*Z"zX/x�K�Xh�"���=o ��q�sa�Qx�x%�(ϚVV���\U����d��e��D�'p��n�ӥ ��֢�.�A���Ԣ�(�y1,)�T��.����tե�d �WX[Z�������}:8�S�(�^T�eӅ�#�n�j�y��v6�z�~�%%�Jw�~�l�h�����K��=W Ы"x���ë�a_��J��b��� �NZ�a��)�lٸ�?غv�C������U��O�i�0D����h�T���g�#����ܿ"�Ոn��F
�Td[4_�|�5tp� Ό��j�r'+��vj��@`��}1m)~	�ح*�~��բ�X���	x����%tU���3hk��6����~�׾�����W޹��O�f���N��1���rU�i���iǄ�� j%n"3�$������0P9�L; �g�/$u�뵬<�$T���0�Ƃ�UI�>@�wP�CQ���8�K13�Df�h�y�df/��؉��s�KzH
0 ����#VK{����oh#�?�Lkh#�2
|sA*��'�~�Ik�-���Q#1
� R9�P���@��B ��p[Mcm�+J򁤊5����Z6��S����9F/ņ�������cz|���%<&����4��򬤓GGB3(��;�S���#��BNބȨ78��G$��`� L#�JV�P$
�$Qu�z������aY���p��vw�����7���/���9+���Dn��CNc��R��9�-�2/�f��j�+�D��H I+Ӝ'X�`�?����S�Π@30�P{�?��R����{���]��9�%���@&p�/tϢ?�'�As��8|�W�)�g�� qmb��+�2y��������~v���i�=��JwM*���D��O��H
��$�"�������bu
�ІO"g�T#	�R�[m����pc���h�����M�Z��:��C���3�Kk�Z�*�8�z�9�e�%��h�F��,�ѻ��+g��q�,�(��P�����ڔ���Gڏ@�b�R��F\�U�h�sl�Gog_�c)���tS�w"�,�гD��rQ�P
����p(Ք&-x���b��9�����hr4�q�Ҁ��"���D2�4����tFM�F[#��v��,��$ ���L��6^�y]z��Y��:�*���B�H��)$��,�yY��o�����(����o�D�|��x
�(�U3teqc9��42�4
!�5Z�7���IN�r)���.��0�\U
ʬ�;���[�(U�+���b9�F��L(R�����g?���{�>֏>��.��Kl1��S������hs-q�� �M7�W�_�у�X����r�7H�&��X�p��?8��iH~�ݓ����f����p>"�PG�3�p��%v�q=���a��z����n�ob���A���: 5�i`*���BT��U]j�h�:m)���
�V[+[C�x���=� =Y�4�F#������ ���gb�����v�mút=�D.%���� �1�|�ÃS�a��ivR�[��C�����*�\��ݤO�������֍�GD�W3�\����&���̗4�s]�6dI��n� �Q)ɻ�h����av:=L��8�.Tb�|P���gQ�u��:����K��s���q1���s;������o����A0o��ݹ��������w�݂�ٞnf<�w"uw!�mWO���uҺ�T�}��h�<1],�w�r�Oo�z���������?�m[>�x�VF�_>�)L���P`_�s0��
d�ѫѻ|�88�z1�J��^P5��J38���>}�xFe�S��!23����3R�̓�JU��� ��%��L�C<|��( �wٝ~3O�=�����7߼y��-_���5@\[k��{�������־~����?ߞL&�6��_ʠ��:�r������A��f�D�MD{�]�h8�+�f����y��̶�<v1}j�����[�	���}+�"��np��,��g��:�
P�)d_���P\�����tm$5T�Z�b��.2�h%by�����# ��ʳ	c�ύV%_������#��C;�'jem�T-;�ZTc����Blu��?`��S�Q�:������;��7��/��.�Kl��o��+���Џ����[<�%KYGYT��(w0x�(Ԉ^6���9���5-=?>���.�9����:��v�H����#%���8�ᵦ�5��&%��r>LH�_��� $��ju�{�st���ID���q�[�]-���د��b!&(���>�Z=�>�.l�i���Ğ���7���g��]�] ��p
(|�v��xK�=^�H�Z}/�P. �U���$9�� ��tH˙����'/��1��vr*'���3T��[���V��&1��b.*L2���@bȷE>��~�(��:�(1��!�^�e]�?�4�i2�ј�b�C�K�{���OP@��@��J���bWmh2�4��� mLI�)"�x�(a�,��Ő���kr�8"������k)�����xs�������imϤ���V�K_���t:�g�86���o������b�`��Y.��=Z28@�3�$9�F����ߧ�A$x�h0`�j �/M�X��徒�<�*az%�2��wV;H!	��
��Kt&݈����!����u"��R��t��p��s!L#��]��暙�8��'?ɶ��J�ajAB��B�j3��Sc�R��ZD�����<��}�>էhq8�*u�o�!�|����K��h|�����56��/�e�] q�l���R�J�/+)3W�R�t}�:XEN�!j�~L%kRx��ʿ&�y�6��&F����shbD1��{v��]uz�L]f> ʕ�ۅ���4B'_:?I�d+�7pn��a�O�nD��ӆ�m�����.,��g{��e����x_b��O6��m�����PHr���Yu�m��r���!]3�ks�;�����OX�H�"ib��BR"���t� +0(�O����_̆���L�x|��ɔ��	��Z�߾wFǧ8F#��v��aE�\��)O���H;�Ҏ�OR�(L\T+Tb�9fe���cD�������?���}�sZ�3ik���C�
;�{�~c8ο����v�忇����*RВjFZ�ç��T�Fb�f�;�Z�Y
PHP�1]��g�o��=pZ����,����bZ��ߴ]V�������ҋ��}@tQy<F�	���C(�.�n���W%iJ�	��% ��d�}N���$���m�f��h�ﬡ��cz��}z��;�X@�f@�@��f4[��[o�E�o�h��?w�Wi����ol�ow��sh3�`p^���VC�?5||����f;�T�D6�=���^�G��#�Op[h-�ι�ō?�-�������T�Id�e��9��)ퟓ� _���~"�I�C�T��.n�JI �-B�d�^��|(�Q�E���1b~ �����ȭ�[~���I��$���m���A��14����K7�~8H`A� b�3�V�}F[{#��������o��������� I#ą)���|�@KI�{y3�d�c����H�eD�����J�Nr����rz�{�wi�`���iS�m�W�r�	PXF���ڈ���X�?�r���;��Y���c���z���x���c��r�k�ƶ�k�`|����noo��`0����|�<88�Yv4��E�4��h4l�#r�I��7��Mq\�J�&�����8�-�.D��z5=p�C���j|H�v\�����l�RA��g��Ȥ�:	����m����R,�?���A�J^���,�K;�A՘N\�Јd,�0�z�	YGMסe�J�Ib��2�LR�������xƀ���`,>*W���4�iRM���!MO�y!�}�倇:IJ��*LkU|�= �X��輐A��uEHƆs#�V#�z\�n{?��W��>���+ƪ6Uݴ�e�4�2.�� Mh^;ָp~c*׭�Z��}=��jT.�'��c�E�.�'�[Gd�?G�I0�@��]�<�}�:���Ԓ8�M;�G��\�Z^z�Ɓ�bE�]�e��p��霎<��o=�;9�s��c��u��������o�ӿ������-����V��>�*0^�	)���,)�=1�&�{4Qmª�S�Ldr��w�a2�<4���tr��c�YZ,���&���cV��LzO�F��i���o�5&� �P}����{?�S���/��/\����>8[ĵ]j(Za�xss�woݺ��믿�sGGG���G�^eǱ�N'���P���3����"������B8�(t�l[��б��D�u��6��q3����ѥ�Gm[�W�b�X)�@=��ۤ �A��KE;�(�^�Z����!��(���p���1��?F���������&W}���Rp�π�B<)�	��g����|�h� ��E�Kp�2��
i�X-�&�t��4d�x��ьNi.)�$PfK�0M3^Ffh�JUA	�w���-�~���D
 ��^���nj�E#ǁoH��k#7}�E \*bZ�++�;�x�R |��qEIG?r���}�ed	m�ե���rF
v{�Vq{�9������!�V�d_�o.��+�>��>wp^�@�-���6>��'��D�\Ttg�>îZ����}>��G�t��O���t��o���M��&���T5}�gm����%{�T
lDف4;!��p�+�_��JG��9��Q�\&��{&�n�<_?9-���[�w��zH>AqJ%> M�d:ľߋ-���~!
�8J��l�>�89���%��$�����x���O���?��u��g�� qmWZ������w��ۿ����~�O�x㍟>88�y�Q�8��n�lù:C)IRc����$e�L����Ɩ��ٲ���C���S��6]�	 f>(,;���L��L��^L�\&��ʾ ��k�T��ՙu�l��$XW�fsO��C��V�&2*��p}l����ňW�uSnc�{߆vuI/⨟]��B�se�I��F�H,]Z� ��iA��D	�G+�K�J/	i��6F+�!d]�����=�!ّ	�;u�,���m����4�:�C��xs����u�RD�(��ot��V��?�v)g����u/mi(��/� F��걣�C%�I@�~mt/���Xp'�=���,��Ts~5"�r-����]�LD�u�')�Mqtq��i{?���;�m�w�Ƙ���� �/��=>|�Z�Ʉ�,�F��(�0|��0�L�t����}@'��/�IN>s�荿��[_6�?;�����o?��o��[������� q"�-(c�0�Hy1�i0�k��� ����7T-�s
&:z9�L
D�x�up��[�=����KW��^z=��F� bqI��������2"�����d=���R��7���޹�Ok{�m���4���Y��?��?������sxx�}||<�Y�0I|��0�<��6��t�\�Ե�����l{c�)��n�29;�nΧ�M#�ڹ�i�A]WUUn�u����Kj[4/�S^���t-��=a��V�����$�D|�����2���4���LP��1(��ajU�IY�ha����Ӝ�D�����y:i5�LS�}�� J�^��=���{����%ύr��T|6�a�.��[�Bj)xTc����(䴹�3p�t2�%M��jTP�C���]�D�voiww�:	��4d�7�1�S�����BPx��D�C~nh��ƍ���A�I� Ci!�nF�uL��#
��c��i������̮Fټ��Bi���H2��֡�ȵ+�1�
)D����s&i�����_�}����}e�C� Mb�@���q�"k2�`]&�m�	���1�M�cPwL�;�]�P*84"(/��X�t�,iu3&4��x{YRy���GG���>>:�f6��4�n~�����������ï�29�_L��w��Y��r@y��k�>�%��5�<A'I8Dף�K��4�jӥZ2 |�	}�G4[0�?�H�?�o�$�e���`��$����z<����^��&���%�Pz�g/���w�yBk{�m�����<<�{���:�u�������_�ggg��e���?�3�(���f�sd��1�2��f?#����D0Ȟ����ڴ�#���Ԓ�t��AL�����r�V����w�q�i�]T<�fP�Ӫ��oN�ۛ�Y��/�|�,�^�P�\������O���� l��J@��� �8W�u�~����6M �T�H
Y��dU���{�~����J��2����nN�-K�rA)"��!_5�##�ҧ���!�":�0���ݡ�^|���N�h� ��ҍ��ˆ�< �#oߠͽ-�FEЏQ�"����̔��$­��Z|!o��ӓ�nC-����D?Z�{�&²9�pLp��r�&��_�(ʙi����]Ns��;0�����*�Q�i�Eɞ�������;��_��Mc���ۘ A#�Ԧ����������m�U�> wB�(������錦G'��h��1�쟑��$�n��4���٧���g��w�C4�Ηo�����K�������r�Y7F���<]�%�/�˿��6����6R��v(��C J���at"֤�4���ۇt�!��T� �:�]���߉*��#�� Q�a�����c��e|�_,�����/}�S_�җ�4��=Ӷ�k���=:�?;����h� Y�)@���^:�L P�����n1�)��l{��'3��s��#G��)Ў}b)��B�:n��
�b$�\���nT�֮M����v|�	��Xt�
��5 �R��vM��I�i%7D�Q!����1��7���7i~6�c��� y&�;��l��᧟��^�w6М5�y;7ƴ����W�ۇtz� q:�&ih�@zdsڻq�6vvi��C���< L]��ɢ{�m)Y8�(�|��]!�D���?�LB[14i�m��K9�&�H���&:�5Xf.E�(0)A{�(Kl	:}tH�]R�(PɐP��W�;�	ϔ$6.z�"n�*��?�+����Z�Q�S,l�qY��(E#t(ib$�JW��ֺ'`_�n��ܴ��u���� �R-$�%@5�އ^��#+̀W���:<���)M��;������>0����ɝ����?�G��_����!��_NO���?}z�S��-K����IZq�~�P3�}�s��-�ۉ��MF9�(�L�S�cC�JĮ����[(v�NO��[%=���=�( ��ZU!4�ӮT�w���߉~�e�A�����5����&�'Y����|�3�����g�� qmϼ [�ՠ�D GttpX~j�8����lA�6A�J�< 'Q���HQBWZ��ۚ���υ�PLWe�k�>7�;�k�^4(����� I�E�JI��S�9��}�yq�o��#�'s��|��-���;��'���zSK
[�b��?V�w���n��aMg4��U������6�-~�I˺k��dB+�@�:@)	��P��U����{t��~}�F�B�}a�~B%���n�S�F䴋�#C�[H��^;���&]}<!�ʑڮ��R���K�m���'�j�sv>خ)[�Jpn����
��(W�#�h�q
�eB�	�F��X��b���i��F�v�@�Y��Ԝ���8 V���Ũ`��%�
���#�Ni. h�IU;hվ8N�O���>?~@��Z��5\� ������ܧ�������w>�8���ӣ��e������\��7*pӨ�!?:����?�
i'�ّ��ry��~�*ʄ$�����]ޡ׾sBoޝ�tjd�
�*�鄏i�˪P�&��y�m�rO��/��=쿇k	�����G���`8���?��Z�3ok������H���%�ٷl��$߂�nja:�6�cU�����:�U�eȯ� �>��&������o�.��G�3��_#R1 �'ZdJ0 ��$��BK��hD[�Mc�{{t�s]���G�{�6���-��"u^$lj!V�s�ƣ����ӹ�żD=C�Q	�$YA_��*J�`M���6<\L�b�$%���Q�b��~Q�IAH<V�+;��-5Y������r1�P7�m��m���(�I�gh5R��Q���.>�X�^xv+�߇}��=��k�4�(]�����'�`4ҪZ��h�"�g��ۗY�a��n��c��R��XDt.�FO�Wx�Q��'"�F;�����P�K_��!eo��iB�V�7�,�ЃA*~,�%�N�4C1��)����TD�����:� U"��K��z~���ɽ�8󇭿�����������W1��]��
�Ū�&�T�B���/��?6��)���)e�P�Ib%3�R[���k2)p�m��IJ�~mB�F� lEMQ)5�/��K#ǶyeF[Ԥ�<c��=�)I��>*�g3��Z��O-�kx0޿u��W���/���[ĵ���Ǖ-6��l������nY&	:���T� �@��V#Kf-p�.���ӌH_RL����j�$�R-gj�Q����!؉;MAJ1@��C��4Z���4��bqQ��+�ӝ�-�{q��Ds� ـ�4�@U"&��i`�E0��S��eks-�E�+�u,y�B1�P��6��v��C)� N�,V!W
�m��BT,|��Q�Z��\i��E=J���"�c�(�MB����/��c"�t�E���H ���&��4�Dh�����c�Q[��R�;>�@b{���f"��"��{�GI�+��{���~�iӺ�=^��&e����<�U|��o��2���MSk!�p�SI�
j�c�V�I�@�� Q�x�6=�e��MG�ڕ"�R�a ^H�HA����i9mhz4���dN��R�w*j�2)�Bt��thp"�\����b����ַ����XE
����>�8����Y��� z�ΰ��9���t�I�m�̋���mj�qo�\��lq%;*��(���K���\��ǧ��ۢy��,��-�<�-Df��J !mpC�2�� ��E41r�(���p�������?�oim	[ĵ�-�1�����7'��?*����Z��lHn�����hW.�IA��z�s���I���-�3O(��*t�F\$Շ��31d�ֱ��O���롩�Os�!�!�;X��T"�sD{��C%<OK��_�)D�L@漌J `�˚i�\��6]K�D���@Vϗ��mCDM�g��/k�n�b��	 �h6�Jo$�e���bp쒼l�H�Σ �J_kxO:թi��D?�S���&.�$�L'���p�$�r~x��Ĉ�`�z��Ed�)�"����B#��Q�݇�/���"����۲N����Q�0�w��L�����Q�ο�D��t,��Oh|��0NWƐ+w�;��m�r�.�ͪ�n�v9Jlm5�� �9��Z��^"�J &%��I�H���s� 1N�.L-~�:���f=ߐ��NJZΚ�D+�$K�������z� (��U~����o<�-�aV3�7����_�Ͼ�Ť>�r�@�����	_�����͑^18���x��}7��݄_�>�cUd"_��o�.�����ڧ��YJ�r��{��c#]f�hW��A]t>��ha��jf|��2"��\���!Mp!,vW�3n��+�~����/<��}$l׶��ol?���w�N�t��WݒvT���FEu��G.D0�[HX\���� v�4˨(�t��HYj B��G(1U�#v��|^޼qc�&��$��P|b\	���ג�E�O�n��F���@Z�-
2�	M�zYI�I�,�ż���
�%��r�t�ɒ�żվ��D�$OH�E��D����t��Jz3Ka�� x:~�𡤈&�dC7��7�xH?���(r���y�J^��4˶���ã��e���3t4�+��2�]��G��;Ǐ?�X�n���0��\�Oɯ�!��D��V�ށs��:�Dx0��	�F~'Kiޯ�J{��պ,�+Io#�N{���RrΉ��^�e�t���IE��[���{v�+{�'�<�ٻ��A�]�pp���-T����K�Y�S���f<�hR>_��dz�l~�����K�������I�����1e`�=� v8�*��Q�v�6)�@��|���b`i044�� �h��,�~�n�Dh�9��S����s�A1(�k$r�-&�e~���y{��0���5;���S����߳���!��2@�UMQ��[b
c�Zb�ҡ֣h=�ٗ�My�[Ȍb�P�4+3z�~M�~픎N�)H1�D���ur�t�>c��� ���  �� "�xtp,ߏ�Sb��_8{3����ɗ�+_��׽�?"��k[[ό�|�¿�Wl?Hg�x6p��=;\V7��Ƿ��ڌ���{�v�j��Mע%�y^z\#������l��ƛ������y^2��&��[���|��/���ǪE�F��\� %����4T��
R{Xo]	x\.*ZV��ypy �-x*���J�4��%.���6|f�Hj�_hVɒ_.iw`ho�a p�HdB�R�˃�T="�K��Hڨ���*'�T�m�i�Wa��z���A"��v�����!x��*n8J���[��x�3�?{od�}�����_�� 	� � )p����-{$��Scҩ��%��)Sr�������S�*W��8VM�8%[V�ؒ�X�e-�Il����}����������nI�@�S�h����{����s��`Ԫ�O.�u�e�e��<�3+�"7����̖+'?�4��^~[kV������*6F�Z���C0���R �nR�fKL��s+vBj����rY��8&ϗ���2^�9M�՝��5�l��(v�8-u�~�����m���d}��*����e���҈3`��D�k;����j��a�� �QVE�G��H��JG���ynj�*�
|
��\��1l�1���\ftm8��4D�e��^$�e,�`�\���	�JD�aY`�3a��~���L�`S��r7M|�����p®���-�3�.�{[Ɉ%R<R>3j##�)�Y��Yݒ� ̥R�.>�ll���>�m>&���� �*w�M\�ҡ�t�Ea\���L~�"�a�i:���,u/@�P�2�?��q;��$��Zj�PZ�98�����+��6�ݶmt��z�T�*�u��߮�+�z�q�{��F����{��l�_�c�e�{}��v��u��{��+��s�h���������\Ym6ۃ&� $nDih� 3�:���A"j���õԴc�kd�"�8�q*�2v�C?�HRC�(Q� ��n��I�n�Dw�jP��+TWf��lacb�E���r�T���nD~�_Z�X������J� ���d�,|���*q"�]~�.y��|_e�{ӿ=Q��VK4��6W���g��2�����f4�u+�m��f���#~����5LT�H���؁��[+f�XH6�(�w�FO�XQ��Id��ھF�bDhà89��O���Ȍ��;?S����T_1�����*����5�7�?f��/�\�93i��3;�(m*�AaL���|aa�zT܆��R9��	J7���7��R����
[h3���tɪ�~
���|Ķ�rI��D�k��rmW:��D�imJ�Ywy[�}�J?`�� �ܜ?�ps�����|?>�D&BLyO�\j.#�B̡;|E����s�xLE���!l{Ђ��9��@�s*|ތ��\�Μ[��Ř�N>>�A�jnI�;FS�K
�(����VkШg��"T��z].o6��*j�Q۵ͧb�u{��M�6}m۶=�Tԛ�
�XTQߢr�����+y��''O���t����I���na��Fn�kj+��=V�%p]gm���q�J�7IT;ڃ��-,C�^E<�+]5O��x�hxؤzJ��]Gc�+����-%a�3�Z�O�
a��,8��5Zq�@�f��E���H��+�n�f�ͺ*��v�`e���KW�m\z�4�.�Wv|���S_ܶ2=u�ge76�8 ȳd�,��(P�Kʇ��M�ۀQ�ư�+7#Q�����&���e���Z����Z+��o�t��g��P��H��K90�����`H���ն��`c�ߗ�=|f���!qޞ�Ϯ��%��W.^9���V��/�9ƶ�gK�yܘ��IyB:#�1�!�G�c��
1Æ�4>ob$*�=
�~�J��c����˟Z�3R�7)8G�D�rV.QL���d����c&����4ּpn�/����A�2{���ꮾ�/�tbLx�\
n �g����!��L�ᗳ��xiD�Ö��3eR�/���R��W�^r�p6���><CǏ/���0�E�5vPg$K���k-�,��4Mc-5�@8t�����b�2Z�s��Y++��,��|:�ÃWn۾��"{��U@,���z衇:�?�Ǹ���g�9�����BB��~�.bj��C咥jڹ�^\$��Y3<�LGE~a~������A̝�s��#-��j�m�=sx�ZZN����te�vl6i��u۳V���)�vLT�mP)�3	��`�`a�7c&�q`�lʣ$��Э28�a���N�	)J[;Vg֮�?�{᛽&'�ON\~���|��b��U��4�ae��bc���;�I��K���l�	��R*�s�2�A&mek6CF>sIJ�*��C�~7�=	n�b�4��MN��2�{��1���ό�q��a��?��������n��;V�V��.<���~0�7U��z�b� �"���k6E?cQ U��<���T�a*_��A�%���c�ğ�SB��6��,�f ���-(��xͭ��0ް������Įl|���-��ќ=���}��.�84r�|y���(�Ni/��5ȭ�Ta�h�"�0�I(�ce�;#5���e�1=>o������&�?ߦ�D���Q�y^K�g�����a^7e��4ULo/��s��w je�SVWW���5묜E�މ�_��hm�4v`��ݗ��7U ���~Dϟ�韎�//��������ϴ��k��kʱ(`�b I�@����ՍkJG �D	(  S�v,Y�ć�o6��	���뢨ES��t��ݼ�N����,����}��A,��T��F��>S���G�`b�����b�b��)mEO(	Z�����/-�^���U������|�������~�S���䕟���z��Le��f6��k[=&Ԙ;DP�?�Pc�I�!�j}_����@�t���T>����T2�!�P <U�ʀV�ub�$ޕ��2@d�mf"��@=��Z������g��ާ����VZ�|�\�a_������'f{�L"�R�>WC���&�L���r���X*$�a�I�y��dP���ہ�7���I�q�2��K�Fc�Nktvnb��ۖ������~d?���3�ju��#n���2�����O��)��
J2�Z�$T�Gf9��3�|	��J$" ��5+&����e�.�t��e�zu�7!꽆P��}!���q����>ߪ�y���p�b�P.@Ԃ�`�ln�7�\r_����j������W���U*�MU@,�����?�p��ů�;w��n�;���Ԅ4�nq���~h w`tR�����=K͎���*ID�r���V-��+k�2y�b�"^�Ν����ڹs�<��@����EV�7�݉k�V��2P�j���р��L��Sރ�������	dܚ�C	~�D�hcq�in}7�>��,%s�>�_Gn{���Iv��wh�����s'���-�aؠ^�$&�~>К���5l���w���I�!̍-O��Q���M8�,�C�� P���MT��LY+��jCB���8*�A��P+����$o�W�C�?�y�=�������Y��}�-�Z�m�WN���Y6���r���7�ĂF<&[Z�r��k~y�1��{��E	Λ��<"�K	ye~_�hcgb�$���G�IyoĐ���y��0���,.�l�/��� f�>w����Y�<���ti��"�1\���l`$>27x�#%ⱡܮ�T�'*�\�Wb$��#TDd8L�Y�{T������K]:sj�V����W�/���R J P�{��:� D=?���q���Yo��q;e�:Ф:�/g��F����o:��C����~�� �E�#\����?������ۭ��'I�&B�9˗���	ӗg��,���8�Y,�.e��E�LA� �X+�����xf.���hthzj�N�i�m�:tۭ5j�Ed���
k�������B��f��pl~^,���Q@���z6R��(-X��=�L��&�Md�l����Y����#�Ky��7�9��#f���DqYx-d�t�D�H<!�vN�.߀��l s8jP�P��\���`��f�T���I�m��?T� *OZ)t����+"�J�������О?������kC�!�?����(	>~uq~��$��I$�ox�sB�K� Oj�t�q�Z�@��$�a �?0@!0�1�0��gQ�I�S��v;�c~� ~�̭��KG�TT����3��̲''�ᘾO5���Z�:���mk�
)o$s�&��Rvq()/�y|+U������ac�7���7���L6?*�Q�E�K�(]�H���)�x��Ǚ�EY(�* v�����E���Ģl���D���h�y��@��� Z@�g����|^�\�������M�y�;~l��6����xU Ģ���}�C��k����wA���� 92�N���f�j���Mq5����"� +7ō� Q��J��c{��kw}ryu��~�Хk>�zl���R��N���{��`m�ǘ�;���Y��	��x�j�X��`�ēڔ�<��D3
ue���ce������vҜ�c��8O�k>{�cg�F��K�|�g殜o%��m�{�ZP!�Me�M��[]�\���6��s���¯˭�6���%����)��lI�����)7�̧=:UܜbZ�uH6f��Q����jc�]��p��#���?���)c�#�����j/�.O=]����}�e;�%�6P�Ñ��E�GjnP�a�� $�g ��b��{��9�ȟk�ߥ
�S�R�$�	��Ƿ��3�I�ߙ����Y��[�'/�k�ൃ|������c���?�g���>�5/��_�L�_�����1�m� ��L\ʛ��E���;�[��[���{ �|}n�<-ĕ�M��)ө3Kt��<--�QY" �p.;y��8�d�'i@�����z�ިڲFoq�(���6���c�h4�������r)\7����];��P7.E�p� �Eu���?x����c���V�.�t
��.���@3Z�D�0�X*"M���}�ϦYV6&Z�張���*�63:zb���P�Ϧu2����Ϡ��c"��sCi~\ �jPcȒh5�k��#&���P��ax*�j呇�;�:Bl_�3Ù���_nO�^\^�7'��u����8$����*��%��G�V�4��D�6��(��
QJ��"Qn��eJ��b[I��$�%B�ʘ[S��KƼ�����Է�sn�˱��N�=�#��nle��_|�Tg�7��;�ܭ��Y`Am_�e峁�J^�lC�`�{�(�[���Ǽ&XD vC��2��b�yUSY� ����p�*��V��ڴ���zs���3�g��q5��0\ ��S�������p���k�j���s�{�RE?iQ�2c��O�bP�aP��
s�lo�3 �H
Ӑ�+B����d0�t�R���t��<ML�����'ch	���~���T7_����֛�(��� ��0�=�����H>�n�#�|��y�so�����r���Թ�E�hT�*�(��O}njj���Y'&ع�Y���j�����K+��R����P3c��J�*�mAdk��Rc�4\�R�ŧ�m�L�f���~�сA~�����<�-�Vx1c6���rd�n�ͨ�:aɔ�- ��6�c ��Lf�w��i��pk��/F�_��t��'5��R:R��Ĺ�-��Q�Z��R�#*���?b�����h;F�v��ZQ1�*w3���O�j^�blh���?�wֈ`�/��J�:��v�l}�ߌ����c?�o߮_Z��O{��5Ԛ�@�������E"��T�E�j��q� n�(b��(*����*�-�}cp����X�ff�s�Y��$#���ݍ����mKW.>�|�3P����= ���O�M_}�V���*�7��a"c0j�1�lc)��nD^٠Z�C}����4�j���*�kX&%I(/fU�v�l�t����\���љ�K�܂���7�s����vI��8���L�ʪJ3����<��:k� ׵�ݵ�$�&���5�Q�����8/�yǞS###Erʛ�
�XTQ7@=��c����0�8w�왳����_o�[o��M�
E,�D�?c�9Cؼ� me�M�+�e)T�i�'HɌUJ�,ђQ�/�S���vl�L�F�-�^Ցc���4C���b	)M#�6��Y�n	�(
��V@s�!�|��l�\.)�
6 06C��B/�VG���^�s�[ ��DD 1D&���FQ,�����p�Y@�0o!��8�O��,�dZ�J1mWچx3D�s�lg~d�ݸ6mTn�\��[>]�3>t�o���὿9�n�3��n�4����ӎo��Kn z1�l@��F�*�G��'��$�i��"-�M>���k���;�Hf�Ò�vު���gؖ(z�L����3��N�m�ʩ'�89��2]b����g/|���������!7I����+�{���8%B޸������S��򻔪�<��~�y��T��C��J�x��$��e�VK;���tu�K�Sa�
Ú!����Փ�_+����,U�r��P�s µM���!�y��iii�VVVd�(�h�7��*��L�(�lټy����~�ᇿ�E�XU Ģ��Aꎽ{�=s��Ξ��ܪ�E$��e��sI�k�z�5+gD�aA7sCm�����,Xc��F���°MN�ҹs>�?�eP1@��O�֬�����?')$6�����Rn	�ͬlQ�+�TX<���}հ�R�f>��Y�TL��R	ql��`�"#XN�'C�.��A����T���.�b^V:��A����!Xa�H� �:q5cyX0N��#�Ma�E��̮���Ɔ�5j�vո���0fâl>�ą����W��-���wU�jF����8�����k�f�T
\5
�cL�,� ���=��a�W�c��	c�Ɔ�`�$)o��цbr���h��hu~��ą��Sg��ߝ����̼�S��ވ'w�i�6!>�3��7od,�������˗=W6^�����
R�D���L��1��n��t��=:��$M�&Ԏ,
p�a��)b5eInu�d��U,cH��s0�_��t��NSQ
hW !@��z,�{`�Frnn@3پc���w�������� U�R�}�{����W^|� �u������^[��9탈�A��B�+���}u���;Z(@�I���-�zΟ�*�_�Kz��m\wm^��W�[㛇��M�ś�bdAS-J�̋_#�F�
Ȋ��� �*�"b��A#���LE�adjfFږ��"T���#���lM%��4��h`ԡR����2��x��P�$�;'!M������0�ʬ���A`01HͺT]Ii�+��;�bx�_����r�5ny_�p���|���T��X�eV�%Pc�l����������1;h�l"D�&�
S����چ��Tj�-��P�b�Ԭ�-��ɬ�D}�J4c����vᎋ�Ǒ������3��x���~��\�]���p��R����c"��s�訃Q�)��j�C�A>�*�q�������j�(�JK����uJ�����l�Y��N���H��A�:%S�R�-�c%&�B��ı并r,0(G�Z�$c�B�O��3�q`����O���Y�lq�>�m�H��924���{�>q�CTԛ�
�XTQ7H��ٷo�����'N�>y����v��e����}���4� �y�`�6���� �ĩYX��b��HS_~�ϧ�<�����J�^�͛����8r3u����7X�"�I�J�Ğ�a��0ӎd-7LH�X��F����#&ɰLA�G�`γ"ie"�O<�DZ�L�u������;�HZ� p^���M�D����#�=�Ej� 52ami��L��bh1J*s� ,`q�69%[b�����98E��'���W��?;з��m����[~a����K��|_g�� �+��]�ʲHL�Sa��W��o2Rf �Y�ݘ-����oh ���~����#�dS��f|���3�( ���4*qki�앋;��ǧ��o����l��Փ�<�t��_��ﱳnI�?���U���d�3xP��ѕ��U�[f��*E�A*>6Mq��2	d� Ά� �p�~>>����.�����>Ò��x��F9J�<�YF;��1wY��_�f�q�ծ{O���Nh%�|��:wh^�ڨ�d�g�}�V�2��~���o���ysW�*��G}�3{mv��+Wƣpf�[r*����,	0X4�8h�\,���/ԩy�:_lH �xTkt�@�(xmi�!�5����U=7~p���R_m�,�+b�8labQ���a��Pڋ�2?�*WI����#j���cV*)[^����?���j���c���k�ڛ��~�����On��Á1��FS*�ebt���L�K*srb�#��	(40����vG 9�OU�̔����y��=���|�<����T�}��m����{�ϥ�����<�~y��/fY�f׈0��� �
�K�=7WE�����_*�h8��$b������G�uH�,C�)��Cf	�2S[��-�2è�}n��=�ӯ�Uߒ��f��];��;�.�𯻋����54���d\ -e���rIfP���f{�z�Cf����̠m�(t��oL�����(B0XV�k]�l�K�t�B��]�o�#h�6U�}�k3k+���nR�x�^'|�aD+��m����=��?��W"6c �M���h #���m��g�{��={�t��7u ���n����s�]yꅧ����tW7��
_D��D����>�Z����t`�.U�o�^�o�J�8�5��b�N.0�C����-u��W���&�|�5�.�e�1����"ԓ�)�I+Wl9\;O%QC���R��E����oDWDшj�����25?	��X���b"->��ص���q7ZԿΠ�D���<_-��~���-U�L�'�Z��y\�jsG$����}k���/և�|zh�_����7�=��ߜ���~r�,��g}`سG�bb�)h������C��� \�������w\'��x	� ��Ɣ��,b壨@����7+��������A8�6�7����+WO=��ŋ/�Zg���ms���lB��'9�I	A����Ƥ<0M�뷨��c�ě''p�G m,mrv�2���R�4B�+:rx�^=<Ks�u�q�Y0����W��<VɅ�9�YXGDP �2n!�ו̽��b�P'�����u����W����={���]�.��͛�
�XTQ7X���oo>p��N���؉c��i�@�6��v8�E�jG��`_B?R����a���N���ti����,[�U��uĈ�)�dVpf~��_��j%���0�VȭT)�@}ɋi�f�p<&^��ϕa����Ⱥ2���vF�Q �|&�p-G|��I8� �T��&��-IX��ŲR񨁔�lL�܈��L�}2$_�4 ���Ԡ���&���#aD��K����D�����]��߼�Pc����Fl��wʲ}�Ɋ�*��mFp��$Z�ȼ`������DT*ܫػ��D@>c8�1�C{�I��gR�� ��P���& sY�泇�(�<p��ya����Q������_S��'K'O?��ҕ��Z<�����9n,�f��$S�����d,�ljuS6/}$�ܙ i+O�LYCE�O���'�f1c�\�l�"��N�ҁ�)�r-��TM���,e�)K.y$�b?�&�p�s�0=����-���p$��E(����1��{�����C��e��oٹ�+�����â� �Eu�v���㓯=�����ᅤ��=���5H�v7�9�^g�փ~�G1��AkOE�J�YEm��g� $�-3�sy!lӹ�-�Uh�V�w84P�#�n� 4<j[��u	s�0�9�8ؠlN�t�@J%l'�δ<��$�m���*�/1�SGT���h��XF�~��"�����®�;&Rfϔ�Z��(fR�5��H�/V����qήn���>=\�{���>~���7j�cI6>~*�������Y�q�a��4����� ����x������E+mf�d�64�O%C,c0+����C���mlZ ˡ�OI}�Vf���M �[�N�������/�{�ҁwgN<4�,T+H��<��#rK6�z��_�S��Q����K��e!I �̐b�ꀦ~�8`A7&j!�o���E� ]�0���y:~b���
�`m�tT*W�Q�˛(�ӥ��K��)#@����랧��r,PB�^�+�{�;	�H_�=����y�����#�}�G�X���
�XTQ7`�ݻ�{�m�|���Ο?���:�Jh'�>��/:j�_]Y��T�5%X�s�GK6��U��Ab��5N��Qn����$�6X�H�%rj�ԉ:|z�/LR�����ͫ�]���
�P�i�D}��K���b������| �Q�Rw	�d�A�K�05�LMվ�����P*k�9:�.5F n����3�Ŝ�@���`�S����s
��?$*�oA�[[S� g,il��:��_�[wϧ�o��Be�ʌa��Mі3�7ʎ�;p>��畩�vg��;Ӥ�	�H(�1������́
ױ���C�-,���3�/�U��U|0�DAbS|:��l*Q2�mG�&�bn�^9�m��3藮�}2�uNO}���^}��S����L��B�_o$����6OI��IG���Q*��:�����P�cA����9	�5�SY�2kX}�}�&gk�z�P��J��eigC�������� ��' ��(��Xw0��c�d�{��H�O�6��ǹ�e�Sp��0�*�����X �}��o��M7�t��;�9���עޜU Ģ��;��~���������f���tw�e�Zd�}���`�i�L�x���$�$�H��5�D�� %Z�W��E˛(fM�bl��E6L����t��
X4�?L۷l`|�@��$�C�00��jYg&�n���s\�$	["��Ӏ|^���DV�P�tx�e`
Q@�@b"��Xf��ZLC,j��K��W��R�9�:��.���ʁhB۳8�+�<h͉V�XF���	���s���3���te��7��Mvu����a�Q	W���ʚ���R�$��V7gUk^�ܡ��.�y20��2,"��J�;�0Ig���f!v�L+��À�6���^����+���Ϡ��O>Y:;���v��n.�z��潪�\�P�N���R	9�i��vG����-�PY�Ʀ$��b�M�B �7̳͓|��Ƽ o��QZ\.ӑ�4��]�B�^��O1����T�����4d>󵦡 v�v&�Q�׉� �t�:  �u�n3�6J���o�18v��7?s�w�PQE�U Ģ��A�������'O��wb��:�c߯g�̬�2J���Au,,:��5,&�Y����Z����L+��,��A5���"�er�45eс�42�R�6B#�2݈\3���K�J�v#���Hl�@eB<�ѕ댬Cs�*u��d>��Fm�!0�OH�Q������~�G�Cyځ�.�MQ�b2M�[��l�0��(�MI`�?q`��p��\�T��O������9����ތel~����גQi�1�'�|��\%�����Q&�,�Z)
3apm�` �1@4�H�T&���m2(��fh�\^&���8B�<m��Q�=?������Jwer����ۅ�������_�W�����U�T6� '��;��Tr��9|L(%s����_C��M����'�>�F�H��Eq%��v�C	c��@�Y��1Lg�wi��+t��,-5�������|t�����5���9Ԟ�W����@O��܅0�et
 ��' 1OHY�P9����Ykpp�՝;w�)�)E�V�*��ݻw�E�J���wii�n����*�@�f�Y6�t^������1|XDz�a��9Ş�Ў��
�h!'6
D| �õ�bs��=�������Ѧ�rl<�/&י,I ���6�%����3��D�u��8d����'N@�<mZ�ť�@DN5"ӆ�"/�h%C� }�r�L��q�"��^~ h�»�p=J�,�2�1K[����������`8�[�f/�_lO���������m^|��V���3̔�@G�ph�t.|&h�[�Pr�M�����Q�Ϣ�g0�PWѐ�0��BQ�g).�*1"͒h]8�_^mM�sγǥMi��߀f� з5� ��D��H@	x���VCjX��1bQ�������2v���B@���llKS?Vb����K��`�����o��|"I,�e;s9q�i&R3��c��������z"���s��FP�+j�)��u3����[�n}��DE�S@,���~�a������O�y�ĭQ����R�D=�(�|;0	zNI�K�j�Q
���Ik���]fD��`�O�y�6���ұSKܖ�V�Z�Am:�F�@Ydȼ����)/�q������^�$��s]!͐O�Ř�~�g#��٘�X�Qy�'�IJ�$��P,C�	��X�`��Rh�I��M"���r�8�����	�Ie�(o�rc���m쭵��7
����3H\����1����ǃ��n/�1� ��I"`%5��D͢&yB�߅� �S�Yrr�����M���JL�҄�:�R���F܁&iP�m��--m;S~�>������M
�ROQw7,U�C�0��F������*��)	>8pEdc��5��`!~o��]ap�z��y�6�8�Qף z�����t,&J�����_�){=���q������ �Q큪�Gtf3����M��ڹs���{���� U�^�w�^��֝�,..>0??�v^$Jz!qzf��]�X,�p $��u�M�Q/:�z��zD��uK�	Zb�m��3�J���F�2�AK+;ޡ��r��[n�htp���yJ�$��!�hU柭��k ��6����<�Gm~���/���2c��itc�#�E_Z���H�02��"m��$؁(3s�j6Q����򨕕[��~ix�'������=ME}��{ti�������:W�m�5y[�1SL���T�l��i6�H�W%�/` �9X��}���j���k�(�#9<L�QNHͅ�
��ql>.]����dA&v0&-�=��yC�*|,���.�=t�����zWE0��e��p+��`�1�+���Pr���`�T�#���&fK�ʡ9z��	�4Q��:�1�<i��|��<�s����wl�t'@o��\q���C@���;��UD��+�5�[>׃6�r�w���?���}��*��
�XTQ7x�{�Ѿ}��/..}����t:�1^(L��¢��B�`�LS>̎�cq���.Xb��/L�ؠ���2�"�iU�R��oˬ�D����2xi��n��w6�rw��;Sn4��Q��Y��F�2� ���ZL#c��,�nB3X������[*4�ѥj@Vِ�����ah�v>*����S$6�
��Z8�J+2�~�o�����w��y;*ꛖ�H�f����)��+�^��A�r�I,*Ɋ��@%�%	��! )$`��L6����IjA��j(�1Z�������}��e�Jh�����P g��`����6�R��Ie{��!o.�<��Q���r���l� U��L* 1ØZ���`���[)3���)��/�K/-��s򣊘i#��7�jo�,��Ĺ�M�{�{|W��k������ܡ���s�~�����
�U�Ѹt�]w}��8Y���� �E��G}t��ѣ_�x��}�x��"a��U�2mf-\�Z-Y�^�Xh��z_�����y�����f���i�S���ˋh���~J��4�uh`�G���t�����b�+{�[ʨ�ˁ��ISy����dh���C+�r�1�2j(H�� ���$ ��w$ET*�9+�2�d��"
��4FF�H��]~���qy?����c2�>����ܡ_t��f+m[����/�V��V�Bl^*,bD!?���B2��	�xc��0�[U� ��l`���(�-�͍)#:�A�+(Τ\d�W`�!ꑲ ��j͢�Q��68T"5sh���y�	� ����  ��,s<*W7R����V�g���-�Zd�*�(��Պ8�P �p��/���`�5s�7j�$�'��NM����2�ױ@��z���Y޸q��18��c���9�E�� �E�(0���;v����MLL��}�V^0,0hg�M�����0� ����}{={����,VM=�VQE,����[����D*���-.�ӫG;48P�qi��N%�)Y.Z��$ZHn3D`�`�h�
�� ����~�ģj�����ؖ���p��,_�͐�N*�� �����(�hď��D D��=��;���Ф�#��]����f�O~����y�_���M�k%�P��S��LO�H`'��:0@Y*��7��P�
^��!��a���YN��D���9"���H�I��$u=D$Fl�$y�hq�?@4:V���&U������yb��L�<�T�����|��>#�Pn�JZ���:�:ݡg����Ǜ����F�"�y̹��O�z2��R�0�Z{��b0�(ER{r��q�6�e���s�PX�)Ъe=.��>ףm۶���w������>���SQE}�* bQE�A�������S�?��C���&���\*��)� j;=�����a�^��L��9\nH�:e{���4��1��� 5��ԬE/Z��� ��Ry�i�K�-H�9u�bAK=^K�6b�R/��e^x]�wC$Y JT?��E�Vi+0#��E���i�f��~�Fڽk�3���҉�|�b��(I[��ϵù�91���������F�U�4#��-"xd²���؈��ˊdv�-�k.�j z���"1w:��T��Y,1���汑ʧH�/%�������K"F�X.��1x
��,V{��$�c�)�d�S]��z
�:�I�<;A�-��r�oWe@��i��*��I��0�@�k���� Em���G?P�����
:}����DXT�������~��F��RԷ� U��6n�8������Ç�n6����m���JZV��C��C�b�)�a0#XL!�P@�������������BX���Y2�%��Y��4h.Ġ���A������K�s__?/�>?GGr��$2��͕���3X�<,ֱ��!2��H�I�����H�o+���r|U��Xkg��??$f�К
��ʺ���������ioǇ/�w^�qo��}�9����g~<�f�G]�LJ,����[���3������b�6��bTJ��tS�[�����T�%�7�;�1f1`�fs��O2�|�'$-~�@��`D�nvh`cL�#�a ����>����8ͣ�H��q.@����7P+�g3z��E����J)�.Ê^#8�8G�X���<۰�r�����@��.6�mm�*B\�c��8H�<��/�����Ν;�|����ڢ�e ����@��c������iv��ӧ7'Q�A��`�PsM1���*F� ݆�3��AԋJg0�V�Z�`�����(S�)�AC}7�L"�K&L����h��
9P��R���*��}�(1B~�P�
xl`�>��I<&uo�b��Q3/Uu��ER
nn�F��$S�33��4K�Ni��1�7f��A$#���]8�x�]�\^�����}G��i�a��/Ȯ��Á��R�� ��z5��C$�dz8��-�1���eI+�qR�x����C�W4f^�ɱ�j	�d��=K���Ƿ�Ci��JL�6{4�š>�� "a��3&��fQM�Z�D�#�e�QɎ����������-z��Y:��"��!_�� ��A(��.�߫Ï/)}�B�F�7���^�;�&�Y�Zh���0��i���F��I~��9w��w���~w���m� �E��_��_^9v�ا���6�/e\.3Uy沰0a��h�ػ�z[�`R�,7�e��4�{� Q�°3�'�Ĩ:�#�L���Th��Ы':DnHa2@{���A^<m�ɲ,�I��؈-i�
GiA��6`*�j��f�"�,���e��U2yI�����f[�R|WWXE�)���B�d�N7��,��|]�������|~p�O�CFE}�26?��.>�b�����a{�����6��m�R���T��E~u������L���*�h����� tD=/�j�5�X��(�]��ß�[���z�Mm���=?W��	/Q����,��
�p���|���n0&?XG�N���s�t���1��T�9�I�\��4C�`,@϶�܇���`��Yېi#ky��>�i��ub��<��U�^�}����J��066��w��]_��UԷ� U���}��'�,..�����*w��=�N`��_C=�t=�+�:6#|u=AD�ڱb[��4SZ�J]���ʄ֗+s\X�1��e��ivi�^>��^_:D�Һa�VBq� V�ۙ�ӔP������-����QA���D�u7CT�	�6+�+x�`v25��mBeL�"���i��I�zg���{��|�l~�}�/�R������o[��������k��U?�����}U��V��Q�r-~[1^�L�D%ڀ�����U$"]�݊��XlRRaϔh
)=q��O�'�@X��;+�~�E��6Y�"+�cְ�&C�Q��=~^6-�&���[�rm3��T��唾��I:xd�&�1�Z����� ��n�eP�Ȍ���pU�^BA�����Έ^�b���%7=���w|j[y��s��Uݣfn�[���]�v}������RQE}�* bQE����?�я�r�ʧN�9��o�Gu�6��B�jqA�
��W^;(����F^�#Q3��d�E>U~�P�S*d(TӸ.�ty"$����H��?A>����*9��,�B}�=6:d��b�&`����Hb���KA�Ir�A�ږC��RX�N*Y�2�+�.�1ev{EI�0l�_�˯9��g��0��H�w]ό�I���Y��Y>v��+�1vd���Z���em��H';��WÎiL���bw���"���!�][l��(3i,�v�6R*������*lg�����2�":]��c�d��6��7�T�˽P���ʦ�4�2e�����VE��d�2�H^�V�;դg^\���-����B�k�P�rlrH��%D<���V.�(T��^k)�*s�d����:O ������^T�,`p��޽{��8Qx��V�*�Z�?�x�w~�w>==3��f��n$�h�=����w�g\�6Fi6Q�^����0}}N3�ֲ�Q#�a0�T�f�$"�$�%��[�8���R�Z�9E���w{4�i��%Jl��v5��TӦR�b�W�+T��9��"�����)��i)o��|U�p�ڼ`�K��F�V�� RJl��1ZM��]Qgv[su�'����_��^׸�e�4��oZ2�x�c_Mڗ�la��;98.L��B$�� �/mG�`[o1J�)U�1��-�m���2����H"���4�ޠ�&m�Q�u[JT�(��|섢|�$��z����^�]�	,o��p��_L���詧g��D�b��*Wf !����r�����ދ���RH�)�=5����mj��)����!6~�s��<�U0k;�ܒ*���v���������t@E�V�*�\�>��/}鉿�T�M�����WC܅X_`�
-�(�eqVQ&�U�0�����k�D�z���d��
�&�'�R�0��ؔ�D4�,DJ�0~ݘ�V��/�E�ʨ��N�VZ�jR/�j�Ao��a���2�ђ��%Ca��A*�|�L�6�j�Z��YdvM���D̳�i2eF-��e��(��L�j%�V3��@� �Mf4�L�[$�ð��f�Y�ߋ�wE�3��,�W����kO>�ž�{��wN-�G
���M��MM<�+GV�^}O�3%9�$��X�GA@��\�(�,��ܥND�A�/Q7����DY�̧J-��MD�n�h�*��� �K~�%�#1_�p%HWd|��T4fWa�d�?� ����9�Aj�}t��O�=7A/�Ԣk0����!�Q��� Z�۔��l�9�5����� v�8����\�0F���x����C�k����h1�y�^�{ H~����۷��O��O���*U�wQ@,��7pa�#��^z�Ł3gO�Im�Ɛ�`��@E�8iq�Nk�s˗��D�T�1k(�E#��0?<A2하ɂ�%_��re��gP*���7�x!���y�a�%�������-u�*�z^8M/n��UM	N�7�A�b�$���l��� ��\���w#@��1θ'Z���F�J��_E��ʾD�<�̤YK�}g�n���.�07y�W/���A{ݎ�cc���R�ٹ���M��aw�̠ʱ�2�
���d�26D2���� s�)y��%��9�{�<�l�K%�L���ɦ�-)T
�O1ü*�yV0�z��fTsw�yG����P�� -���Sz��:|�I3���J�e!UŲ׎�(�d�Q\�;fc{�_�/ǐ�Fe�c��)j�Q�j?C�*j�6��K>k���C���nݺ�|��/����SQE}�U Ģ�z�����������?LNM�==9�����@�,T�����j�-T��1��5�JFk�P\z��T�W���~�?���p���p ���
6hf1�V�K>#�vs�<�N[�|�Y�fv��?�j1��G�%���:��
U"��r��p�Ϳ[ˠ����rua]���cc���fs��̌)m��5��'��*et 5��d��[��;L��?O�����m_�8���҉�x����9��ތ`1�Ɲ�KW�������h͟�+��Ӳ���2_qS"`�T@[��F1

�vJ����
U���r�y���`p�Mu�Cd�6�f��)3����c#�R� �`��s �%�K$�>�06y�Ԡ�9��k�s/,��+M�]4�eǜ*@�c;k�>����>��<��M���}��6�V�Y&ׁ=�f�:��)���k�m�<�M�ŭ[���<p3�TTQ�e ��������}��]:~����������J���^�<hK�`  aqZ��A��g3ʾ���M^�K�V)ϒ�ǋ?/�fB?ӫ�X�����U~�1ľo�6m�Q�i����4P,�%i�d傽��2Z�k������ �MiO|�o�b��Vbfb�b�%��G`��V�������T\[j*�\gf�(q���o��PbXo��{:��ts��������6�?��^�Ѣ�Q�C�U4�eO�43�f�W/}�v�,���y3��JF]#��R�M5�I����0�<���F;*�L�H�9;��Ae�=:Z�uc����Ɛ���c�4T�TY��#%� ��:61z�e�_�f�����Uz��U:~<���ߍ�O��2��\omnW<m0�g�����̡X�د�<i��4�C�'�!=�\jAJ�s��c��ܹ������?��?��m*��D �����?��?>4=9��kW�yE���1@f�k�Ɖ��LW���>�+�o���3�����2*0����V檙0k2z������S:}��׭R��у������V(����B)��%�����I;Y�Y��fR�d�sc���]�:�|so�o0�	U������B�v��U�����(���S��u՜��+��Ԃ��fc��}���ɕ���������r����}�֗�Z4v�nEK���	�J�˳��×����Qw��Nw�����}aw�6+]q���PW�x��
�̂Jz�r�M�(�C���(m�bkS�0 +��OՑ��6�T��ꍌ*}���:�+3�2�a��]Z�i(s�RX$�%�l��(Q'���� ���E�;t�O���a�U���=�w[�-6>i��V��׏s�7����%�Ғ��5������ &��`�:ܦ�v�_���-e�vκ�nspp�������{�ᇯQQE�#� �E�&����.]��3O}m˵���x�YoZ����n�i�C����a/�A��l��Q���@�f9�ݎ��E�-�����&$�ɰ��R;����6u��ԅ�]<D;w6h���u�q	ڔ��x~8���N^V�ڕ����Ƿ�uq�w^�NF�E,��!v8�rb)a�%Q�T�2s��$�ԷB4J��!�4�_0���[����O3�Sm��^8a;�//���έ��:�ߦ��M�Je�nz(�Q��C�x�\)�su�$�S��灰53�7g7�����n�ݕ%����h��2V�5�������x��H��Ŝ2H!�b�|��r�eNe��N��WK�Z�M9#��c� �-Rz `�����|��T�M% ������q�/]N���6=��2����"tT�a�p���i��2?V���)���T �^��k�����26��f	�]M�zB�z]#��1��������zT��ˣ;v���w�����E}/U Ģ�z�Z�����V�A��Օ�O��R7�<I�ș����F���J�5���@���xę�!p�TFt
��0=X@]��H�.]]�(hS����R�D�>y/�%S�d1!-��"S)�����2�6-&�<,٩����AaŢn;%��
��fI��W@� ��}Kb�c�8/�,.̼�O��i�9e �� g�egT���4�l
�}[�(53�<畆�{}����NWϿxa����U�U�F|r���e̲}]s�k�.�z��*-�W�'��?�2{v{ڙ��Wn���&;���7�n��/MB1��E0":�a��=�X����|�$Ry���%�;U��jC1���9e�R%�R�?��P��RE4%��Y�qC�_ƛ9�p�8򩑧�k��ie��._q饗;4~��ǜA�-�"�Q`Ʉ��T��	<c�����x����uJ�u�ލp�%I��hp����i��A�$��� �P>��1��ʭ����|��Gy�CE�=T�*�MT`���w��䕿>y��X%��Q������}��^q��g{�W��YF�{� 2��'�H��X�lC)���*����2��7i�ӦV���[��>�*U0P0��(�l"a�0�h�⏈3y�fV2[D,H���-�l
Xm7�?2E`}RY��-��i��6~�)�{�X2�N�L��
�m (�2�D	3lm��I2c N��017�V�o�._�g���E��v��w�p�K�Yi�ni�\�Ϟ��G&j��9��~�r����Mu~u{��v�1UGO�t��rhy]�YY�V��N%�N���}�O�_����$
ki�eq<jg�1;ZX�v�kq��,u�}C $��:5#�J�37�3O%O��:6"0h�ۓ�D�7��s�r���7�R_�M��V=�X;w2�(�yɚE���8�AH�?ihH48lk�����y����+t�xF���;z|l�T����$�Ź����PިJ0���-bak0�k4��HSѪd��1s�������q5��~�h1�u)�g�Z�~��;���֭[�����* bQE��
f���?|1�-'�����έ�N �(0�~��3�ՠ#��َ�W�Z���ի���eQ�����!� c�$F��e�%ө�߉he�M�1���eZ\��[��ؘI���Bƚ�ڑ��(5%J@�)`���QD�8��+��T~>އ9e[Xİ;�n3��R1j�{F��LHy%�B��
%k�����w1G�y��xT��B�o3 �F�K����| 3�yٱi���֖˥�ԲS����[^�0�M�����_���ڶaD|���/غ4KLS�ٌ�F���⸧>���j�__9I�
��5?h��~��`p 
�I��%Mw*��,�L�i�4�Ȱ4�Ŏα�XJ)�$k��Ĥ�gm���q B	�|� �'1���b�z�խT�s��gQ�^�U�HG�w�3$���Z��H]�^�2B$�x�h�"M��խ�`��&\zy|���C:q:��9���"��F`>uf2�lD�c�X��V$3\>"1�.����� ��ܵ�?�ǐ�y��M��.F��
�f D���gq{�ʡ���ʕ++,�۳g�'�}��v����* bQE�	���������������׮]�K|�?K��Xk�P�/�nAkƱ7K�1��@���g��,�{�]ߖa���o��c�:�;�s�Z����dsW�"Ej�6j��dlI��³�L`&��/@� #�XJ<X�$��L�������x�y6��Ƕ�8q$Y�Z��M���f���m�9�w���,J�G����pQ�uo��K}�{���غ>��K97HQ�B'�����%X�/���sP_h�����9;.�����E��񸭈�A'j��.��[�*ŏ�,'�dυ�z��)��Dq�2I,�-�v݃v�-\(�Y.T��t;�p{6��}_>�f13+9�f����f=�H�u����ft�D��B�u��:���b�H��Q3�%��gĲ�o�u����A�,�2s��{xv�/�dI1�4�m�b�eH Ө@��B�@.H8��}�3c�N��F�����dr�1Y�{%�vI\zH"�؈��0�:٪�D�MY�<$�>TG
04���D$�R�w���w��-�3CyH-1$"N���7FJ�'�q��!!�P��86т���/����"��+�y��a���)w=�H �5������P�<8Ƀ}.�b�.ʿ)�HOtz0�h��|ҭ_$о����%�L���z=C��ؼy�O.������;�|V�o� *�AP*��G=q���o���5gϝ�NV+�9����&2��ްb�!��b7��y%Aㅼ��2��5e�p�0a�P�V�C[���ð��`�9�����4�̹q���*\����6~�pg��R{_J_F�!~��q�ٔ3OG���%��(;eo�B9D�Ъ�k��(֑d���E�c��
�t5��oM�};"�!x�d��[��wK\͙��# �y��yI�q�Q'�!2�&^h�EYo��,��D׼���Kq�He�Ĝ.���	M�m��E>>+�tM�!�]�M5�L�Ɛ�&-�5{a
K��cK��7M2��!�&xa%�eca/+Ci�l�!t���/q�Q93Im�OA���
̃HLf�F,V���ٹ�^�Þ���u8}
ۆ1E�K����p��"+�����DO�D�u��������]����Bz%�'�-���I�Z��n�<mOik��
���j�Z���^w�u��m����g>�(o� *�Q�y�>�'��z�������$U����&����LP���p�F��g=EilDVp��
8%�4�$+�?É;jUazf��4`�|�gG`�*\qyV,ˠPZĽP挻����]3#�0�#�cVB�|!I���Ma� ����"4�"h#A\:����X둄�3ɂ�g:��R�]&�0��m#�r*ִ�#�=�PC���߳.��,�膎�f��̌��Ǐ��h�'c/j$0)p�&���8֚���,�I�a��M���̐�nڜz,�n�iHq�ޔ�]�I?s=�7�M�ыq�cN�I��)\��2��*U�-�<�.	�󃃵��qI:��Ӭc�4S�=�ȟ����=�Kx���Bs��h����ç����<|p��J]��c��5-�'��./�͸�kM�%.QB�HͮD���}"�C�t2r}H�{({������(eŊ�Dr���?�y�xC�Q�x����������������hG��$]�
�<Qj��2��b���̳���m�����F6 DИg�VNIy�R���.�,n R�^���(�2��Jh���߄���L,��
p��e�iC��5�7�˴��ݰ�X$f�C0��3��F<c�����O9���yx	R�����+�Hj�H�ԗ�7L;���c�������DR|�u��̗�:DJ�v|&9TH�Y����Q�nԑ�43!�V���d`�{m��F�q��(爖g�`��dC��5|�Q���J5 mR	{Fmn���%�!�и�0)�lZ6ˬ)6]yQE-���2T��P��b�r����g[r���g�J����$s����E-��+�5%�p@c�#9���p�\����:��86Q�ťܐ�8&A1�Bj��st��B���HE�E��^��mHD]��D�h�( �=�/�?D)r����(Z�l"���GNi��Q�ϧ7o��77�|�7?����!A�⍄D��=JK=��O.,,���C�Gqr�'��&����n�O�8�J�ˍJ��`P�7--��
c�4���Rs�R�`Mٲ������x"%�	��A�7T*�W�@���p��Ku�>߁��mعs�l�KV�A�Z��	�MS&Y��$���Z����dƤ�g��M�&��	K�@��2�� )l�|��3h�<�v=A���H8�DĔ�D=���B"?V	�!������U'�m�v��-�#�HL���"zJ�L���ŘBv;�E�T/�yl�mܞp?j/3�C��6���ث05C0iz���a�a"�����O{&�_ı��� A�42)�^VF��{-P�8���L&,`1���)��Ԛ:ӹ$3>3LZ)r�ː�a;�V���dϿ8ϿЄ���:[���C�� �B��P�rpA�{-�z�h�I����MƢJ�KT�΅��tMSk�7#Qyz��E:������[�����x J�_�׮]�Ѝ7���/}�K���~��w.� *
��g?[�������O��O���Z�qNp����)�{�=�l�fY\QJ?Iq��}�FC2��P�5R�r4-�^�D
�	ŐR�!�Q����	
EhwLM)��
)�}Xja���.�����{�\wM��a�҆�M$!�q�ᚺ�*��Ԓ޴�zf��Z��3��zd�gZV|�{l�\%�f-�-�y$� �Ӄ����>�ǅ�.&�ܥr������D3SC}0=fc�$�B�A)|�N�{&����g����7mkK=#� ��U�	��H!�K��,�	l$�:�H�C8NU�{�"�	�G3(W2FRX*�����B�Ќ�I{#�N2��~&���P2&�|Y&�nD+,z����ecɇ��9��˯���W�p�d
K�Di�>�H�u�!�8����t/P��t����L�&���CH��x��)�~�vz�.��k"��^:�9�[�+�H���r���F#��ٴi��+���?�����I%��7J
��{�]z��z���ӗ_|��>{��$I|�i3�Z/b(���r&�l~Vp���}M�uU�
�ގS�ǡHU���P�N�AX�>�ql<��<Ն��6̜K��\sU	v\^���8��u( Y�P}Y̑��.8Q�5	E�8�h���ԦuM��"Y����.t�)TG)P�Bk�V �N�H[��"2�IE��c�D�KL�N����A�^r�O13@�<S�Qf�sfȒQ�z�����]C�^
���`���ȭ�[R*�����}X��g
&m8�v!��Ew7<B�B�M�K�H�5�����H��ᚾ,�L �� ��%�h�zW+V6l螚z�b��Y���%ܞz ������M8~"�W�v`߁6����CV�М�a�`����coD��4dDZ��@�d&�T�@����"��t�{D��e�aHU��D�1K����M-���+F��4�[$��S[�n��w��?��?Rr�xS�Q�PtA��?��?�����_�T�}
��%���L���w*��"H��t��ɯke�L����#U���N��ѫd���X՜f�ˆ-�Ca'S$�C�����C���	�*�..@�@f�7����̍���K�fuV.�`E����i�V)�|�	NL^y�\Px��s��8`�E&��-�R`�n�"����ePmxH}h5S��ZЮ�|ܤM�&�Z6D�F&p��'m���)h-)2�h,t|k	�v�VQlN���9m�R��3*�L��F��01��$��2�����p�B��.'a��P$���nt,�"�M��6���&�M��/��/1�k���a�Y�D��x������1�q�� )��ЊFaj:�c /�܁C[p�p�k�p9�d�=*(�(���i��Ҙ:��Gҽ�1��Z�� �¾	Q��M)��U�Άȝ<P�vD$����Mq;>�oI�Ҟ/�D6�OMb��M7��G>����/|aBɡ�͆D�Bч?��?�C��@�ѨNOO�Nvkpr�)��Z฽a%E&���&��n��!�b�sw�t"�n��Ny�_��h���I��������0�����gjp�X.�p���ᚫF!Y��H	%�vL��D"�۴7��S�Fn�F)�(��W�JAJA'�V��sf-|�6�	��- ��pE!D�I#�#$��	cͥd��j��$f�����iiHiϔ,�RN��,!$B���m#g�=�'i^M����f�R��26��5��N�(��G$��T��7�PŇ�J	ʕ2K)[�*��R�5��	~n���SOhB����x�p�_��zF�lwH�a~��r�C��7(sC�]��s8q*��^]�W��`r��%Xl.�vz��:KR���i,��Z�G�0���B߳�<���w:	�FD�%O����A�Z��{J9Kt�/�[�~[(�.�T�i���k׮{��o����|���~֎9
��%�
��Pm������٣�>�=z�����ztt4���DW���"��Ӎ2�̤�ګ|Y�Z)j9M�c��FH�V�R�����)6�g�ԡ�07Ն#�f�}�Ka��\�nF�b(�-����N�6*D=���+�kq�Hh۔nC������g�7��/ct#�*#��f����y\�ئ�E��Ƭ�&2!�Z�$��0���|1eep`:�p�ɳ)f߼�������)h1&�^�[shR�+y)*GA*&��_P��|�"��2	K
L�&�"QJ8�L���V�q���m��N�H�ɲ&�;Tbh��ֽQlqX�홶{�g�/����1A͂"���ZH��pr"�}Zp�`mé�1��粔)�`;��0�^$/C��Ǧ�s/�mȩt�܉���m>7u��s(�7e,-���5���<� ���W�KF��{/���<v�u7���o�y/�S�B�@	�B�� �������~���a611�k�z	N\�������Ǆ$�ɶD�8��O������o�l�S��a��>a�jR#st�^Hv���؆�8z|������b�n���K0Z25�~ͤt���.)�C5�	���	Y�60&�fp�ڦx��ǴMN�L`0���d���a���6�0j!� ��JY���z�Z�I���&��D4iL�����R+������#�m��1uu����%�VwdX�LÒ�f�%��d<$�y5�3a���&�r������:w�!e:�1���Y��5���H��kqC�ԤfO�"��az��� ����u8t���|h�������!��'T�-�H�Du���'BG�t�'	f�.��kײF�a�}�u�!���z]��"rH�z)��6�6-�P*ο�liq�Y�V^�l�ևn��=�v��B�A	�B�$���ݻ���?��O��ӧ?��j j��"�Fv�:������C��V;���"���YL��5G=���l4ȧ�n���	��)M�� ������;�/���yۖ.YY�eä8^B�dj���֤���C�{���E [�@S�h<SV'ܥ�/ش-�	��SSc�1ɍM�n؆�s=ID�	��Vs�I$/@k?� Jz�(]*��;���F�R*{&�Ɗ`�UL9mR��N����|�=4$B�#�uͻ]3n
vk�pY%��Zf;�$ƿ�[,&1�^ĶM3k#�"m2��(jUh�8w�	�&p�����p��<LNG����oV��*Cµ�)����\�"3��;&�K�e&�9; �7ŔZL���
��{�{/r�$I�߃,bw#&��  �V�A��qmo�="�k�J�V�Y��o��ʧ~���y��w�B�VA	�B��(v�ڕ<���qB��w����cǎ�*Npˤw�B����-R���t�DX��J�8Y̬�Bt��&�D-�<�o`��W�h�W�	�����A�q��3K059'&��-ر��7�a��q��#(SG�"N�i�←��b��zn4�HqGkU��t�Hf�3�Z��s��y����ZD2l*M�/F�B�]�F�P��K��Ό
9M
�:��w�	��7V?���2��e {���x�A��F�pg�̤�=c�V0�:M�@��"I,qO���%�t�8�nsf>3�d��dX��f�%���*����Lw��W�gp�T��`a��)!�,s�ߞ;��� zF5��m�����Mu��Q��"w;�T�e��%*N��B�P�Qz)���$�,�$j�D݉6�7ܻjժ�7�p�w����T��x��Q�P�&��	I�3??�rii�C�qխ���L����MG_,b8���0���b��"�JM��,��.�g�f;"��L�� #E6�� �m��o�ɉ�?�ÆM �.Ka�z.�T�5+��l�a��j!�h�8�ڝ�itbl_�Y ��SG3
k����Zö0Ah:�p��T�Iҳo��f�$��'�'�~IZY��K��Zp�mZ\ ��]ߤ;��Ǥ�M��:s�O"�ֈ��7M#�5%M��8�p��cQ���%�Q���A�p�2���/�`�6���߀c'�09������EN;{E��;�(uo���%�#Z<�j��&�ƈ�ȣܛ���o"��R&�H`�M-��D���}(������گ���H�wR�nqdd���´�����;5P(�b(AT(�$�����O�����W^y��h4ni6��ݒ>���P�R�E��L�R���b���I� %&J�5���4p����Y<Q*���4��Ȥ��$0��ԇ��놠1ۀ��&:9�����VF�X�u�>�-�H��Ď�EM<rې(�&J�c&���(T=7d�A%�5�f�����	o�vIa�b��YkS�g��1�M�1��"�SH�bE*�魜u_���록�:A���|p��^o���kIM�s���b��H��ӳ���̱�e����+�G]��ڂ��$��Ѯ��Li��sp�t
ǎ7a�|�m�Z-�fR1�vR���Ɛj))�����N:&%O	p"����LҨ�A�DG"�r��##���L�٤�))���QH�Y�
�zDW�%b���2�}̮[�o���m۶=��� 9TŲ�%�
���o��o���}���O<�D�V��ĉ�$=e%�"�����BW�I�$�(RzZ���d�"��+^!�JgW�l&zc&m[i0�	}��KY�k
��YX���FdS����x{3��R8JB��!I9�#)��/t��uE�~Y	�a�ls֭)Bգڱ�	o���w�2����(c#n	�U���1�Eӧ8�.9�9����$�G�+���}iٗ��Zbi^=3 ��f���Ƽo�(B@�D�z>���YJn�gk��؃��#f��)�B!��ڛE"�!�I��жY	Ig���)����M���8y*��'Z0�@;�_�"��ئ'��&qM�~�G��'3Y�D�I���1	O���:Q��B�:AB�2�m�ܮ(t?�Z�>A��J�нo�OѦ��>v���l��t������ի������v�������%�
���@!fΟ?����l��_� ^��tJ4��#�Dh&�Vw�	V�\�`�[Ġ4�=n_:��j�B��E�8f������.!i�'Jǒ1�(��]Q<N�2I�qE��Ӥ�z��(�� /�� �7a�Z�o��%�K�v�
$��j�$�~�OXQ���c�nb�$Id��Dr����\�ǵj F�F�[��9_j<�������ڨ`b��I��M�P��2���)4F��c���n7��y�i���R�HѺ��!I�4��-p���U$�eX���jqm���M�<}΃�� ��4Z�H
@����/��!��q���)� i���i�/3�)�E�I�#�b��a���]?O�7t{��a��&_R!
~���A�U�ӱ,�\_9���o��?��+7�tS
�/J
�OK���w8٥�-��n�ɲHD�&=Qn�d*�U�9�q��D&E�"��k�-�����F9��X������2�}�Zr�����z@�����R&�!���s�D%$Xh���Y��)�>[�e�>���6�_��%X�2���U��P.5!(7X	L�+1gS5���6V.Nr���3�� ���I�R:��A�S�O�/�}i_��^T�ޒ�w1�n��fL:��,}�FN�>8�K">?��!��QIߐv�n6�d2�&��3��:Pk�09���&�b�?����,���Ch�c>��zm�����+6��C���Y�MB�ԈbRύ@�s��@F���&3vϔ?�=)���^�kW}�xrD�����2��r)�~zH�{�#�>�ťb���W^�n��֗�j���m%�
��g�US����������O�:�;�Z�6���1&������MBڙ�d�F	Yq�/�x���w	!o�@wf���������D|N��L����bnHg�g�Q�aCi/��* �	G��H=87ۂ��P.�`ll֭��MCp�%ش���KH"Ga����D5rm�[&Q*���+����&ukR�&����M�\f���a��!u���������Ey�o��q�ӳ&Z�ٖ|�KR���C��4B#�!�B���͒�Nǭ ����>[���	�;<SLM�/ ԛeH�a<~�/�B�~��~�p���+$p��U��i��ѳcBs��|ڌFr�؄�C"n��� JjXH�Q�[��,몠E�Ͽ�}�H���s�q����W�Ӷ��������*FQ���Q�P�\���{�|��o���?���~��F���7���G"M�DE�"v&�W�څ����5�n����Sz�]6��۬�}���R�o��ϮgS�ԍ��A�&-IV4����4۴H�����$q,C��HvbX�Ep�h�*MX�� �V��a��_[���a�J�ё�ô_jbҚ��t��k���{`��R�gɎ����b�xG��|��OU֖�7d�%���g��_bӸl(��P*�ZFj��scd���%�7BX���05Մ��1�>Հ3g� ��^�.��>i�{dsQL�6mVvSt7ߪ���A�I�tr'6��&��Aׯ'�.?�Kz�s�4��5iz,��N�'��
HIj�G�P��EH�*������u������b��
i�G��I���Ζʥ�w\y���׾�_mlo7(AT(?7��n
�<���~��?���3g�|��J�`}��I$BH�ISlC�QRq���]���r6ۛ��V�a�OD�3�!�/PRʜ"#T ?�ix��[�cd�E��55xG�(SPZ��	3ꀒB����`a��g8^����Xт5�0�"��cX1�g!T*�d��b��IJqIP��F��q�/0*�%b���/����.�( e5�9�Բ]�9��Z���X�c�uR�	r�V'Er�A�0���/�+ 1l�ܼ� �����X��vs�X �v���.��q~h�ڤBiU�ǤT,��F=mR�A!d�#N�w�e��muRS���ߏ��%|@	�P����Ct�
{!~"B�{�U5����A�L��E��P⿏�?1>>��W_}�_mݺ���C��J
���m>  $%IDAT2x��������O?�t�ȑ#�'��8���Z�z.�R�U<�9��un��ঠ	&�g�Y�_���ˤV���Q��1M��h���c�cɳD"��Z�Q$�k&h��F5>D��4����ӌ#�/���t	`��8�j`t4�5+K�f�(�//���FG2X9^�ec#Q��;P.DH^"<v"L��P􋍬��3!v��
[�[��{�����k�2BϚr��H�N�&��$9�݉�I�Ȑ�Z#����R&��f|��J��BS�\�A�ILolVV�C��R�c g�,	YdDc�p�����(1��8��������95Jq���=b/�{d����a��rW�BQRI%)��#G�%�Y�6�\�Ha�� 0��k��7���z��m���\r��;w~c�ƍԱ��!� *�7�g6y�����o}�[ͽ{�~'��J�L����Q��滫�}i	n*O�rh����g!H7->�&���q������ S�Fb��τ#f\��(f��y��q��}f[�ڒ�`a(4��(��^�ܚ��e��H,�	,ԑ4��!�w�	��Q$��F�|�e`�� V#�	��
����	HH�ˌ��E���A)4͞�DL��1�e�����?"�D�(�f[�Ԓ.� J�v|h!a��c�_���l�j�[�`f�ss �&I�jp{ꝼ:�"'�9G�lƜ��*�Y��^L�cl�_���E��r�� ��� �w;�Q�����Ȧ}�k7f��R$�T��u�mm���#��6�����44�n@f]O�,�O�W���"�0D�ѽoͰә���j���֭[��;��?��?��(��5� *�7��s�i�$��{�<r��}��]��7�� �:l�	� ވT�%4����禞}�n�\���Y"��9�l�XlO����ۏ7��:DIM���_��I�6��w&D� ���p����Oh_$��2Rb��K
�9�G�Er<�:D�1��P�"�	�)�q<<��R$� � �U��h���P,��6�Ԭ�����X�n&�V�ҤH�n#$�jWG$/�Z=c��V��q})�F3�u���C�H���PE%
�P�h�5!GuM�>3l�:���S� z�j��>���Lk��{I���2�,1C?3>� Yq����J\V &�R&�H$�S"�p"�z6
�K��ݳ�UJ�G8N�F��P������(����h����3���k���+��+��8���ɟ�	(og(AT(o��t�R�ە�?~�������\�q]��t��\w#��	�Dr\�)��nh���>dV��>�3ɻ�>����z�z�h�Ӯ��?�EM�[+jic��;?�I������Kl'�ڽN�
���x虜�����K
�" a|�� �P*#)f0\F����
ŀM��fѴ��L�ܘ'�kU��ln�LŜ�Z���I �A$~D5"RH�"\P�1�s��ϩT6�~�u���v&ޖ������v=i<���@�e�U	��>��Ϭ���aɪ��G0��Ț�|���tr�?rл����eH=��n�c��#}�����/>eHc$�+W�����^�������O�
�; J
�
�6���M=on�+�LMNN'��8q�(�BK�р�j�;)�D+�C7�h�ۭO��W:����u�ٮ��\B�b��va��z0Z/A��v�=kW&�>Јi<��.��(�8ŝZK�N5fڞ'qЌ=6Φ%��`�1Dզ��ER�"��9
g�{&����+���^�v�r7`� ��q��1F�V��}�����B�.6�D�܎:��|_oi�(�^E=/�i��	!���xB,�Zn���	{~�]�l�7E�)Ռ4�so��Ccccߺ�����?��w�uW�w� *�74>���?��#�?��'N�<�񥥥�p��	��H�k���'Ůp�0��x#���$�y�}�������u�Id��i:�\Gx�%2iK�w��:U��(�#152��Ȉ&�"�Ԅ�lB6����ni&؎3,���!�s7�]�
�,tXTfI�3�!� ,���H8O��$k���I�^do�o,cN�P��n�;����5=����-��m�'��QF�q�K�D�"<�Z2��?[�V�{6o����o��?��O�q���H�x�C	�B�x�@-�pB?�_��/��?=��������jށ�֑ʹ^7�6�؅\�$�Z���6A&�|iP�'O�^+Z���bQ�����Ai�[~_�B��Bv��L�$����Y�B��l|M$0ɐ@�"O^�]GjkVg�5��"ft�}�5��1$�L�~t�2H���p�>2����-��/���+�<A/�l��X,w�a��k\��C&!����ߗ��{��mܫ}���1P&�~���"6My�d�ll�/[���/������~�s��S1��%�
��M�ǒa8�����M�{�{���ɩO��W!Y�t:ύ�H*�&^IG����u��aq��=�@�(�غ|q�z����b����G:	Ɲ%鋐y�\��g&m�N!�<�@7:m�����D�{���sf�V��v���8�xݘ^֬�"��;�l*��d7G��|� :O�]E�����_������F�Wz�0c�v��J��.�uG�����*��v�{��&=����._�����v�W����?���7q��%�
��-���ݻ_���'����/NM������;���V�Z-�&{�=�؄H�A��.�s	��j��\����"��Ϡ���������HY�%(�CX2�s4/��OL��D��'��׈Pz���$�����0Rz��d��~Ҭ��6z�b��^��Gb�c"�)���5�]2k�ӫ������@��	[rc%�@�}Dέ3t�v�Ä�BIs��{��h��c��y�;��ߡ�*�9\�re?;�/�Ab������9H�sP(��P��P(�2x�����_z�����L4�~���������6�`Kn�ȵ���Y�����T]�����XD������.�������~���I�)�G|V����-t�S�<cc�Wj�^f[���H�^+&�Lۦ�Jِ#{�.�e���\ck�����(����%ukA���8��K�4�%u�Z�QݟD"�^�U �=��:CW%�O!�������Nvkڎjj������x����Ν;��/|ᬍ�+�h(AT(o9��ݻڻw�~uy�����_��C��_�gg	Y�&6���ˑ�.4W�*0T*�-u�d��	5r۝�"7e��m]�Zu�$&���;Y��hؿMl�?ߦs=0Jh�&�^V�5���1\ /����=�C9w�5����[�u}�0�X�y��~&��|_�ѐ�ش�K��"7����m�zc��Qn-�lK67��R�(�΍.��c����=�|]�A!��F��Sl�E������u���#�~�#y~׮]�{��w� *�_v�h�4�y�g����KwMM�ٵ�T�'�a�lHtG"<3����|���|�>��%2n$k��=n>�z���[�0�z���=�����Y�u�\f�v2ٷg<ɣ�wZ�I7g�-d�M�o�' ����O��	��[�V>s�ܱ��%p>u,D��8�}m�\!ˠԴ{��Y��F5�����ݯ�7��i;*{�������!9��7��m۶��YSʊw� *�_(,Q<������W_}�={���c'>Z��/+�J!N�)D��K�<�$�OK^�.�]�ֵ��O7��n{qAK���nc޻�uqi�|�'�`$��.�m�hI��ua=m��w{M�G��4*]S�螃M7���lf�"�و�Hf���#���u'}$� �Jd*���,*bW�쎽D� �k��:/<qS�n]�����SH*AZ@�(��U�S�t:m�ߩ5k��`ӦMs�m����(�P��Q�P�-p��wG��wߞ��ꯞxꩧ~��K/���g&o�Iz.N䞤���a�gaB�G��\L����$.����b���$�"5�R�L��xZb�Y��g1��s�
T�Km��?!��&�����ufZ��'Ղ+#�����e��4��6!`�ߠ�K��H�����.ATвo���Ä��}O�Th���6��`��s��n��v��֭{���/����_��U�V��7
ŻJ
��H�a��޽��qҞ����_k�k�E�e�Fc'�"�6��J\��������!�h�}�VN��t剝+:�^�#���g����{�m�g�[�,���c�gB�^ϵz��c8�Iۗ9��	m��{ &�V1A�=��tR�'J�;�B�{P��C�֏@B��f�&B�����e/��3Hϓ~W���������}A��4N �4y�X�P�+}��mGQ�f��]��;w~�����u��w�qG�w9� *������G�Ꮾ����z���=sn既(ڂ�.>N�۽$/.��!�T��Z�d��O��S�����A��}`;�X�Ag�A��#�zņ�rF��˦Jz��~�o/5����K�s��zV7��T{�6�������T�K��?�H;������k~��p�&�5�yCٗ��E���Dj ��|�R�47\~n��M��Нw��=��3�BY��D�B�mMF"�G:���}o�8}��333\\X�\��*a��	1R *f�h;o�#�f.Q̧D/F����\�f1��Zw)�#�^���K$L���]f=����`&B��S~��	�c��c;��B�Z�>����~R�����^�S)���]k�<)tE&�{�	O��eP�ߌ঑��:y�H
dp�H�|��]��j���Q/�J6o���l��o�������Z���{A�x�@	�B�x[c׮]|�|�ᇿ����?��SO=�w����ggoiG�U8ї�o�%n]���0q��$�M7�I
!o����Cهl+b���%]�f��'bɬ�$c���[�X󛞄��ng^�s��7 ��w\s"�>��K�2WC�?I�)c����/��W!������U�R7��P��rrݡ� ���/�K���?�qӥ�}��?�����,�C�*�sP��P(��N,�2�}�UO<��/��!���5N��"�	�(-ֈ�q��@��t�	���Y�Au�.��㹶:��g>
���d��I�͜O`}��z����u��%,��r��+��pq���4�3ݞ5�6m�(W--�R�W��#�B؂B��E>��+���{�ﲐ�v>�}f��#������T����r���r�d�166vlŊ��^��髮��;w��B�D�B�§?��:�<����������8䔫�?�D�}H V����R�P:�Hj�UӒ�U��[��
^�)g���#[�-A���I�n�������3����|�bQ�Aiq7�w�����kS�~cq�t���#}��<_����j\���1H`B�@��,K�:�^�c�w�6q�q�^y������+��b��nS��{J
�;��ԧ�v���C�����'?y|����455u�+����N�S&�122�aii���H��Gp�\��<!t��
\�=7R'�Բm�Í��ۺ۸��VZ����:��-��%̓�#�[�a��ݱs��%�A���uSƴRK�e!��Y���KX���\��6.S�J噫���w���Ԗ-[�~��]��ò
�{J
�;և�,��]v��cǎ=v�ԩ���|�'�K�<���J3�)`�&�
��h�tu�4����#Y�>��{7Җ�����9���m�'z���o����H��%���Q�K�KT��a^�Lp���H]���Mg��q���Q�T�Z�|�sk׮��M7��#$�G>��O1�:C�D�B�%�3H���}�g~��/܄����z��Z��		�(D_���CU
�^"��e~�g/�][���I��s۶�� �ˠ(���X��b�AQ�|�3��|�݆��� �*��=gw��p�5�>�i^d�F8=����>�A�C!�ǐ�;~�S�k��d3AR��j4�Nq��K�^���[�����k�9����ٵB1J
Ż��M���b�w��H?t���{�~�݆�q;�����հ�{��\��M̕�}E�F�G.��+p*�1\�@w�|͜l���̟��ύC9t<��5���w%RGp&���~��^*;�}�ݷ�-c!u����ύL�X���ĸnztt�Ȗ-�}��x�wo��C�b���P�xm(AT(�:�ta����{l������C�x���¯!q��^�_���p7�5 ��%:�i��tb�!@y�m7F�7������n~]>Z�zu����b)��߃�C0HA�'}.��ZEw�]����D�����L��D�Baڞ����;S#��/�Y�v��m[^ڶm��K.�D��B�SB	�B�x��
��pI��C=t�{����-�����/�Gѕ�(Z��c�h	�,�via�lw��!,-�ӫy�yAJ��O\宻}^��OU˶����k~{��m_�;�zWP��
��N'���P�]c�<i����'�NG��Y�Y�T�'����lt���v��s뭷���'?�z*>Q(~&(AT(�	X�@e��|�W�{n�ĩ�kOOM~�V[�:Nӭ�n-.$>�Z�z�8���9D�!B�d����!1DlD%�'m��E��u[�j^wB���s�'������%��"�y2Kb�W|���F]u��A���"��az/^�4=t�+�5<<��~���3��š��7<�q˥��ꫯ���/~qAI�B��C	�B�xO�����$���/���r�����;u��ϝ?=EGFFV���N�5H��K�o_uh��#�F��#�Cp���D"M��ŭ5$�D��F�!Y.��s��� ��扜[#x���������ʵҸH
Z�(���D��S��č$V*����?#ߢ3�##G׮]��m;����{ｋD��>P(??� *��4l��A���W_}��'N��055u5���Fc�?s��f��	�0n�������J���I��"��'Z�=� ��+I���=���=��%nyCٯ[3��Iʵ�ᴜ�����#���L����n��'�W�<�E��
I%I-�p���Z�#�Z��A�~ptt������7lذ��+�8������o��7���@�P��C	�B�PX A���.�h����]9r��Ȟ={޷�T�����V$;k
��e�bq�*��".��A��l6���y�'�%l�T���?�Kʤˈ��uͨ_O�"� ��!u"��(i��Q��Sܢjv[��vt��UC�j�a����&�3ccc���G���O�^�zߦM���t�Ms�v�Ҏ'
ś%�
�Bq|�c��".�?���Ν޿��\w�����umَ$g�*�5�j��ȣ�:!�B��I��Ϲ�F�l#*^ImKg1���UM�xJ��5�����ēa>mM��h ��]rL�F�C6C�7}�y����$�!�=��'׬^up㥗��+~�cǎ�j��@R��B�C	�B�P��뮻�߆��>��$e�|��፯��ʵ'N��t��n-��H�(=��CH��D�\宛J%"%ii����U�`�u~����� e��0�my�7��(�{��w5�7*(ۋ7af�*��M�G���i��J����������'֬\sb|���KW^:�����v�
�[%�
�B�3�
\�#љ��W����g�k4��fqqq����J\�!z�MH�F�0�w���RҁD٤m����4
��\�๤N��R��GJ3�!�㦑�̼��.���b�H��Z�������5k�Y�l��B�_�����36l8�v��ő����*�X(AT(��V���e��E|衇¥��ґ#G*'N�؂Dq���"E7�6���$Uː���<��RZ�U_L�����Ib~�����m.A$���%�RGH�	q�Z!K���p�����K��I����׿�$�Ȗ-[�oݺ�����[��=�=�B���%�
�B��3\:v���y�=���E$[C���+N�<�	��V���ӹ4���q� ;�~ѸPzz��!E7:�&"Ȃ�9�OL}�χ(���[Hg6�g���F��pGN��5��ES(�ڏx:�
E(�z�>�'rH=�q?m��Z���v���q5\FFF��c�7o�@Rx䦛n:�nݺ�����?� *
śK�v�	�C=t�������e1�.6�Z�6R������fc��qW���Z�����$��8I�0|�h�j��R����n��Są�9�瞫��y'�����<IN�Ec�r�4�M:�M�S:��ʕ+_޸q�5k��-[����i!Ql�9�p}?o��o�f[���w� *
�[K�$¸��)�c�=���l6��W_���#SSS+��ٹ�J���Q�!��K�b'��H6WtZ��H�J�j��x��� �l�(����$IW�Z͑r�L�`��Q���$B�94�*��- �P��I�H�4M(!���](��xn���-���r���^O��ziԮ��c+�W�X1�aÆ�;v�hn޼9���ۉgy2���|
�;J
��e���)�H���C=�Z��[�z���	I�w��9��j���z��b����~�D0C"�7���ѣ�<�ba���#��իk˖-k#��qߴm466֡!n�C�8�-sJ�����"
��xtt4��Hh[<nv饗2�;{�lz12�P(��P��P(o3X��sæ���{�z�Ї���O���/�*�Y�;ޠ�
�{J
��]K��T��כX��B�p�Q�P(
�B�%�
�B�P(�>(AT(
�B�P�A	�B�P(
��J
�B�P(}P��P(
�B��D�B�P(
E� *
�B�P(��Q�P(
�B�%�
�B�P(�>(AT(
�B�P�A	�B�P(
��J
�B�P(}P��P(
�B��D�B�P(
E� *
�B�P(��Q�P(
�B�%�
�B�P(�>(AT(
�B�P�A	�B�P(
��J
�B�P(}P��P(
�B��D�B�P(
E� *
�B�P(��Q�P(
�B�%�
�B�P(�>(AT(
�B�P���	�N�d�s    IEND�B`�PK
     ˡ�Z�C��R  R  /   images/b905cced-8669-4310-a345-cc026e3fb08c.png�PNG

   IHDR   d   ;   �:/v   	pHYs  �  ��+  IDATx��|wxUU��{ʽ����CB	�t�2����J�Qfut,��gEGǮ����"D�4TDJ���@�����'��=�{�?�0�[���{�=�{�{��]k�}e��:T���~���� �`�7@:X����7�ļy�зo_���a׮]�}�4�r� �"���PTT�7�xӦM�ԩS1p�@t�v�r��a��/pʠ�x~���a|���hii�/� �\�2
���o(fRRRt֬Y	��Ν;����֭�SO=��K�rp&M����		�'�|��>��w�1#GGVV:6mތ�'��(JI�NINN���Ot!���PSUզ�,�-uN��]�9++k�s�=KKK�;＃��\s�5x��~���P�̞=�~�K.�'�ꉴ�����ݻ'��dOlhl�隟]�v�[Ô�C{͚ 9��iY֙��!����ͻ���gм+Vl�ֵ_o\��������O<������'�_�y9ٝ���	��tu�ڵk���/�,��� ��$sDQ�e� �``�����[�l�)ض��0�;���n���/#�yy�/�*큃�p�����o���'���<! 5�l<���ڣ�,+z��^���t]��z=���5ft��m�  �M�{#v�%� ��vb'G757����]B�>>g��ug�g�:��̽�������r�X��Kt�R�䀿Knv��-�c$� ��M
���@�#��"���O��3,HtN,pHL�>C����s,�Se�n�ini]Z��U_�pЀ~x��W�{�_.�uh@F�}N;mr;g!-=��U5喙��rK�'p�͌l����6��U���@�b ;C��G�'�thɨ��P�_ƮJ�j���B� I���$Y�O�Q83�#���fw�+(��P���^~]t,X�����rޘ1����p��w#�S�أ���|��#���ɘ���k������S�y�� #�&7����� �R344����k�X���MnȮְG�3�a^C��|۶m�]�
'�X�x�g:�|��v�w�d��+���>������767�c��jM�8Q������8���0�l��5ǂ�pH@�IA�I�a����\����L�T���C�8�*�����>|�ʏH�IrB!��0�a;w�Z���9����|��O��Es��v�{�����#�<���\P27��94S���%�Q+0eD����n�RE�<B��\%�刄H�-A!��0e�$�d	d`��S �'�udv1��UC�BN�1|����Ƕ�^�-��x�(� =VG޼��񣖕-O����ڽ��ٳg"//i�����ώ'Դ�?�z��AD-j�i�����uDjE4ՈP#D��ހ	oІ��r��O}՚����b�+ɩ�1�E��r	���ЩPG~Og����~Ͻ�c� $��h4(�-j"~Ƈ�{~��74�I.�rE���Cr��I��=�%e�Q��7���+�s���M(��;~�ᒑq.�?("�h����F�r5��YILO�7=oXS���v�<\�M��t	�Op��V��KL�.�=�AC���	dx��^s˒x�����1�M�U�}�ц��WUa��E>�}BW���;df��ѽk������z���'t&S�n��b�	� \CU�I��+�����U���i�!o������,=���v-�[�(Dc�܅�>/�v�!�
ݡ�����(nN ���?_C\�`�nR^����	M{� ?��P8�>��v�C��ګ'�wi/�,-�/++{��b_�:~^�L��ܡqa�#��H�N(�M���)��w���`�$�>CѸU�w}�`�8d����O'�y0dر�&[k�����C�����N\R�y_a_7O��@��-;=��� 8�Dc��U5��L�����ʖ�s�<Ӗ�a yHOOAuM�5�D�d���܂�j �,���+��SR���<��Ռ	�]-_F�g�����4$�|�x5܃nQ���1"�=��G�BP��e����o�?AIa���V��|�c�/����| ЩTō�񴌰�T�^��s�ܹ�&ϙ7~��v��/Hk�߶o�=��eH�T
5�a;�YU��d]�~�N@�{���aQ�&2�P�PȈ&�NH��v'/�9�ȥw��"e�8�g�B7B�2�ru6Ē՞�W �9I�z�&񂕛�>�?�>	qi4o��өh�a�C��b[�EڱQ�7��ɤ�Ɵ��;$@���B"�
I�J��0.l�D�� ٷo��z+�u�郖��23ѧ�ɪ�R�H-�����l��B��ؿ⒠������oSO2��%E
�jA���I���U��mC�f�&��.�DaKB�xw��:��*�UKz<x��'B�f�d���.��X��W
��"S��)���=�q�Ẇ��p�s��9���5�'��h�ߨƞ����^T7��3�asN�F��>c�޽16�r�u׵Ɏ��#�݃!�G�����������|D�ţ
�@G`%%6�E�v�-�]ý�\q��O�*`@w��E~~2~�t'r��Oah�g58��~�\��%6lK"�q�bk=��Fznx	��?�>�k)x`��1�������&]�8�_��w�۟y[�q���=J~]79Ŕ������\pyD��� K{�ڵ�/yˆ�Ɔ6۱� ��Ϳ�5�OE�����5}�H؝ ���������ɽI��	$'���h��C<6pɸ����CJQ��>�y�k"��(L��M�[l�!}�v
���h�P,����� ٭�	�ڦ'��b�P�Q�g�(eCNu�~צ��O��J%%����6�ħ+M�4�_Qt���0�ӧ��f;����Z��y���+(8�O��EL93�}�6��rr�s�x��� II##ÄG����V:�#v�$$��zQ6�CVN	
"+��es�:æ��(vk	����8��Pɳ|�r r�r����c�{��%�����odT�N�k����K?���@�#;zTFAg�
l|W.R�hs�c�<����������v���f@v��s߅�΀7ʏ*JQV���:a��g��Y���_^�j��ɘ.�n����s$Ie�q���=-V��gD�?��y�q6������k-v����Su�[ʗ,k���z�/�m�J�NQK�D;VZ(9 !�<�W��ow��sI���(@��������[m�=���B����G05u���t�<�;tD�~܍]j
tC��X=������(�nRPl�o{�QM�d��Q�{�e��Xh:z,�)�����̢�H���q�Ƽ��-LJ�t�y9��H)��h�����=M!���[BJ��h=�����"�h6�lEӵ�f���< �з���p�U�MZ����^NCDɄ/�@j���u���lfLF�lzՠ��(u��yDcH�f��题N�Tp&��/���4?���7�M2u�<Iw.��0<g#��C�{���V�<�����K e������m��*o�{��)"Ro�/d�`9�n9j���H$��!I���Vs��x8�7ʾ>��fJ0)Ȋ�X��A����n��@"��bܸ�@y������L����zO�3$~ߟ������?�8��`�ypqfM���`zz�S	�:��^�ck �_�Q������2](����h���dX	���8,��)�%� 2'R�U�Q�-������YVd
mnmd�_`�GrNT��H��nj�� )�%�pf��Q��3X�,6�JƓɆ2��sS^�P83-�u�;a�I�d�Y�����O��N�K�5s��R
�[B"R�@ZW��'������"��%���14jF��ax���-����-�z��&�Y�S��3/���iRG,��4-mmmD'C%,1��-�h4���}-"rRTNqܘ2�O��T�cv�Xm�C>_:���c��/�Z?~�W��yA'p���}�s��wy�"[�rp�� ��T_��M)@Y�B���&������~CL�ĲN0β�n4u���΢4�,8}k��w"O-�L�D[[��3xʞ����h5����#GP��E<a��=�� ���0�$!
����|,����E�D��νm��Z���3A�$��@�[Ø�),�9�H(���Bm��- 8@�������7��kV�cY��	Ŕx^����x!~�]��Ѽ̙\��� p��}��W���n�Ų���N�d��ނ�����پ}��|9��A���EjR��ԕ�ܴ�T����C4�8Y�fI�Mj�nIk����g$~�;���g\cs �/��P�*Y��΋<���D�
�A"R
��݈V̏54AR��P�<��C���)���)� �#D�1��R���C#�E���x�*�P������c�bDG�lI۵�G��P��G����@QEd$OЈp��������a��H��1�E_O`�y�W���l�x�Dh-�p��S�q�y6��%x��_*���H�	�`.^��Eܽ8�8A^\�ww�ɾt&L���$NT�<�y*�-C'�1�R��꘠hkk3 �� 8�4%�]��CF�ᐎ�ڀ={v����Y9HFvT���`ʅD�a�#�Z�e�)F��SbM1��F3�Gv4T�F��x-��r>ȏI�����T�c���W'���z��R��m2�]km�M7y����|�=:��eI�=0���Lx�PdV�e<w~����S��=֮]�&{��K/Ï�N��-�����U7EB*rD�&O9R�e/#v�n��1�GYp�������̠�Q_�%P(?	��M��gD_��:���s����)8��SIŹ���<�`��ú������j7�	���CJ���ͺ��1��!�1������B��E�LYV��}R[��~�Ŧ�f�7b$�����ͦMG��ؐ������mYF@�$�dX�K�p��3�h�v��r��2�(������.(D.�N��8��	L�@�D�)��l[t� �"�X���cN�p�'�L"	<�p��%�&�۾o�#��	wA��C�f�UR��Y���(	d� 'Yض^Be��B��[� !����:ee��|G���n�L7��x&�TTĎ9��֭[����s��$�[���B<�K�ͅ�,�%�WY�`:��T���5#�P3�7d��e`�R��HS��Sp{)��V#�<#�He��(_��l��%z�J0�}�8���j4���H��$Hn>B�`�[ע�aV}��C;f�[����t�v�=I�<��Q��UnF�\�)��܊�G:u������C��zv�܉9s��LcǞ�Ԍ�H�{��o[�D��I��J> ;���X���%Sd�r~A�>s�'9�/Z��n����E[�!.;C�3�M
'MؿMB�Q�Lޞ�e������n�F��Y'����h���Я��5H/j+�eS��)��������f��I��<�m��|t�;x*�us��T���'e��M������V���[A}=�bY\�~����^{-n�����u
�gϞ��5Ѧ/Q��k��g-EЛ����=;+�f�W�U�C����6�����$������,�z�����,���K�no�x���^xZ���1$�t!�^B��g�u��p�-x�&��^䧾3ĜI�]���U��Z�a)j|��}ܣ�_�	eu/�]�^'�"Ҋ܈h.�=�Bܙud����`�2���,.�B�qW���W_��O�o�����Ds����ܗ�V'��7ܸy�e�|��K���u�1D���]��ƺw?UC��	haRJ�;���w�����Z�у��/CΈ���)���*�zٿ&�ɺ�m�͌��H�6x��J�����L�����X�2��.[�5ϏU��U�%��HPN�>����6L��Z< �V�n�}:̪��g�����7`_FF��]��B��� -aO����G�(���G�6�	��I�+��
�+��������!��H?�~����"++� ��wgi��i�Q�B$�@fW�5�q���j��S�&�O��M�x�=�;2�˒�֝Wj^^�S,<��]���~�]��a 0p ƌ���|�����_���Ds���S�v��-�����]6Jώ �T@�>����EE���{�ٞ|�$\��!���S���f'|�ŨVe�%��O��GO�0���b�v!#���^�u$g�X�]|h�H|M�U)��آ>��3���|�K/����׬m;t@X�6�&\{�5h��oq�ܷh����QD�HI	䚯e���O�i�$W�k��*�Xm�HT�/ͺ*e�.�fJ����W�wp��ӝ���B�0�-���g�-�%17�^���i�AIIܥ���s2�6��r;�+&�)(�Ǐ�۽��=.Y���lС 7n.��bdP�����rr�1�1C��ϻC���7�x_����q�-����RB,d�0����c�G�r��ӧS�c�V!���Ǉ�����{H����0�rJ5$�舨.�$�x�D�2�>��|?�?1��eff�q޼y*��^{���/������G7|������W���T�䆗�&�t��iq�87��8��nf�t46Q�FS�������Zt���p�C�ō-%�L1��k"��@����ow����
�ֺyn�V8�'��*������	�hl����p뭷⬳�j��w8@X����p�}����c�ܰ�OSht^z�L��+��		o��b�ƏQq��h�*R��6_6�jܙWɻ<>2t�o����Iʊ|��'K|�RBc��9��͋�I	������ظ���a@������	�%�]�'�|���:>���I�1���%A�fRjj*/Tjl����S��x�-fͷ0�$C�'Ы���L6�m\�g�e��JB ,� ���w(X�Y��r�a�o�y%>��f����[J] �2jY�����9#FRδ��{�����C(l�h�:thr��;Iz>D*G�Y�U4��Z�8l�Nc��ūz���HKR���~Vzr+��"]GB��D,�*H|JV�Vog5[�� 5�2�-IIIS�؎�Ç1r�\��r��_���(7�t�,+À���o��'�
���ZZ���{˖�8��2�~%IN�1���u"j��)bk���3���i�ݹ"�ٲ&O��j��R��_�������Ё�1t�Plذ�W�ߎ���:4 ����+�Ga�}����t<���_�v�-�ߚ��X<>=��f����f�|������A�غ���� ����|�z��� ��)fqUJr�c���u����e�	&��?�����am����XXTHd���ys�D<1�G��v��}�(�,�<#�&��^;�~��O�;�H[�9�W�y�`/����%\�����R^Q�y�Ҟ���_��p�������U�zB r�����x�Ea�[����5���ꪏ����a�$�!C���#%��`���J�l���� N`�%t]?�Q<߉��UJJʊ�[��*,(����r 322���UXI�_��P�k,����R����%�ki��4mnL�Υ���ƍ��aY��J���*/�U%��5�n��>}�Z�lY�SV��>�OFCc#2�ұx�b<���z�NH@������s^؏��v�l۶M�TI<^��Aנj2�V�kz��՘|�D���[�v�4\x�8o�y�5{��O'4 ?o,ga�m�y�;w.�ʰ1r�O��c�lق��u����k�O��@������9����h��v�    IEND�B`�PK
     ˡ�Z`$[ [ /   images/dd9bac2c-35cc-4be2-808f-eb026b88f611.png�PNG

   IHDR  �  �   q�y   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���y��u}�����;g2�"aO !�		3眙(�l���R�RAp�
�֭u�]������Z��V�K�ZŝE\+J�K����@2����uiUf��3�|>�p��#�I2���|�3��U           dV�           �w           ���;           ]��          ��`�          @W0p          �+�          ��          �
�           tw           ���;           ]��          ��`�          @W0p          �+�          ��          �
�           tw           ���;           ]��          ��`�          @W0p          �+�          ��          �
�           tw           ���;           ]��          ��`�          @W0p          �+�          ��          �
�           tw           ���;           ]��;  ���p���*wƯ�R������gkDl끗�����
t�NDl遗�ZD�I�+ ~�#���й�IJ@w��G{����"�rG �� @71p �%.����� U��9��3 ~�{G���h��v~�ގf��/���r_��G��?U��ϟA��򦭵�F���}��m�0w�Ϲ��⏶u��AO�u�Z;w�/��Z<�;�7�)���~� 0t���          0+�          ��          �
�           tw           ���;           ]��          ��`�          @W0p          �+�          ��          �
�           tw           ���;           ]��          ��`�          @W0p          �+�          ��          �
�           tw           ���;           ]��          ��`�          @W0p          �+�          ��          �
�           tw           ���;           ]��          ��P� � �<o�w��G�v|��sDJ?����Fl���E����m��<         03�͉T�G�eD����E��~�1�NĖ���綄�C��9z��;��ܝ"�W��{F����[i���v������%�����n���`t�IăD<�@T>����{��GwE�GwE�woD{t�>?         �)k�����´����o��x��1o��c���tvl���@T��������g��pǶ�?�0��3�e�}E�oi����ϢH{����S٧Z__�n��m���N;����~a�����w�����OV         ���/���Q�@�����k��=�����;��*�H�.��uADD�_����������]Q�sWT?�~T������?�货�21pg�H�z��#tH;�h�������������t������G��M����)�o}#��~��         �^�k�H��bɲ����n���y�D��K����m���߉�{wn��q{ĦoE�m[�N�d����v��ly�!���1�X�_i�`�+���G�ۣ��עs�7"6���        ��T����}Ox�A�;"��=rWM�z}��x�A?;L�ӎ�;��s�ף��ע��W�z�'9+a���}}�;"�U�(������Ey�_��p����[�lݺ����[��/F���]         S&-^ő�H+Q,?,��/wR>E逃�<ࠈ�Έ���ߏ�Wn�궛��/Glݚ9w�Z�s�(VFZqd��ss'u���(V���(���޿|Ktn�|T_�RTm�]         �7�?��C���y��=�}��}G������[���������ꗢ����y�+��u��%Q�>&���F�gQ��5Ak�G�v}��ht�rkt>���������]         �Q�y^���(WiŪ���u\��"�82�GF;Nw��'���OE���殃_૜��^Q6VGq��#-=0w��S�E1؊b�նmQ}���|�����و-�        ���Ŋ#�X�>��H�z=wь��]�Y�Gy��Q}������'����s���;�</�c��'D�dY�Y#�����ض-:7.��pT_�-��ɝ        �lTQ��b�I��mF��&-�?��D������h�#Q}��Q=�9w���;�.pP�O�r����9�sf�z=���D��������?�yT��(w         �@Z�[Ǭ�b�)���;wά��,���/���gEu����F���"�*w���;�c�.Qwb�N��Ϣ�5�wv[��gGyꓣs���F�˷8�        ��UQ�jD���HG6#�2w�$��F�F1�6��Gt>��h��G"���40pgJ�=����3�<�Ĉ9��sx,�2���(�����������El}4w         =,��V�igGZ����Ϣ(/xV.����?�3��G�,f0w�D:�(O>3�5�GE��)�o�^ř�F���%:�Ǩ�/w         =$��5��N���3#-�-w���Hk�G�����vS��醨n�z�,f w&OJQ�Dq�9Qth�&Q��k����I�G�����>�{�Ν        @7�c�(�8'�c�Q��a�E��QGu�ף�O7D��/�b1pgR�GF��ߊ�ly��Rߜ(�pj�N����Kt��Ψ�'w         �d��Q�vv�O�d�>��������ۣ���-�ϝ�`�΄�C���H��ȝ�t*kQ�?%�cO��'�%:�����/w         ���F�ĳ�<�L'��2����v�+��oD���::_�R�$z��;�R,?,��~˰}�����.�yt�wCTm�]        �4J;ϋ��Q�pZDߜ�9dT,?,���::_�-��������I� w�$�{��>=���E��;�n1�?��ώr���~��D�#��sW        0��"���E��gF�uA��H1�*����/|:��Q�sw�$z��;�Mߜ(O:=�'��n������(����Eu�͹�         ����(�vq��ȝB�J)���Q�����E���#[rW�������(/�4�{�N�G�}G��WF��/D���-��~�;	        �I���7�s�����)�9Q�~v�G���w�Utn�XDU客���+������Ϗ��S�Q��p+��޿�����͝        �x�jQ�~Ng��^�]C/�ma�.�"���b�/�(���_�"���;�UQFy�iQn�(bN�z]�冋�8��}�[�����E         �AZz`�.�<��s�0��QݟF�=�7�xOD��;�.c��/H���"�ly�f���Ҩ_����ć���"�G��N        ����Y�Gy�YE������/���Q�E�o���o�.����^��)O���'Ge�f���r�)Q1�oKt�v[�"         �i�`Ԟ��H{�;�,-Y�k� ��w���7������DZ�_ԞsU�u�f�����WG�#����eT۶�.         ~��\��3M�Z�g�Ecu�����ޝ����+�l�R��O������L���<錨�����? w        ���������g�3���%Q���Q�|fDJ�s�ȫ�,�v]�+^峞�7'w�XZ��_�&$        �\~z`��o��dY�f�z=�/����EZ�[�21p�������揣ɝ���t�+"v���        `��e~Ԯ�ց�t�be#���H+�̝B�IJQ�~vԮ�6Үr��QG�k�8Ҳ�S         f�������Q�j�N��j��E�E�Gy�����l�W{����_�y��ENw[�{�_�(�?1w	        ��U�]�k� b��r���VQ>储��e�v����ib�<�}G��o��ut�xl���]|��[��j�k         f�T�GyѥQ��+#��r��cR�D�o��xI�����W�����o��h��)0f��S����FZ�[�        ���v�=j/{]�'��;�,�(���a�5�S�b�3Xy�Q{ދ"��͝㖖���iɲ�)         =+-^�k� �A��N�����_�Y��.a
��DE�g<'�/�(����n�G������;        ���Q����;&.�(�rA�.�<���a
X?�0�nԮ|EO85w
L���Q�5Q�?%w	        @�(�;!�W_��ιS`Rǟ������S�&�����0j/]G6s���(ʨ=�yQ^tiDJ�k         �WJQ�u~�.�]�\3cGE��7D,�=w
���}��{Qԯ{c���.�)W�tFԞ����K        �QQ��Q>��%0��~K���7D�k��)L�� -�/�/{�w�0��N��s���B        ��W�Q^��(�y|��6i�=�~�"�4w
����ǥ�F�寏����S`�G��^D��;         �Z-j��$ʵ�s����� j/]��]�����ly�_����ϝ���Q�������N        ȧoN�^xMͣr�@6i�yQ�"-?,w
`�ޣ��WF�e���y^�Ȯ8|e�/���        ����F�E��∡�%��N;G���G:��%���{*�啯��ӟ;�Fq؊(�xyD__�        �����^š+r�@�H�s�~�uQ:�;�q��`l�eˣv�uN��*��~J�Ϊ���R����ܛR����E�O���D�O"":�Σ�pJiAJ)u:�2"�GD�(��UU-���>���%�4"v���x����]�{1���#FGs�         L�T�G���9�zj�wVUugJ��EĽq�O���-��`Ji�������e���tv��{�]SJ{D��UU-,�baD�_U��("�<���7'�+^��4�;��]������Ҩ�����vΝ2l���k)��"�+EQ|��noJ)}��ln�����nڵ(���N���X+v|{@D����g���fԞ{u����Ft:�s         �FQF��E����d&�"bSD|9"�RU՗���}۶mw�^������o��zUU�EĲ�(VD��NgeJi "��<i�yQ�b��/��?��;�����G�}E������K�^�͈�lUU7�e��o���ܰaC;WL���IDܶ�q�O����w���oF��)�5UU2e��b��]�1��7�        3OQD�9WF�<*wI��?">SU�g"�ӏ>���k׮}0W̎�y7�x|��Ͽ�]�*:�C:�Κ�8:"�D��y*{�.���W��+_�]?�]�c`������&b���������>X�'���~�;��q����GTUU�r�-+��:����SJ�DD_��Q��(�l��_�i�        �IU>�Qu\�^�hJ�SUU}����4�ͯ�������~}����v۞���몪:9"N���3&���`��#�뮊�{r���w��;E���"v[���ܚR��v��ϭV붔R�;h�v\@����_����=��ÏO)�gE�nY�\y�i�����;w
        ��(�<7��'����F�{RJ��j[�j�C��&êU�������*�|�̓UU��R:;"�̜����{F��ĶW^�Ȗ�9��ݬ(�v�K"�4wI7�zUU7D�߶Z�o掙j�#�#����w]�lٲ�"✈xjD�5�K��=#����g>�;        `B���Dy΅�3���)��E����ؚ;h*�8���W�z�K�����}Wxtָ.��,���$���u�v�~�.V{�s�8b(wF7�?�����F����1���ȍq㷾�������RJώ�u���u���v��1�����o�        ��Ё(/�2"����NJ�c��������_gpp�ΈxKD��_�EQ\DĮYúLZՈ��/����'�S�ܻTyƆ(֝�;��|����m۶�5kָ7��Y�|����7�|�AUU=;"�{�-�}}Q^�򨮽2��~��        `l�^��<�^�]�M�����fsc�n3<<���x�M7�tUD�SUե)��rwu��	�Fy�]����s���0p�B��c��pQ�nю�wWU���V��czA���vD��������Ͽ���Dġ��rK�w��U���5WD����9         ����~�u�v�]�-�o|���zݺu���v�f��������o�yuUUWFē#��[�_y�oEu������N��w��xI�.�]��x8"��n��<22�)wL/�q�~[UU��[N����X��+��Ϣ(��}���N�        �_�(����#�O�쪪�dJ���F�SJU�^�h4>�|�_\V���zVD��ݕMQD�+b���|/w?�������_1�?wIN[��z[Q˛������R�4��5��c"☪�>��)�bp8�'��;        �7*�~Z+�3r�\J�V�u\����q�ĵZ���F���z}iD�."f�I��s�~��#v�9w	?���[EԞ{U�}�.�e[J��;��A�V�ҡ�������捭V블��qk�\�'?5�#��3         ~���:�36����檪Nm6�G5��厙�V�Zuw��|qQ�F�;"b4wS{/��%�G����ܻD��F14�;#���G��j4����4h4�o4������(�|�Un�        t��E�+f���)�K��p�����1�����w����UU�����ɡh��g��`�.�V5�|�y�3r������h4Nh�Z_�3ۤ��f�y�#�<2���Gs7M���(/iD__�        �����F���E�s��%���z�~p��x[J��;h�i�Z�l6����Έ��s�L��"�82wa��߮���eWF��bKUU/����V냹cf��k�>�l6_)����NŒeQ��ٹ3         �Sy�%��;cZUU��v�=�h4^�jժ�r��v�F�}s��="��{�H�iSQ�#��5wɬ7�V�]'��]|�l�B�TD�Z��7��m�c��f�yG��8!"6D�=�{�K�S#���         ��yTǟ�;c:�8�ti��|���Ȧ�1������F���������3m~zpuJ�Kf5���N�b��;c��$".n4�5���ï�l6o]���2]j����]�;        ���n�G���sgL���;��8��h�-�T����l6�h6�'TUuYD<��g:�U�(������{&i��Q{�3sgL��ED��l��E�7�^���f�ynl?��ǹ{�Z�uA�~�
�        �Hi�A��v�]2���F��ԡ����7K)U�V�ϋ�X���3jO�8�~Ksg�Z��z=��\�ח;e��VUu�ƍ�6��;r�0v�f�(���dV1剧��         f��'GZ�ȝ1媪�lUU��V���na솆���q��u��ؖ�gJ��Q�슈Z-wɬd��Ay��Q,Y�;c��YU�ѭV��6�s�0~CCC�ٴi���xeDtr�L��ό����        �,��ņ�rgL�vD�|ӦMA�o�    IDATǴZ���c�6�����:�����=S)-=0ʧ\�;cV2p�fŒeQ�rf��z�>�j���;�ɱ�tMUU�Eďs�L�z=�K~7���        L���ڳ��^�]2��M)��l6_��ܙcxx�31���e*��=%��sg�:V�ө(��g�{��*"^�q��'�Z����1L�V����8����r�L�b�aQ�;9w        0�'����sgL�/���V���p�&_�ټg�ƍ�D��b��t�)ʨ]�E��dV1p�F�ig�~ǖ���i6�/�����l~7�t\Dܐ�e�����H��;        ����=��pQ�)�Rz�֭[׌��l����ٰaC��l�8��Ԉx$w�THK�Ey�3f�i��^��ϝ1U[�ֻs�0=���ÍF�ܪ����2%v�9�g>/w        0������ssgL��]�f͚-�C��F��"����;sʔ(�yZ���ɝ1k�O������G���.�
��n�[�f���!L��R�j����겈��3ي�V#ksg         3Pq��(�FrgL�mUU=��l^�R��az5��ϧ�����s�L��9Q{��"R�]2+�O�b��;"wƤK)}�����Cf�V���񤈘q�+�vqĜ��        �L�?7j<+w�Tx8�tz�����!��h4��n��D��s�L���H�N�����O�]1�RJ��e˖�W�\���-��l6?P���@�ɔv�=���Ν        � �'?5b���Θl�SJ�7��!����{����SJ��2�j�?;�oN���}��gl��p���*���G}���k�>����144�ɢ(��n�L�O���^�3        � �w���ȝ1��O)��h4>�;��jժ��ϟZJ�r�L���Gy�Y�+f<�)���Oɝ1���zO��֬Y�%w�ghh親�N��4r���g�         f���gE��sgL����k4��B�Y�|������D�?�n�L��gG�m��3���*��̈�����#,8```k��W�պ���<!"~��e������3        �V�2�֚���')�S�Ɨs�н�Ν;wCD| wˤ��ŹO�]1��O�t��Q�>&w�d��֭[��|��Gs�������gD�C�[&K��K"
/�        �8E�^��b2m.��F�qs������֭[���R���-��<z]��ɝ1cYkN�ڹO�H)w�d��ܹs�\�f͖�!�f�ycQgF�#�[&CZz`�G��         zP���H��;c�l��3���>�;�ޱf͚-�Z�Ԉ�1wˤH)�Nq�*�S ��t���������800�9w�ghh�_#⢈��n��s.�(��        @/)�(�t^���I)]�l6?�;�޳jժ�����"⛹[&C1�*��W�Θ�ܧ@y��r'L�{RJ��\��ǹC�]�f�xi�I���(���        �!�1���Ϣ��"�te��xo�z���ȽUU=1"���2��N���'Y18�A��Θ[��8��h|;w���l�."�$w�d(�:?����         zAY�r���^U���ƛsw��Z���N�sZD<��e���âX�ȝ1��O���<{F��^UUu����gs�0s<����G�GrwLT�k�(�Y�;        ���'F�s�����6mzN�f����/���U*Ϲ0"��3���$*�GEZz`�	���5�V�ݹ;�Y֭[7�n�Ϗ�;s�LT��FԜ�        �j�^���8���eY>mÆ��!�,�F��"�swLTZ�<����3���$*O;;wUU���6mzE�f����{��xR��mE��{Fq�q�3        �.�֮��ma�RUՆ����s�03mܸ����UΌ7�t�IR�"�A��Θ�璉��.+�����m)�KswLTy�S�R        ����O�]1aUU]�j�n���̵aÆv��>?"���2���#-?,wƌa�>I�S��;a��u:�����=�C����_���2w�D��K�X1�;        �BŪF����Θ�?m�Z�;w3���Ƚ�N炈��2�=�%��a�EQ箘��ҵ���_����Q��~'"���c"���ʝ         t��ԧ�N��oD�sG0{���W��qT���͝1#�O�کO�(z����;��u�#�]V�Z�PJ邈ؚ�e�Ҋ�HK���         �HZz`��̝1�:��ӛ��ùC�]6o�����grw�[QDq�+f��^ew�4�(�>>w�D��,�7l������h4nN)]��c"�S��;        �"�g�N�����1w�Ϻu�FGGG��n���"v��;���OPq��}}�3ƭ��+�����544�ڪ�>��c�����4��        @7�� ����+&��w�q�sG0{���l�������7'�cO�]���'"�(���߄�h6��3w�[J��R�4"��n�Z-����+        �.P�����;c��v:�gmذ��;�٭�l�-">��c���'E��;���O@q��H{/ʝ1^[RJ����!�l6�RU�rw�W��#        ��R���sW�[J��������RJU����x$w˸�(�CrW�4�	(֝�;a�RJ�4�o�ڼy�������Y���sg         ��ˇ�~����5�#�FFFnO)]��c���'�N�i��5o�(�G��oTU�����֭[�HQ���1^�:#        �͊��{hnUU�l��?���7D��[�����=��}��c�Q�������fs[��eCCC����1��1.F        0[��%����Rzw���h��e�fs[J酹;ƥ�/Қ�sW�,�q*�;!w�x}��h|(w�*�v�ʈ�w��E9&w        �A���^=4��N�su��U���#�ù;ƣ<���	=��}Ҿ�#-^�;c<�UUue��uFFFn�����c<���͝         dP�9.w�x���jm��NJ��-w�X��F�wqd�>E��2��V뛹#�7)��U���cU�"����         ����#th��,��玀ߤ�h|#"�W��(���N�I��У��}M�x,7������<*w        0�ʑc#Rʝ1�۱Ղ^�x4w�XG�;�'��Q�dY�E�������l��������ܹs�?��1V��        �*��cr'��=�<��玀Ǫ�l~���w����xI�E����9�c�Fz�������ksG�Xl��7���t���;        �i���-ϝ1�Y�v탹#`,RJ����sw�U��	&+�1*zp��Rz��ի���c5w��?���rw�IJQ��        ��Q�F��;c�~�u��?�c�l6��c�����N�9�c��i�E�3�j4����0������c��s'         Ӡɝ0fUU�ɚ5k����h��o����c��]i�}sg��1H����ㆡ���䎀�j��o��Grw�Eq�@D���        �T�i�H��b�m��No�g���l���������;����Aك���ޜ�&b���w���&wǘ�jQ��]        L������;cL����իWߕ�&���!w�X�G�r'���jN�!�+��S�V��#`�:�Λr7�Uqd�!        x��;4�*��-�#`��������1�#"��rg��ǨX�^ϝ1&)�?�� ���j}5����cQ��n+        ��R��r(wŘTU��������I���c���a+sW���(�l�N����zo��D��0&w��x��        �(�? ������(zk��֭[�?��1iU�m��1p����޽��U�w��|�9	I ��ֻ �V�V��?�Ul�u�^��Z;����3өZ�J��U�h��VE�A�En�!9{�*!@ ����������~�:��|<���z��k�?��~ᙥ&�+V�(�ettteDl-�1���zB        Nzz�6�w�޽���#`�{�;#�K�;&�Ӿö�1p�A��s�*]1!9gOZ1�<���m�=���        ��y�Q�&����a�h��U[��GE:���`�>�ΓZ7R]��g?���0�rΧ�n����        LJO|J�	�t:�/� ��c���Jw-�HG�|�V0pBOa>�t ̄+V���Kw������        �K�|t�Na����|f�t̐VmfS��.��}-�0}�t ̄�R�����$O[       �|��M�i�m�`ީ�]���]����Y�8��P�bh)��+�+�3he选h�Y        ��m�4M�6W0��K�tmDl,�1�t�#-*�1��?��O�-�1��s�N���:���"����x�
        �N���s�1JG�L�9�^�aXiѢHOxR�9���A�#�\:aBRJ�n���R�m���G=6b��        �4H���*�1��ҹ�`��iS�i�6�����JL���zֳ�*3-�|~醡��1�/]        L����"R*�1��iZ5���8���GďJw+=��	s�����<���	q~J)�����k׮�#bO�a�v]G        �}y�a�&bWJ���0����^P�cX�]�oa��@FF#=걥+�ֶW,�d=��Ͻ'"�U�cXnF        0?�����V�X��t̆��������E�������@z�c#F[�ʻwﾴt̢KJ�Ӯ�        �>��^:ah9��l�`�RJED.�1��hQ�G>�tƜf�� Zv��=��;JG�,j�	�)��         �"��<��+&�5+��+V��Kw�e�Yg�� Z��q#bAٳg�ڈ�S�c(���t��JW         S����%KKgk��m�z�#`6�[��m�Fy��?���G�NZJiM��M�{�Δ����J�zl�        `
ڴ)�9�w�q�Jw�,k���Q�)�0��?���\邡5MsE��mMӴ�f�>�t        0�E�B��u:��|���Q:aN3p ��܌��X�bs��m)���զ�        �^�h�RZ_�f۳����F���Ci����}����e���J����RS�f[�����2p       �vkӉ�m�V�tI)5)�kJw#�h�\���>�i���t܈X��\���h�5        ؋C^�`X{�.]���PB�����>��I����t �p�GkKw#=܍        ڬ����
�}�QG�)��gSk�O����<iu]_]�
�T:`(��X�_�
        `2�,�8`y�a�cS3���fS�����}:=�t��:���K7@AחJJ�Zt]        �U:�U۟vl�`����|�zp�9��}_�X�`X�믿���P�����s]        �o�A���s��t��cǎDĠt�P�)��}i���W��u�(%�Ԟ7,o�+�        ��I�g���tڳ��iv�q�"�G;4w����-7�V�{a��|<m        �Ԣ!j�47�n��Z�+4p�7�}9���C�9�\�Jڱc�M���f        �ԖCs#"/[�̮����B����,?�t�PRJ?)� %w�q�"b[�a��G.        p?�%��z�QG�)��V:`Np�7���DZ�銡4M��t����       @K��p�Vl�`���{�l���)�����i�҈�Jg�_B�Y����v<8        ����J˦�/�ԎMa��di�9��}/���	ю/!̬v�(-]         LBZԚ]�M!�eSɮp����e���������hq�        `��H�a�B�]���۵Y�5�{Ӣ�GFFv�n��:�Ξ��h��3        �O��p˜��PZ�4��֦m�g���޴h��snŰfRι7�<Ҟk        ��r�e[��Ԫm�"��1pߛ}XZ�%��ӊ�Ajѵ        �����lS###�847�	��b�7-y�*"����|	a�����=hѵ        ���l�Y����GnϵeV��Mj����Ѧt��4͠t�PFFJ         ��iǮ0�T�n��RJ��FDt�
��W��V��s�M���Rگt�P���         ?՞�M!^Jiq醡���$��Hu{`j՗fN;�nD        �N-�7Mӎ-̠���qhnDk�-���}/r�F����͈/�܎��        �R[v�)�vl�`�����oǵe���M�>,�N�͈�-7���S:        ���nي-̤6mkSݚkˬ2pߋ�<i�s^Z�Jk���=?r       ��k��gY� (�5�6][f���^��.�0���9���Cq#       �vj������rέ������	s���^�ݻK'����K3%�ԊeyO{�-        ���[3po�a�0�ڳ�mϵeV��ͮ�m:i��"V:`(��)]         LB����	�jϰfN;���~��]�+�$�}�ގ!j�^� 3!眢-��1p       �v�֚�{;��0�ڲ���l-�0g��C������P�W\�ЈXT�c(-yp        ��9�r���*%��ڱ�m�ue���K{>4�/ %��~��nV���V        �F-:47RJv�,h9��J7�Mו�f�-:����PR�4��nZ{�        �E۟�iZsh(̄�R;���d�-z*��6nܸ�(�57�7#        h��)��J7@)�W�^����6��}1p߇Ԣ!j]�^'ՖW�DD4-��        �O�6�ўCCa�-Y����j�aܳ��}��NZ�4O*� ����,�0�zqם�+        �I�wl�h���jǦ
f@k6����g�<���!�vk鄉xz� (�J#�~[DӔ�         &�����C+6U0��i��][�Ye�M�>4�,H�����G��J��)        ��j��1�֭;�t��Rj���e�q�*�}H[~ҦӖ[�e�i֚Ͼ        �[�6@)���n�Bڱ+l��[n+]1g��C��#�uG�a=���e�#`��[�����        �m�w:�v�|amܸq��8�t�0�["��s�����'��5�*�-�|L醡���-        ��i��Rzv��m�w�^m�F��zRB;�'����	��P����֮�	        �3ڴ)�9��������sߦ�I	�������f�B�aÆGG��Kw%�hn��t        07��s�a=���G���Y����j�F���[��I)�sN�;`����_)�0�|ۭ;w��         � o�qǖ�C�9[�fK�9��tǰ�M7�N����n,]0����?�t̖N�Ӟ��ܪk	        ��M�/�0�9�����=-".�1�6�]����w�q�ݥ3��s���0[r�/*�0����K'         � ��=���K7�,j͆6߽5b띥3�4��[t�r��7K7�lX�n��qd�ay�
        �|��&����Ǘ��ِs~q醡��ME�?�6�N$���������t^R�a"r��#        ����˜�J7�L۸q��)���Vۮ#%�?��/]0Kr��/3-�Ԟ�������         �A��-{���Z�N��I/���Jw�i�6���l�v�	I)��t̤M�6Ǖ�V��`    IDATsݵMS:        ����MP{���5k������s~Y醉h6�tg�� �n�|����W�Z5Z:fʎ;^�Jw+wS�        `�v�{��E��C��)UU-�����V�zWďo)�1��?��#�UOJ<젃z^��))�?(�0��V��        D����	�RzE��)9�_��CJw�m׏R܇жS]�nF�Kk׮=0"^T�chMM��        D�����)�1/ݸq���#`&84w~2pBӲSJ����r救��ߎ�%�;��o�1b���        �4�۷E��-�3&b�`0xi��n�7o�/"~�t�D����$�b�>�믍���CSJ/+�-��_J7LD��v��        N��]۠�s��W0����w"�!�;��gO4��\��܇������n�	i�濖n��TU������sU�        `��\]:a�^�~���JG�4����l�v�`P:�܇���N����o���?�tL�?��T:bhM�U�KW         3��XE4M錉��u���#`��[����JwLD�خ-rI�CjZ6p��N�4nF��V���?)�1�{߉ؾ�t        0�;�ו���?]�r�H�����-�A7��Z�U�cK�7^��;JgL�ݴi���0Ux��#�Q�;&��        �k-�>������0U�7o�/��g�;&d��o��tEk�+��W�����G�ڵ�U�#`�rί+�0Q�ƪt        0�Z�)�N�s|����[��qD<�t�D�6�b�>m��_�sN�;`���ƞ�T�c"��[#�x}�        `5�}7b�=�3&$��챱�cKw�dݷ�������Nh�	�W��h��������(��Rz}醉����)�        ̤��������M�T������R��zC�V1p���}[�k�,�1a9�7�n��;*�����tהN         fA3���	�R��n����0m���7F��Q:�U�'�^{y��xA��}~���N��h�uj�h�J        �fCy���5�RzS���n���)�_-�1Q���Nh�vG�<�����tƄ����tLDUUO������"��/�        ̆=�#���W�z�_(������hzkKg�������"o�X:c2�SU�o���a��PF�Q��o�N         fQK7C���KG����zIJ��+�1aW�G��^��uZ7��vތ""ޞsN�#��t��cr�/+�1Qy��h��P:        �E��*b����{UU=�t<��s'"�Z�c2굗�Nh%�IȽ������q�����JG��9����#�uc���t        0����{kKWLF�����\7>>�'qt�	���_W����'!o�yC�tƤ�O��jY�ؗ��^�-�1���N         
h�\Z:a��SU��}ٴi�9�w�����ow(��}���.(�0Y����KG�ެY�fiJ�]�;&�[�����        @����o�I�II)}����U;w����xT�ɨW}�tBk�OR������������/?k�����l֫��4�3        ��&�o^T�b��s������"�����n�|����e�>YM���}�bi��c�#��֭[���xC�Ii�6�8        �A������RzcUUO)���R�XD,)�1����z0�OA}i{Ol�9�����a����9wFFF>-�5뻑��R:        (�-�\9^�b��K)}<�J�@DD����������4Q_��ܩ0p��;�D�j}�IK)�4>>�������2"~�t�d5��/�         �m�土WU՟��M)��t�d5�[n/��j�ST_|n鄩8�����`a[�v�c"�]�;&m���l앮         �f|,�[JgLZJ����*���wRD�� �f�7J'����5��"������R�O�n���;X�rΝ����E�A�[&����MS:        ��:���t�T<�i���S��n��#�KwLV��-���Δ�OU�Ds�Y�+�$�����W�������mD��tǤ���I+        ��h.>7򮝥3��UU��t����cSJ'���3�;ܧA}���]:c*��\�r�tGUUϊ������"o�V:        �C��m�\va�)I)�k||��;X8rΝN�sJD<�t�d廷Fs�E�3���gw��[�b�~�#�8�t��ի�Gė"bq�I�ќ���        �T���S��k��7nܿt����#���;����_"��)�1/�O�悳#���S�s~{������o9�dɒOGēJ�LE����[n+�        �E���طJWL�Q���S�#�����s�o,�1%�~�����9��}��wE�U�3���s������K�0UU�����;��>�k�        �9�>���	S�s~e��{m��u���R�rD��n����"tƼa�>��3�1�Θ�C��9s͚5KK�0��z����Q�c���u�o��t        0��뮍��^�)�9�wll�y�;�V�Z�ddd��8�t˔ԃ|�����4ʷ����Θ��x��O�S������s>-"FK�LI�Q��+        ���rjDΥ3�j���\�n��C�?r���lD]�e��K/�������4������~���G�^�-�#�֭[wH]����n���Z��v        `(��k�Y?V:c:<|dd��+���C�z��;SJP�c���������4�[n��I���M�n�/KG�n��B䬈xR�)k����R�
        �EꕧD4M���ݻw��y���J��n�n��"��JwL���s#��R:c�1p���WF̏S�#���n�����Sι�|���E�sJ�L�f��o�~�        �E�n����tƴH)��]w����s*�B;�z��L)}�tǴس;ꯟ^�b^2p���ۣ����eQJ�kcccǖ�]rΩ���E�+J�L�����_(]        �P��S��)�R�OUU}�t����~%��Ո-�2��%b띥3�%�R�K��)�1]��t:獏��(B{�����R���ӥ����?��t        �B���������&��W�n���;h����_�9��J�L��ۢ>���3��}���ۢ>㋥3�ӁMӜ��v�V:�����%�����%o��WO-�        �X}�);��Θ6)��VU����}�n�i�N碈xh��2Xy�|:{�1p�A���D������Д������(��UU��)�7��N�W�q�ݥ3        ��[����JgL��UUuB�殱���RJD�!�[�K���h.9�tƼf�>��:�?�t�t{x�4��z�_.�ܒsNUU�/"�Տ��Û�����        �<P�Vďo)�1ݎ�v���9��!�-���+:��e���-ө>��M]:c^3p�a���l�JgL���/��z/(�ܐsN�^�C���-�mp����t        01��?���v)����z�9ۥ����4�%1�Nn��h�+��j�tƼ�B2�SO�̻���9系��o���U�V-���K�ץ[�[��yc�t        0�4����^_:c&����>�iӦťC(��뽼i��#by�i��G=P���gA��-Q�uZ錙�,�tFUU�.Bk֬9���FJ�J�L�=��>��+        �y���G��U:cڥ��Ӯ]�VUUuh�ʨ��59��#bi��6�ڗ"�������,���2�-7�Θ	#�n���U�V���a�t��',^�xMJ�WK�̄��S"��ǥ3        ���[��ڗJẄ��q����,���Y�r�H���pD��p��pC4�|�tƂ1�>@s�`�O��4�KfDJ�/8��3��:�t3����RJ�"�ɥ[fB���h����        �<V���7\W:c�<��������� U��+���Gq��9��Y�eF4M>uR�`P�d�0p�Ey󷣾���3&�������zz�fF�9UU����FD��W�4u��#��a        `�h�O>1����ه7MsqUUǗa挏�?cϞ=ݜ�K�̔�_�����XP�gY}�g#��^:c&=1"�UU��K�0�6m�t@��;-�}}Ȣ�=3�9�+���H        `in�>���*�1�F#�^����7�_:��UUի��YG�n�)y�m�|������l۵3��pDΥKf�҈�l���Ț5k���a���3w��ٍ��/�2���7��k_*�        , ����G��ΘQ9�W���u�^�J�0uUU-�v����/DĲ�=3&�?yR�];K�,8�4�h.:�tƌK)���ŋ{�n���[���s���5)�+"�)�{fR��c���F���S        ��dϞ|���A钙vT�y����s���-��v�kSJQ�e�5��U�3$�B_�t�[n*�1~>�tEUU�sCj�6<z||���81"�+�3�ꕟ�|���3        �(�p]�_�|�ٰ_D����Ϋ�ꑥc^ι����6�ԋ����i���G}�gKg,Xǥ����k���_D�||����񧖎��S�����`�1���{fC�z}4�Y:        X��sΈf�����7"�^��9�T:��~��#{���9��D���=3�ߏ���yal|�$���-7�`��Jg̚��M�l���͛7���ۨ��#���0����8�tϬ���|��9�.        ������ؾ�t�lyH���^ﲪ��R:����EUU_��U���=����"������{a�ygFs�x�ٴ("�ߺuk566���1�k͚5K��zSD\�R���=�&��|b�;��.        �|��1��Kg̶_���^����V�ZR:�{����ZDl��"b�jܬ�F}�9�3<��r��G���[K�̶�u:�K��:���>�t�B���^�x��M�ֈXP?�sΈ<��t        ��Ӭ[�g�ΘmKs��X�|���n�OrΩt�BUU��z��)M�\?_�g6���O| "��)���\��|����~�^�R���v߱z���c����UU}3����8�t�lk6m��i�+�        ��N�T��n*�Q�cSJ���z�t��g��YH��:���"�ڜ���u{�����q�ݥK�9#_wm4�|�tF)KRJ�dɒ���[֮]{`��l||��UU�l�f,�}��³���?�.]        ��Ճ����w�^���秔zUU�=66���c泍7�_U��q}D�N*���G#�p]��c�>�ԗ�ͥ��(���қGGG���z�]�f���A�IUUO��z_j�檈���X��p��~�Ozg价�N        ط�����QJ���"⥝N�WUթ�֭{R�����eUU����?"N���K7��\tNԗ]X:��1p�c��~4���Kg��s9�.^��ƪ�N��ꑥ�ڬ�����N���sί���oN�x��}�t        ����^�S?U:��ND����ȷ��:���>�tP����?�ۿ�N*���w�>���3�z�:�~?�|�B~���=,�}��uUU}��W�[�r�H����n��&�\��8"FJw�V_xNԗ�_:        `h�gG���3�ND�4�����ս^��+W�\�au��'�z��7Msc�{b�Ç�������.�g��`/���w�)�����/]3,���622�ߪ�꥔N�9��bŊ��暵k�>ftt�"�G��K��%yc/�S>Q:        `���O1z�â��g�N�+��s~����UUuJ���g?��ח��k6o޼�֭[+��9�_�9��MsƮ�1x�[#߹�t	{��9*�|c��=M]:e�9:�����AUU'���=�tPi�6m:���WUUu����O��2n��|�u18�]�O        @;5u>���?��t�\�Ȉ8>��������+7nܸ�O�9�n�{LUU'mݺ�G�2���a��S� '�3�=1W9�}k6T�>u��.�2��t:���ꦈ83"N?�裿�Rʅ�fܪU��x��/���߹s��F����|�����v�N        ���;b��7Ţ�}0��CJ��5��xQJ�E�~WUU�O_�l�GuԶ�q�all쨔���z�W���,�3�N99���Kg� ��f�7�~�c�%�W:e.{\D�:"^�������ܜ�y�~��c�=vެ�����4͋#�7#��s��)�����.��
        ��~z����i���9sՒ�xiJ�;w�����.J)��s>Ŋ7���.UU-���r�/N)�8"�P��꯯��sJg� �[���g#zh�<��S�������_/^�xgUU�L)]�4͚�<�!ՑG��t�����RzND<7����i~�tS���1��?z%        0������w����iѢ�9s��;9�߉���jSJ邈X�����˿�˷��ުU��,_�|E��ؔүEįFĒ�R��h�yQ�+O)���۠i��ĉ���/:�~N�6Y/�9�(�[�n�]UU�s^�9競o����;nP:��+�|�`0xz���9�c"�9q�X��b�wD�ic�        �i�\5��b�5�;b�t��93::UU}/"��Rꦔ�J)]��g>�ґUU-�9?9"��L)+"b?���i�^�O~("��)�U�-�:yO,zݛ"=���5m�_D<�S�#�˗/�SU�5�)"�O)}?�|������뮛�s��z���K�,9,�|xJ���a)�'E���������s����G���n�        ������c����":��9m�Ĉxb��?����UU�W�7�tS�R���]�nx�s�{�t���V�]�l�cGFFK)�s><�=���Ԕ������f�X>����)���d0�������H?���5���������ޠ꺎�˗GUUwD��9�-)�-qw�y[DDJi[D��/�9�RJ��8(�|pJ鐈84"�{O���>=�)��418��h֭.]        0�+.��~��蟿:�&m�<."��[�%K�DUU;"bKDlI)ݞs�3"�望��߷+��E��
#�t@D��'<4"��0;U|�4Wo����QO�y����ٳ'��ys,���Gz�Q�k��#������5L�ٿo�>�_�t4�_\:        `�4�^�E�c����S�e������҇�2���}'��cD����0s�wR�ў�1xϛ�����%07���O��3K�         ̺����g>�4�S`Nh�suNxc�];K�0	�-�w��{��U�S�����'?��g�.        (��蜨?����.�E5�\�{��sG�&���������MwM�(���#��K�         W��$}_D=(�E4��b�79�����n0��I'D����%0�r��g���)         sFs�7c��wD���S`V�����AS�����J���ع#���9���%         sN�~,��S�Y0�K΋�G�����|�41�䇢���MS�fL�sK����ٴ�t
        ���\5�����-��N���s�_�B>���y��}���?+y��+0/���7�.�וN        ��l���r����/�3�X:�if�>5�VG��;��[K���i���[��ӄ         �������n��>۷E���͚KK�0�穼��1x�"��ǥS`ʚ�Ή�{��sG�        ��ɻv��o����K����[�7�.�o_]:�b�>����7�6�+{�S`r�:�/&��hDS��        h������}�    IDAT����J���䍽��o"����)� ��n�=1xϛ���g"��t-�q{�v|�g�t
        ��Q_r^���#߹�t
/���J�������J�0�����ԃ�=�/5-�|������F��ۥS         �|�51����f���)��v��������}i֏��M��|�S`��K΋�;�!b띥S         �|����ƨ��J�ا�Û����E�]S:�Yd�����7�>��.,��ֶ{bp�;���G"�A�        �������gb�wF޾�t��%�E�^���Na���`��];cp��Yߍ�?����Nb�k6m����|��S         �f�[�|�����F�+J����ۢ��?Es�7K�P����������ƪt
U=���_��	�Ǹ        ���w��o���'G�kX���7����ʸ}�s��Bw�i�E�#���>̎�Ûc�O�|�u�S         ���9��ϊ滛b���鑏.]�BQ�>���rDӔ��0kf���t��������'�.b>k�/<'��>�{W�         ~F�������3F^�c�w� b�ܔ��l�vԟ<)�-7�Na�p����7�����y��b��,b���I�3͍�G󩓢�~s�         Ȟ=Q���Ƚ�1�篎�#K1����_���3��οa�ο�4Q_r^4W�����yƊ�E�{vG}��Q���        @�47^͛_#/��y�E,^\:�y�Yߍ�3�y�m�S���٫|ۭ1xϛc�/��4�R:��j6VQ�c����)         LFSG}�W�[��W������h�|�Q���h���t
s��;�^}I��51���o�"bѢ�I�D��-Q�<%�u�K�         0�?����!��~1F��/#=�q��h�� �ύ���G��Q��9����{W�g|1�o]#��K�-]���o���ӣ9����~�         �Y�zC����c�/������e��Nbk֏E}�'"��ǥSh	w��o�aNzWt��1���q��Nb.i�h�\�/|:��J�         0��A����Kb�寊��4��)]��o�Aԧ~2�+{�Shw&����h����y��1�?��G�N�����Ѝ���Gs���k         �M����ODs�y1�ߏα�7t_��m�F��ӣ��MS:�2pgr�&�u����F�������a��{d�*fY�zC��ϑo��t
         �o���������_�c��R�,fQ�r[4g���D4u�Z������\~q4k.���0:���HZ�������>��ͥS         �C��7��wE:�I1��gS:��vǖ���j4���/]�<`����Q_r^ԗ_#��k�y��Fz�cJW1��:�uߊ��3�1l       ����ٓ�����Z=��5� 	� !��#���>��s�R���!�IU�r��s��ԩTrqNm��c�mf4�$@ck�[S��j����a� ���g�We�T�[n(V?�O?�[�O������Daۣ��O�C�}!�XL��=�_��_�5��5l�2p�ޚ���;�G��7���{�����w_ո|f:��ߋʟ�5��R�         jH~�x����5bͺh��?F��ѹ$u�A~�HT^�}d��D�y�ꐁ;#�#����Qx��h���E�/E�R�q������|-����T)u         �l�?*��?E���_�S��(,_���;U)G�����_"?{*uu�����9����E�?+�镟G���uSgq#Y���Qy�/�}�+�RN]        @=�*E��%*��sv<M?�u�{��U*�ه�F��7#��R�� �Y<�Qy��Qy��Qغ-�?�U4����ֶ�e/���"{�ϑ���        ��eY�=��ܳ?
+VE��F���1bͺ�e/���|�������I4w��Ϟ������_��hz�Q|�(l�Q(�NkW�"�|Wd�YϾ�,K]        @�G��]����/
O<�M��aDGg�Ƒe��<�O����EL�R���I�4�7��7��rU4=�r�r~��}!��Evxd�?�l��s���         ��,����Q9�yd--Qx�(���(>�BD{G꺺�_�l��}�N�}�s "ܩ&#�Qy�Qy�k�E��g~p�f�b1u]횜������|فO#��R        �-���������mQ|��(>�r�x:��;u^��*��8��=���0����E��T���ko7������OF�����#V�J]Wݲ,��g"��YϾȏ��*��         �ۙ��l�G���(�X����SQ|��(�x"�ؔ�����c��lߞ���|��:	n������LG�ww���Q)��yk�x:����Ï�N�<��҅�N����퍘�H]         �^�E~�TTΞ�v���eQx�(>�D����G
�+�*M^�?��}��?��;�%�#?�����/QX�>
���#�E�Q�oS}�ǩR���ܗ��Ɏ4h        �!���nd�{�::���#Q|dG��GvD����\`��H�ǏD~�Hd�G~�LD��΂o������E>����Q���\�MD���o���m��F��#u�]��F".�Fv�7�"�x>��#��S�        @���y����쿶),6Ea�}Q�s������k���e��r�}�#?�Ş�҅�O�||,u�S�ԟ�S�?��#"��T1
k�Ea㦈5뢸f]Ě�QX�>bͺ(,�JӚe��G�G��?�>ؿx>�R�.         �Y%�K��_���/���"V���/\��ڟ�]��"��$�1U�bO��Ŧ�?b�?���m�<M,"wC�E�%��+����?߹$
+WE��;�kiDWw��Ft/��Zz���ֶ(��\��ķ�D��E�}�^�������|z*�\��4Q��(MF�&#�����c���DT���         ���RdG{"��?���+#�-���b�����/�Xzm_�����k���-���}��l����'""������|f�ڦpr"�ɿo'"/MF>2quj��P��!�ڭ�W���5        @���#�����s��$z�           �*w           ���;           U��          ��`�          @U0p          �*�          P�          �
�           Tw           ���;           U��          ��`�          @U0p          �*�          P�          �
�           Tw           ���;           U�9u   ��(����%�1�di�,銹�%1��s�m�5�D^,F��%""�Y%���(dY���D��L���F��dtNMD��d�M�����    �wyD�vv�t���A�c��-���c��=�b1*�͑�""��<�,�by>Z�f�uv&Z���}�S�95�s�iS   w��  �Z�m1�f}��Z�WGiŪ��캧�y~.��G�{l8��Ǌ�����    �f�.]c������1�|UL.[���{�1گ��{l8�G�b�p,�3z  ���;  P5�Y�1�7l���bj銈��ޯ^ni����cl���m;#"�ef:V�_��WzcՕ�6suA    ��1��C6����1�o�X��9��3�]1�qKDD�<���Ī���ʅX9x%
�ʂw   �	w   ���)��o��M���[�|�o&�6��;�o˶�۲-""��Gc�����h�ZJ\    Ԛ�ή���`�mz��e|����B������Uq~�SQ,�c���X�{:�����J9i  ��� �$��.�K[��������9�TZ�"N|�q�����Kq��#���(dn4    n�X����C;�����bꢛʚ�cp�ܸ%�=�R��p:6�<]�C��  �d�  ,�������gbd���)w-/bx��1���h������O���|�4    �JT�[�¶�qn��1ױ$u�]+���Ňv�Ňv�ʁ˱���X�w!u  �@� ��G��}ę����u�s�َ%q���̎�c�C��ġh��M�    $Rii�۟��*��;5�vc���ݣC�������tRG  u��  X0yD�o�gv<��R�,����8��sq~��b�ɞx�؁h��I�    ,����8�������(����Y�+Vǁ�~�;�c���c��;  ��� �1�|U}�G1�fC�EQni��;���vƶ��bӉCQ���Y    ��#���G��S/�|{G�E1�|U|闱�+��gD��p�$  �� P5����ܔ:������c��RW�[�����ٝߏ�XL���ʭmq왗���Ď��K�R'}i>"�_��ݵSwQԳ�yx
T�+��% �@����n�O͕�8�V��#��(�V�O�����ɯ�Cl:y8����s���t$+���Φ�+�K
 @5����  hp�yĻe��w���j�}���O���]�S��X�&v���cӉ��v�Ӫx�S	���׍�x�웙  X<�y!z��k�cS%�����rKk�z���ݶ3�/��^^(F�#OD��[c���c]���Iq1+8 �g�  |g���8��+qe�éS�J^(F�O����{�ˆ�S'    ����5q��Wc�{Yꔪ2��^�e��|:��~4�ͦN  j�oY  ��Ҳ���o�~3�]����ƹOGuܵ    ܍��=��θ�6=���(�X�:  �q�  ��vy룱��CL-[�:���b���c��~�m�s    �;Pni�/�2�<��Ȋ&�3ս<v����}���)  @kN   Ԟ��9z��i�mٖ:��޿5v-_O�Ft���    nbr����?�̒��)5%kj�cϼ������F�RI�  ��^  ܕrk[|�����]Kc�/~��7�N    n`d������θ�;������'���w�  ;  p�f�;�ӟ�w1�vCꔚWin����:�6?�:    ����[c�a�=1�vc���oc��+u
  PC� �;2ݵ4>}��1�buꔺ�75��~��L�    D���ǁ�YSSꔺ1�le���oc�{y�  �F�  �UZ�:v����ڵ,uJ�)��s�ę��O]    ����G�~y���^�^����Qr�
  p|U  ��t����'�s��S�ک'���>�:    ҅��SO>�:��͵wħ?���� ��2p  nj��#���b��3uJC8��ѷe[�    h(}[�űￜ:�!8s  ;  pC����m:�*/���6�N   ��0��8�E^(�Ni�]K���&ʭm�S  �*e�  |CV,Ɓ�+V�Ni8y�)���jL�\�:    ����5��G����)uJ�)-_�����  ܀�;  �G�}%��oJ�Ѱ*-���_�\{G�    �Ks����_G��5uJ�Y�1�>�r�  �
�  _ѷe[\z��o�cI|�Ո�/�    �^��8���c�cIꔆwiێ���#�3  �*c)  |�j��8�܏Sg���u����O��    ��rv�3����yZ�<u  PE� ���Ț���������*'�x.F�ݗ:    ����q��gSgp�JsKx闑57�N  ���;  Ǟy)&W�I����q�?�����%    P���;�����`*QmJ�W��_L�  T	_�  1�vc\|hG�nb��+�}���    Pӎ=�b�vv���&.l��6��   ���;  4��X�#ϾQ(�N���<�=�:    j���qe�é3���Ͻ���  @b�  ���o*���H��8�쏢�Ԝ:    jJ^l�#���%5`fIw�~���  @b�  ��f:����gRgp�f:��܎�Sg    @M9���(��f�䉸�ty�   !w  h`Ǟ���{�1g�?�K�Sg    @M�Y��w~?uw!/6��_L�  $d�  jt����ܥ��9�<�-z   �N�~�y�|Ԡ��[bt͆�  @"�  Рθ��f]~��q�;    ��̒������|Kgw>�:  H��  �Ċ�1����|Ky�)�=�T�    �jg{&��YD�ڰ9&V�M�  $�+9  h@�6�PH��wp���b�cI�    �J��qi룩3���<�t�   w  h0�e+b�Rg�eMMq��'Sg    @U:���"knN��w4p��(-[�:  Xd�  �`��x&r��ׅ�rk[�    �*�ֶ��mg��B!��p�;  4w  h �m�ѿ���#�斸����    PU.?�HT�[Rgp��o����3  �Ed�  ����55�����mG�    �*ܞ:�{(+]�  ��  �%v�Ni���X�&u    T��Uk��bu��1g�  �X� �AL._�e+Rg� ��lK�     U�o���zTZ�*���L�  ,w  h��J���۴-��    �X�A�Y��-  4w  h��?�:�2��+&W�M�    IM�^3�]�3X }��q @�0p �0��;���H��ܰ9u    $5�~S��Բ���  ��;  4�!��7���;    ���-�X`��u @#0p ��n�k��߷�!$5�rm�[�n�k*�"�    �=V)�� ���+�,R���-�布Cs  ��� @�+��hy|͆�!�b1�V���/��`   �U�[���^�mF�Ծ�5�o�kʷ�g  �~�  P�*�-_�Z�흋TCJc�y���    �����t�%a��3�����ה�  X8�  P��o3Z_}�[��㷽�    j��m�n_�vqBHnl��/��N�  P�� �ƕn�`gr���	!���|�'os�    T���m��l��1�l�-�vg�  @�3p �7y�����o}�O��o�Λ�|��   �5y���lǒ�o�X��*����E
  ��;  Ը��F3���E��t�oh�Z�    ��nuyCiيE,!�[��FD��  X8�  P�Fo�`'+c���7zS�.�����    �fc���cz���!�َ%�o>wq
  ���  j�Pq�g;3K�F^p��Hfn1p�ּ    Ԩ�[��g�n~&F������9h#�A ��� @������<ܙ^ҵ�1$7}ˁ�ov    �6���N砍�f�#yD%�� @�3p �:�w���\[�"���\��?�n.   �F�����E,�����V��   ���  ��������7���o�`g&"�=�   �F䅘��9�\k��Ɛ��>�3g�  P� �\�ɡ��{�ك�Y!\�   @��"��M.pp�x�o�N�\�  u��  ��ś,�����!��M>�n.   ��]��x�fgbԯ��}; ��`�  u�\^�J|��>+z��h���i7   P�N�d��;m8�|����  ꂯ�  �����7����T�7��ts    5��M���ɲ��袏3Y!��   ���  ԉS7057�}�'�>7   P�.e���o���~��v�ϹK>  �~� @�8z�s1�$(!�}Ώg���   �Z�ōG��AO!��[��L`  �^xu  u�p�����]��!?��P��ü�n.   �N����Fcg�[��>��8�], �n� @���B���5��J9M�4��s~��E    ԉ7���FgbԷ��}ˊ1�m, �nX9 �-    IDAT @�_��K����D%��2;󕿾�b؃    ��`^�+_;������u��g�*no �zb�  udO��?�i��`�Ѵ|��Ξ�h    ���J�W���9hù����̻X @]�
  ��`^�s��[�\�p��9����>    ���]���,������  ꎥ  ԙ���T�^�LXB
S��s~!/����    ԗY!.]w�u�������n�� @��*  ��ǕBT��Ý���Q�]]�H:J_���ʾ�   �>}x�;v\-%,a�eY�_����rD�r
  uǫ|  �3cy!|���,����E,��/n.*G��_�   P��V)F��?����_��T�JDD|^)��� ��X;  @z��k��F��غƯ}�?�=�   �nM�����{l8q���g��gf/  P��� �:t(+D���{��8�f�F��tDD����    Թ7�8k���֙��kX,]_�y��G�� @]�J  �Po�������Ή�'��    �WǲB��]��h��x��?��"K�  ,w  �SfŘ�#���Na�,싈��˾�   �1�1�,lِs�F�|�/&"�c�� @��j  ��l~����D�]-��a,�KY!�f��   �1�ɋq%/�
���v��S���rŞ�  ��  Ա7*M1׆�ԷB�������J���   �0�<⿖����2s2V�V��X^����  u�+~  �c�y�_�M���b�����<;{=�   ������\,H��[�w!^�c6O]  ,$�  �s-�x�|�ت+�?���   @��"���X}�B�R�G���x�l�  �Ϋ~  �ss��3�56�:�4|�7e��   �1�b좁{=��ߏOG9u  ��  ��ʊ��{6u��4�M�    I�s�pt�&Rg�@�z��g.�  ����?  4���1p�W�NǕ��:    ���b����,�7ϜO�   ,w  h�G�#I��x����	    P�9s.u�22'��Sg   ���  ���'R'p�M���p�    �
}CCqux(u���ζ ��� @9y�Dd�r���    ��zNO��=T)��̙ө3  �Ed�  dnn.Ν;�:�{d~~>Ο�`    �w��队�O��=r��٘��M�  ,"w  h0=D��3��=sss�3    �����ŉcGRgp�yGz��   ��;  4���p�\���r��N�    U�hOO����|G������h�  `�� @:t`�[�kܩ�bff:u    T����8}�x���Ç��  ���  ���p\�t1u�R�R�#=�Rg    @U;�s0�,K���t��|���   0p ��s`���3�N�թ��    PծNM��'Rg�-�<�:  H��  ��@��;�:��4??��K�    5���cnn.uw���3148�:  H��  �g{vEy~>uwa���b����    P����#j���\��tw�   !w  h`W�������3�C�##q����    PS�=�#é3�C�퍫SS�3  ��� ��=��N-��<�|�Q�Y�:    jJ�e��O"���)����h?z$u  ���;  4�<���]{�S�N�<���3    �&��řS'Sgpy�ǧ�>��%  ��� ���w+N+�&c�g{Rg    @M����15UJ��M�8z$�����   ���;  {?�C��3��,���ߋ����)    P��fg�o���*4<4{]�  |��  ��/��{/���R�p�}������    P��c���Rgp�����ཷ�R��N  ���;  �ɉ�����3�¥�q�pO�    �+G���Sg��]}����  @1p  �����8~�Hꌆ75U��>x?u    ԥ]}SS���ؑ��{�l�  ���  ����]q���knn.�{�17;�:    ����L���7b�\2}�/��Ow��   ���;  �Y������SN�R���~3FG�S�    @]�w��F����)ghp0�{�Ȳ,u
  P�� �*���������)#˲��o��@__�    hC�����Fnh�h&'&⽷ތ��|�  �J�  75;3o��zLM�R�Խ<�c�'Eﹳ�S    ��\�=�|�A�y�:��M_�o��瘙�N�  T1w  ���NMŻ}#��^M�R��<�}��S'��N   ��t������#�4}�j���_b��B  ��� ������ǘ�O�Rw�,�=�|Gz�N   ��v��P|���"˲�)u�49o���blt4u
  P� �;2U*�z-�R�ԍJ���N�<~,u
    �nr����\.�N��CC����1&'&R�   5��  �c�33���˗.�N�y�������ϥN    �s�Bo����cvf&uJ��r9�z�O133�:  �!�  �])���{o�gN�L�R�&&���?����S    �������O�R�N�8��z��ϧN  j��;  pײ,��?x?>���({8qW.�?����K�    ����h��?Ĺ3�S�Ԕr��?�0v}�AdY�:  �Aͩ  ��u������g�b���9U�R�ľ�?�c�{R�     wh~~.>|�ݸ|�b<��K��lfq+�c���{����h�  ����  �N&�������<�|<�cgꜪ411��N���N    ��3�N���`��'?��+V�ΩJgN��=�>���  �wf�  |g�J%>��I��]���bttv�N�
Y��ўCq��~u    �ƍ�����c<�����vD�XL�TJ���ٞ]q��|�  �N�  �̅�����x���b�#ۣP(�NJ�����t��1>6�:�ѓb2�P��� ,�]�b��f�����=�b����=����3�_�+W�NJ�R�đ�Cq���(�˩s  �:R���uy�  ��<��^���V�Z�����v���)�jzz:�}�'Μ:�:    X@�B!�>�-�~�����H������ĞO>r���3��?�}3 @#0p hi�x�{OǪիS�,�ٙ�8v�p;����s    �E����w>���mm�s���`��{{S�Ѐ� ��; @�0p'����œO=�7ޗ:垚���G�Ʊ#=177�:    H���%�=�h�|�����L�sO��ő�Cq��|���; @�0p h�T�������{*6l�/
�B�o�T���=����Q.;P    �inn�m�<�w>]]ݩs��<����K�sp����w �b� � ܩ6K�.��~$|�����H�sG�,�Kz�ԉ�q����s�R    7V,c���bۣ����7E�XL�tG����̩q��񘜘H�_2p h�  ���jU(c���e냱y���֖:�+�,���+q����=.fgfR'    5���=6oy �l}0֮[�*����ą��q���Y��N�o0p h�  ���ZP(c͚5��M�a�}�jժ$�MM�����|�b�]������     ԧֶ�ظ��x��X�act.Y��y����p\�t).]��C�F�T=w ��a� � ܩE�--�f��X�vm�X�2��X�K�F�P�gcvf&FF�c|t4��c��?��J���    p+K�tŚu�b��5�|��X�be���߳��eQ*M���H������@Dy~��}X�  ��9u   �͔�����Kq��/���)�����{ituuE{{G���Gk[[���E!"�MMQ,�|@37?�ss1;333�155��ɘ*�bff:��    ��;JN�)Ź3�������X�����ѹdɗ�-������.ɲ,�J%򈘝��ٙ��������(MNF�4��ɨT*�~w   w��  �)�J%���b|l,u
    ���������L�  �芩            ��          �*a�          @U0p          �*�          P�          �
�           Tw           ���;           U��          ��`�          @U0p          �*�          P�          �
�           Tw           ���;           U��          ��М: ���:6�ʢ~̙����^ԏy7֗ƣ�g�3�����-moI�       T�ߏ^�����zf�[b��kQ?���P�B��΀�������fRL��O#5���qlf~Q?fwww<�nŢ~̻��ž(�˩3��mli2p       ��_ǧ�����z�.][�V����ˑe.�hm6p��S           @��;           U��          ��`�          @U0p          �*�          P�          �
�           Tw           ���;           U��          ��`�          @U0p          �*�          P�          �
�           Tw           ���;           U��          ��`�          @U0p          �*�          P�   ���%�������=��_���MhҤ�{h��)�Rڌ2J/)Yt`ņ��a� �"BHl*6��Z�%* ZڊVC�J!iQƹ��̌=3��>>�簨 ��i�w<�?�<�.�����o.��'       �Ъ{ ����'b�Su�ؓV�����0r�����~��{2�����W�      �>�~�B��cO�=cO�'�������3u�ؓ�kq����܄�� i6�7}�� ܂A�����n��	       ���xO��O��:5;ݺ'�c4�            w           ��          ���          ��           � p           �;           )�����������=���^t�J_3�j�F�7�Jϳ��~t��!.*��jEQԽ       r�N��n��I�$ԋ�։T�ch����_��Y��j�z����J_������x��f'V{���w�c�+�1�E���bfz��       �.��|��7���Ʒ*�NkIc}`���z'�wʷN۱�9Z�3�:�&'��m֨{            D������磈�����v\�v����f#>�ܯT��~��ra��4��z��Oƙ��*}���f��r�����XX���i��=�V����X��[�       ���(��g��������^��d���_�t�?�������� �Qx���c�P��+��X\]-}�(�XX��V������f�[��b�������	��ܣ�=E1���ҥK�{�|��SSS���|��S�'!pr9��Õ�g���q����狢�G��U��      �BQ4�����ŋ���X����t��ir���;�̝=R�yvhi)VΝ+}��l�����H��           !p           	�;           )�          HA�          @
w           R�          �B��  �抈ߚ��=�mzsGb�#g��m4u�'�5w��     ��nn����gp-|��hm\�{��|�ۊ�A�+  ���  �ъA���뿞v�'c�����mt�ر����{    @)�v;����{��{���1���>$��  �\��           !p           	�;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
��  @fWVV�o^���gp=~<f��=    ����z����=����{kqWQ�
  �K�  ?F�ۍ����g      į�{<bJ�  7Ө{            D�          HB�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          �Zu`��O�3�SQԼ        �f��s���(|�+ �����=���~�
w         ���C17{(�:������ֵ�~��n;�&��O4z�_z��%;��� F��J����Z��e����wU��i��      @YE�=yw�һ�ɢ[�u��T\0��Z��ի����F���^W�t���܅ů��c��϶�����*}�b�J�E �7��G矿T�|㾻�س�tǅŋUg      ��4ҵN���|�+}�be��"���՟E�������{��3�*�qa񭪳c��           @��          �$�           � p           �;           )�          HA�          @
w           R�          ���          ��           �Ъ{ ��웗�/�m�3��?�{@-���      ��8��������b�랱'Ůgxf��������=�[�      �8)v�'د<��F�            B�          @w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )��    IDAT�          HA�          @
w           R�          ���          ��           �Ъ{ ��3�1?1����M����U|xf"�f�3`�-L�       ���f&���6��ܭ�Ss�Quπ�v�։d��{��nn�to	G�^         ���<q���3�NG�^ @2���k           �	�;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          �B���W�vz��Fzg�hĕF���~7��h�� ow�d3�h�=2       ���w��Z����݉��0�~r�ǴN$���ZP��u=^����Çǽ�.���*^~����zuπ����G�SG��       $��X쌶�9r�H�sO��饗^�~�_�k�[8g��{��n          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )����}�h�|���g�Is�_�N�3 Fn��w��O��{ƞ��;1����{       ��։;b��}��|����?[w����{ƞL����o~��܄�� ��Mǵ�{ƞ�����X����������      �R�s���=�z[���Α�����.pO�Q�            ��          ���          ��           � p           �;           )�          HA�          @
��0zKV��ko�=㆚�n|��V�������[��v7v��o��W����Up�g�����g       @��t9^{�R�3n����Tl�ֵN@Bg�;��/;�߸W��N?��11!�>h�C��N��m�=��^�z����7�P���F�+�g��n�g�n߿L      �C���}��j�t+�NU>,`T�w��N��;q=ɳ��!=��c����0�{�^t:;�Ϸ��o�d�;��w_���Vu�P�x��x��J��(��P�C�ggg*�*��w���Dtw6cg��      ��E��|t�wt����)�:MDﻫ|1񥿏Xߨ:`��{<>y���o���E��L�²wv���1�jj����{�S�EQ�!SѥK������OMM��g��tǟ~��H�3��ӟ�L�����q����狢�S�N�ʴ�֯.���w�z       �Q���s�<�;.^������OOO��ӧ+��G_�w�;���.N�ӥ�/--Źs�J�o6���O�ʴ��V_�+��Q�            ��          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          �ػ��ּ.��������ޗus��@�F���k��kVH$h4Q� Ĉ(	
�1�(`1�A��`0��E%1pg��˼����O��w�t����#{��鞪��z�:�����Ϸ��:�T��y���          @�          Ȃ�;           YPp           �  @�z��K�������<����f���M&K�4uQW�{ro��8���*�o��B�z.��4MDU��ٽ�����Zu���=gn>z�#i�2ƽ�}Ѽ���iƿ����1����?G����׻ь}��Eo�9bM]=���{����s�{�Ѽ����s1Ϸ�{�������s�\7%M���3�e  ��?�  ��w/����7S�`���w��7}K�3a�����c=��~��	�i�������p_ϝ�گ�����N�N������;�s>�S?G����P��^����g���>��g6PKU��Q���9�}������	%j�˟���7�빇�?G�z��O�r<���������-���gJ�.��������޾����<��ğ:�D��ܻ����c=��;�����_�P�v���?�n�����c��~�'j�������z�;������\ۿ�������s��S��~�`�T���*������O|.^��0�D�QݿW>���zn�C�C?���������~�s�c   dŴt           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           �0}G�~ >���c         ��CG_�O��z���
 ]���A��h������%        ��7^�p����� �CLk           Vp︵ӿ����4o�G~�|�;��3c�w�ʸ� &���;�������wފ7��ύu�����i����       0QM3��ɛx�h3�����w��X��ݼ>n,��k~�'c�W��ȏ���Ǜ_�g�:���Pp︺.SGxB��"�6�{R�d��Gl�1�h�hDTc���{<       ̲�����}u�0����1��(t�����            B�          �L(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,,���y���x��:��U� I��~w����2u       f���w|O0�^�قs�`�:{Ppo������Z� �á-�p       ���� ����v��N��K            "�          Ȅ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,,� /�H/�H�7�c.DD]�S=�8�z1?�	�$�A       �K��t��đ^/j=Hj�[��(�3�~���9py;�qG���&        ����;�NO�ʏ�N @f�R   �[��[�#̄j�f���M�n��M��ͣ��1xcxt����x���F4U�:�L(où�֝�GQ�^O�]��2��ޝ�   �(w   ����^�3������E�k3���)[��h��
���X�(��1�Wo>���K�c���V/�Kc&>;d���h�%c8W��h|�   w   �����k��O��](B��d�|gNDS�S�Ȟ�U������1��_<Qשc����+�l�����1؅{��'SG`��F��  @*
�   L�տ�ox�\ԛS�`��Qom�����*cpj%uvS�Qx}��Xv��Y���\ʧy3a��J�Y����Wע���:�(�]������\  @
�   L�����>H#k;�"Yk�*�S˩cdm�z:�G۩c��ʽ5�a�O����&�|&�M9��Ldɛ���V�X���^�עZ��:   ��  �t5�mڟC�'�*{3��g�8��`�:{(�ߋ���1�U�<�����1�Cu�N��.���5� ��7
�g2�ތa   RRp  `�|I��b�x�<G����By:{��K�Te��*����՛cp�b���\�����s�l��zk3�Χ��s(���D��obo}c  ���  �:����_�jc=u��8iu�]٥a&X�yoJ��A�rw��lP��]�.3A�uw坍^��:�1�p6���1��^  ���  ��b�T4E?u�,Y�o64�aVO������Ũ��K�(�<[SUQ�\J�(q�Nqz6��۝1<�����F͆�����g��ߋ��˩c   �a
�   L]S�r9u�,)���ճ���]f�UW�MYov�����������J��`x�JTw6R�Ȓ�fCSU���pO<;|�{��ұ��I  �Sp   	+?[��eV(B<��gG�J+��=;���(o�H#;řvʙ!��Ok�"
;����g��nf���l�O   ���  @�D~Zu�N��l>+���h�*u�옼2;��cx�R��Q�-�E��)�f�U���?�Q��c0"��Vom�����1���J4�A��1y  ���  H�8�M9L#+
i���ފ��s�cd��u#����c0�ʧ'SG`�b�S
��b�秙,7[����_>Qשc0�f8���J�Y���bx�l�   t��;   I4���=�:FV�yf�b哬�7{�V����Z�w6R�`�;_����b��,^:����1�bE����Q�R���h4{|�{Rq�ne   ���  @2V~�2��Q�|����1��d'��3��ս��cdcp���1)�	MU�@Yz�(t?�����=��  �(�  ��2��l>�|��$�VfOy�F��7S�Ȇ��j�(V��N�+��&���Ξ���v���=���������1�˟�  @�  H��􅈺N#Ŋ/�gQu�v��.�������^��:�P(u���l�������_���!פ�T���*S��Bqz%��0u�d�����0��'R�    w   ҩ7*��?
i�ˊ������4�c���c���(o\K�}P�}���l����觎�VfS��(�畃#"���RG`�|&�8��`�:   (�  �V�����3�!3�g���c���kpn5�G۩c$W^�՝��1؇�Fqj%u���&���S�O�s?1�
�]DD>�  �	w   �R x����-�g��cVP�]õ�Qݿ�:Fr����j�2��S�H��h�2�`ףY�s��Ѭ�/�#Ux/  �w   ��/��:Br� �m�kV̭w���j��W�Dqb1u��yf��OAz��v�u��v�u��{Q^��:FRMUEqr)u   �w   �6֣\��:FRV��}]��~pr)��L���1\om�����1x��v�u��Kє��1�R�m���1���:FR>�;�����F���:   D��;   �z��_��A�W5�g_�X�I��E�u�����rD�݉6���1�v%u^��P|&h��O6�h4�:?�;��  �w   ��r9���ǥ<f��b�� ��op�Lԏ�S�H��}MQD�z2u�d��_�ڢ�o�:�C�w�h�(V��N����:  �w   ����׶ o���Qo>L#�����J����*c���Q����:v�^�M������?H��_��0�+kQݻ�:/hx�jT�R�H�8��:   |��;   ��.Fu�^�IX5�%�:�+�,gNDS�S�� t�X�E�;��w�t�����Dڢ��^DӤ��D�'��Iy�FgW���5�m�]����坍�1   ���  H�i:�R�2O{]=�o�F��bV��RDY����/�QשcL]���K�S�� ������1��A{t�~���D�6�   ��  @�Z��j����Z�j���Z�.������6c���wW��m�_��9����6��=����  �<(�  ��.��8�b�6�9M�Oc��:�+&i�ESQ��Lc��V\m�.���ڥ�cx����I����u���(o^O�2�x.�͇�cL��	   r��  @���~��:�T�@n��Fqj%u��^:���G�um7��*cб�m�uqW���oۮ��n�Sg�Q��.Fu�^�S��2M���SLUu{=��R�   �'(�  ��.��yڧk單��]е�t�z:�G�cp���n��@]�    IDAT���f��z��7Sǘ*�>[�i��X9��;/�]�a   r��  @6�V��ڗ�]еb�1�>���"�:u���wp��+�l�����1��r)�,S���u��]�<���3�cp�����K�ٮ���(]�  ��)�  ��.l�N��K�T�)v�����f.�Ocj�V^ꊢC��.�;uI���]�w�.�����]H�6X=M�Ocj��  �٠�  @6��
���۩K���]���F�L@g
.Mŉ��)��.]c��JrWtiw�.���dp�Lԏ�Sǘ��c��tES�r9u��0I  �\)�  ���(��z2u��P�i���X٥���+���څ���K�	��5���t�|�5õ�Qݻ�:�TtiBJ�4U�S�8?��թ�u&i   �!w   �Rt��֕/˻�+��*���y�W^]��;LVOG��(u&�#;L4�0�S+�c0!]�lԕϯ]�s   ���  @V���-�ۭ��^DӤ�1q])-uQyg#�ׯ��1q�p�u�ܕ�������h�~�LH>�ui�.*N,ESSǘ8�4   ȕ�;   Y����]���~p?��/��1Q���Q^��:Tt�Xم߱˺P�����e]�e����߱ˊS���]�\�(��1�����s��cLTS�M�    [
�   d���wa5î�/Ka��|�~m?O�7�G�~3u&��c8��+|w��왨m��1Q�]Z�)���8ۅ�(]��׸�$   ��  @vZ�%r�?�_ 7�ۯ����7�p6���1&f�v!�R�`��������1&������:��{b�Z��q���  �lSp   ;m.B4E?��S�c0a��wSG����E"�k�����:�����TU-.���)���|O<�t>�͇�c0am^���$���1����{M�:�Ĵ��  �lSp   ;m^Y���Pm�G�~3u�����bx�\�LA��u�|��}m.��w�}m>W�|��/���Rǘ���3Q?�N�	�܏����1&�$   r��  @v���Q޼�:�D��;��Z+��-*񤶎����^YK�)h�����.(N-�vbd���O�Wom�����1&���I<�����SQ�<J   v��  @�ںb�-�����������z��/}!�iR�`
�����c������o���4E����1&�X9�:SR��~���Ok�纖�  hw   ���"�-�������^8��f�N!�;��0-,�������w�^���z�LI+��&���S0%��wSG����  hw   ���"�-��e�v1�{wS�8Pm-��lMUEqb)u���-m,o���-E'̵q"+�k�$��系jc=����c����   �Sp   K�+k�+�uEov������c0Em�lT�<�����c0E�,��}����ǣ���1Tۮ-쭺{;��WR�8P>�uOۮ��K�~� u   ؓ�;   yj�(Vڵ�cW�eom[e��EQ�ֺ1|b1��L�)j[9��/�W/����[�Q�]H�@�'��nwO�^��  h'w   �ժ/�m�Im+��=�H�WZ�jawN��Ë�R�80��cM�:S�Ӣrpu�N��L�蚶��߶{|��m���\  �,Pp   [m*B�.���g�D�h;u��TU��S�`ʚ�0��+�c�6]W]Ѣ�L��6+�*��M��jc=����c0eõ�Qݻ�:Ɓ�l�<   �I�  �lϯ��\,K����AKJ���Qom��A�Y��,�8}"u
h�Ć6�.�nТRxk�)�ex�JTw6R�8��wSG �����b���q-��[�c   �s)�  �����8��:Ɓ�Zew��W�쮶����J4E?uh����bx�l�$P�و�+�c��Ֆ(�rMa|���D�<  ��XH    �r�s�:�~��S�xa;����Hd���k/_L�VO��@"��/��?���c���Ƶ�H��{;���ߏ��l�;��|MU��A"��Gb�#M�/�K�D����b�w?�:����{Wm�ףZ��:��,  ������  �z�sgbp�L��o��zl���L��)��03����������E�:���1�t!uط��m��   0Es�           @��;           �Pp           
�           dA�          �,(�          �w           ���          @�          ��B� ����{q�N���|����'>1�c�c��jTe�:t��y4���K�c        �;kw��`���W>�j����S=�8.�9u]����Co��U׉|(�3��M;u3�c.D��\� ��&�)�M�'���        �]�C�w�i�n��u��JoA2��U          �NQp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���: �|������c��^Y�ы�R� ���_�G��s��������      ��=9����J<z룩c����0^�t#uv���"��?W��өc������;�I;o�6���C[�|p      `$;o|d��'��=9�M�o}4���9���M��ͥ            
�           dB�          �,(�          �w           ���          @�          Ȃ�;           YXH��{+��硫�L�Al?���Gu=�4 ��6(����;���zu��F���X:4�:       ĝ�c����1�ia���1�N���P���8f�i����Ȥ���_�X��uj��wo3Ξ��:�3͕e�������A/�F?�w��A&��O����;       Y�{o+߮�`w܁X+ʱ
�����0�s�'��M�Rp�C�G/z=Fӌ~S677G^}u����,"�*�@^�#��2��W>����d����bn~!����q~       ���1��:Eo����"��]<���#�u�j]'&L����{~xb'�������p��ȏ?r�H|��Ʊ��[���q�̸� &�k��{�۾��F~��7�رc#?���ŧ?���D�潋q���D�       ����������1nݺ/^��/��r|Ï}�X����~6�^�4f2���K�����|f��_�z5�?>������S���~������q���D���̥            
�           dB�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           da!u   ��q����1f��&u�e�i�cx$�ы:u�2׋��1<����Q�<�+�7��y?u��Uۛ�0u�����\�\��Vx���H9�#��H�^/��!x�\�xT;��~�<C�Ѡ�v�   �Qp  �/}�x�����1f���9E�z���1<��!��!x����1<��+��3u�OU�}�écd�?7����|�W�K�S��^ugC�=S���k�'F�9?�:�p�嗌�~㿥��3�����=�|Q�  �K̥            
�           dB�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @R  `:�u���I�bo�S      蠿�P�0u��X�N  ��(� t�7�ש#      ��oZ�=  ��K            "�          Ȅ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          ��B� L���|�����1         ��]�����Q �)Qp�w�~#�y�������        ��'�y3>�Λ�N �!s�           @��;o�ڱ���f7�x�՝��Pn�������ѻ�>n,���_��7F~��^��>���q�ظ��2lM��      �Țf�ߓ�x���ȏ?<���t� &�w~3k#?|��/�ko��u�Eo���A�9џ�t)�w���k?ơ1��e?��������	�Y=խ��?��?���׌u���L    ��e�΃,�����2+3k�꽻��VK�VK�}C���-�%˒ !F���cc���0��L�f��d �e	ہ����8d�`kDWu.���{e확y����ѠV��|���w���gwf�oV�{߽�~�9  ��k��}u�Z��w����z�uP흎������������5�]�3M6�:            D(�          �	w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          ����X;c7������1Ve�l�� �����П�7,��#       0$�nxN0�&懿�4vc)u�@��F6]����WS� `6_��      @cxN0����[�]L�M            "�          Ȅ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          ����`�~��{�F�Z��l��ƥ��5��?�|G�T��o��RG        2�wwu�:#�q%��c��H��p��u"3
���6�ƽD���m        ��kt�n6>�: �M            "�          Ȅ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,�� ���sq��]���Ll�����k�c���1Z�RǀF�����m[&R�        2�_��s������u�~�\�TU��h��oK�y�x��u
���-�b_�^��ܾ}<�ܺm]_������t:�c@��g�D�-u        +�m�G�����s�D�"��<VF�g1OH�}�6F(�����            B�          �L(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YK    7��wc!u��Ue�7R��:���e�\�K�[��^��������d�{�j��F�����ݴϝI���?��I#{���RG�6�s�떥׋ʿS����-W�ʥ�����Bt/_���SG�^���&   ��',   ߤ�y>�ۺ-u��-ퟍ��J�[(�L���M��w�[����C�cp݅��?O=�:J���]�#p������7����rv*un��w:�}ǟO#{������bzw�������ѽ~-un�u�`DU���d��v�5;�:�P�[�>q46����d��ޝ:  @vFS   �Mk���Z��wS*Uf�*�(�M#{��dT�n��F��]��s�H��F1�}r9\O䫘r^�z��'�G����1��+_U�k"�2�����b�܆	�wW���:`�  �7Sp  �&U��ޙ�1�gu�d3�&    IDAT�)[�]��(k�wWL?o�F�Z��wսz%ڧN���m�������1�W�<�:�SU�>���+o&ݝ{߼�wW�N[h  ��  nA��Ϊn'Z&d�C��o�7���^��Υ�h�9�:F���]U�:�SUQ(�Q�̩��]H�;0)��\s������yk�NE�i����b��   ���  p�ޙ-��WN���R�Ȗ-��׽|1:���|'ޫ�W*Vޑ1�?+;ߙc<�1|G�3'�{i.u��;ce�;�SC�zK��:t u�����  nI�  �ʙ��vR�Ȗ-��כ���GR�Ȗ-������Ue��=�cp��wVLZ�2w-��;r��u�@�o���-�Z����h�滭ֱ�ѻ~-u��d�۫��(g�R�   ��X� ��jt4���'���Pڦh�:��G���RI����b���׼.u�,)B�rjWL���1�T��1��]��CK#K��鈎�X��~y{���h9�:wQ�UY���M��d�1���ۉ������w���%��C1�+6��cdIqz8ӻ�O~:u�,����99��rgІ{t�78�}��R�X���"^���L`��?�3N|�c����b<��~;u�5UL�Rp�[��bjwl��'S�ȒB�p(���nǪ�ás�xt.����������ӎbv:6�����d�{�JtN�H�e(�v+�߆k��PL�?�:E����PL�����Q�c�@���/�|O��2>��|�sr�y����8���JcU6^�����;�cp��   �ʃ�[k?b�!� {kU�����d�}�dt/ͥ��%�Qã�3�:B����au�[+��{��G�\�Z����9�:�P��M#KŌ�aлv5�Ǐ����¤n  ��Rp  ��rz���-�V�݋�s�t��i9����1X&%؛U�N�L��1|K���P��5���(�NGt��͊I��aѻ��#S��N����^8�:�T����  �H�  �6�W�D����1��l:\�Xy3�&����f�����x#u���Y�nG�w&u���3U��:Fv�ã*�(̦��cx��lt3cx��,�f�ǣ{�r�   �Rp  �Lof��q3+��ᛕ�M��]#n��7U��:�TK�:�?u��XMy����Y�>a�����{��RL�a��q�  pg
�   w��KuΝ���Q��Y�g2u��>v8z��S�Ȋ2�p���(g�R�Ȋ1<|�i�ߨ�3U��:}P"|���|��N�>X��f�u�Kw�BtΟM#+>s  �3w  �;P�x)�ç}�-��A����\�K�~�zQ̘��uUe��RJ{)�����/�>���^/u�l�ϛ�1d�W.E���1�ѽz%ڧ�{׀/UL>�:  @��  �s�Lt.�K#V�BUe��o��6�Jc���Ǐ��2���U�n�{�h?l��]����1=|z�Ѳb���é��w�c��sU�:}2a�EV�  �;w  ��P�~�ե����/�b�p21�E&��r�LT�V�Yh9����1�So�z�OK#U��=�c��'^��b8��y�{���^�EŔ��   �f,u �_Q�bq)�jcE�;�m�ٱB���^_糅���.0���{ϖ5�S�c�>�:Fr� ^�/2ae8���DU1�qS�(�)���ݎ��=��oM%��yxhS�����J#��>V�U9�+�;?�:FrUYF��l���{���N�Ǣ{�rl����Q�s_п�h�b�����R�]�����k}v��/��u�o��I�5���@��\��}'SǸ��N'�^]��{�vm��gr�K��ߔ�#����������زyc� Y)=8��?*���u(��j��۶���T��h�9�:+��D�w&6����$�=ixӻ��f������O����Ië�t���(�NG�n���
�Ϝ��܅���é�$ջ��#S�`%�*ʙ�c˷���I���;@�N�������h��}v���� ���7Zq���.fqr.�g�u���56N�����<+  �]�����k�c$gu��Uu�Q�N#9cx�Y�1�;w!:Υ��
�/(g&SG`��^�X^�Ks&;�1<�ʙ�SGH��3U��Rɇ�b����>q,u  ��Y���>��?�ۚ�ڵ�q�e���X����t_��~�'�����F��~���#�ಿ��+1{�H_����O�kYvܳ5FGGbq�l\�th �0t�h����}_�$I)B�bjwl~�{S�H��6���	
�����*�3/��F6lH%���ѹ4�:+ԝ���gc쑝�����E�g*u
V����/{,u��\S�bzWl�Sߑ:FR��p���}�ֳC9�J����ǿ�G�W�^����~�qb"���o��5~���Z\9s��h �����g?��e��������6GFG�W�j%����[cdd$n\?�/�k����ѝO����
��.��k����7ƃ�|u_�1�iS�� n�Ï�u>ko:g�����H�|�+��l��J� ߨ����{oi1ڇm>̔�!�]kv*�n'F64��,cx��n,D�衘x��Q�)&��bjWl�����L����-̧��*S�b۟�H��T�N���4Ԗ����r�C��x#F�lM%��}�*�9���q���e��͛��:m���o,�����}�ϊ�1q~��6l�0�sx�te�?��5�:   �0(��K!�r������1X�rv:�V+u�dz��:v8uV����CR�H���EuPN7��b7����BVӏ�:h�d�����[\~Q���������1����(��I�U���(g��Ja�  ��(�  ,C����--���LӋ uP������"@1���5PN6��ݻv5�'����*5��<��^�j�1\�Sǣsi�+��Mi�^/���S�H�����u��	sU����S�   

�   ���V�3�c$c�z(\,TH��F����U�:���	c�Ks�>s*uV�}�Xt�\N#�b����:)�L���L������6&��C��𞩨:��1   ���;  �25�`��h�C��J��%料�M����9�:F-��z��(�rp����6x��:i�uaU5��_'����ɂuR��̒��:  ��Sp  X��n���7UY���(g&��vS�XwUYFy`6u�@���h�8�:FM}��b����n0���bVS��:j����ށ�NZ�FU�c���ۍrv*u�@�jEk3Rp_  �|
�   �T왌�tR�XwM-1�Q��B��Lcݕ{�y��UK����hܟ:k���J���hj1���n�����|�뮉�PuUu�Q�Ic�5�ح�&��_u�Q�N��  04�  ��*�(�
�2O�4q1\/e��٩��&i�E���poa>Z����i:���c��&�uUu�/L�l�&�I묉�8M���lछ��   �R
�   }h\��׋r�-�뤉��*����������zi�>�Ks�c��bzwD��:k��v��m��a���h�>�:k���M���f�����uV�LF�����a  ��(�  ��i+��l^;M+BT�N��Bg�u/��΅s�c�����4A����p�4��UL�uӴ���x�Tw�٩�:��1�U�g2u�Poa>�G����\  �G�  �e�V ��~�W.E����1�M�Ё�-�H�5֨H;�(�ΤN�k��k���Mд1ܴ߷	���Z��1�Mw�����b�HcݴO�N�v�i�r�A׈�^3ϧN  0T�  ��[��ֱéc��F�H�I+��Ԩ1�OTe�:k�Ie��,�<0�:k��;U�9+7�m��ݎV��M&�S��u���6I�&��������1   ���;  @�U���x5�!r��VK�t��p��s��u�P��S�X��TD��:k�j�S�-�G�A\��I�M�vj�&��4�wm�&���&��  ���  Ч�!���� ��ƬBZUQ����ǏF���1�ES�s�׋�!�Ȭ�Z_M)�3�Qu��c0 My��]���R�` ���U�:ƺh�$�&�^��3'S�X&  �O�  �O�)�4��l���Sѝ��:���O��˩c0M��Рt5�Xi���j�n���DM��PL�jL	�i�2y�{�BtΞN�)��y�36  ��)�  ��{�B�ϜJcଐVoM(Z!�ޚ0�[GEo�z�H&�U�N��Τ�����7�\�c��z��>z(u��k�5S�5��g�ք�o�����!  �o
�   +P6�$P6�!c�5a5R+��[�QMx�i�r�LTe�:�@�����1���|��Nc��v;ZfS�`���^ۄk�&k�=��F�ֈ�p~G  �APp  X���0չ4׈Uꛬ	%���M�:����Yc��:�(�ջ8ۄUe��rv:�V+u��ﵽ��h:�:����RG8�4�	�����  `P�  V����V�?"ZGEo�z�ӝ���gS�`��n'Z{gR�����QL=�:�@5aU٦�{a���(��-�LF��� u�.D�¹�1�7=ZǏ����������5   ���  ��SǣS����� U���S�BZ35^9�	+R�2OUE�g2u
����5c��Q""�{�btΜLc`��f��
����^/u�ΟAu/_����c   %w  ��sik��e%^P�UW����/�P{u^Y�}�ht�^I��s9��v��W�BxA���|�ϋ�=�����:e  ���;  �
�u5���|��N�uP�1Q��3/*f�":�,+�5Coi1ڇ��1v�h���ڇDoa>u�A1Y��U��=�S���u�7^�>v8z��S��u   +��  �Bu}HU��1Z�FU�c�����h�8�:�*�(̦�1E�W1�j{=Q��37�k9���&7�����7S�k}nV�]S�������1X�^3ϧN1v�  X9w  �j9X�U�y��괣��Nc͕&i4Jw"�^��3'S�`�ԶX���u�u���Y����^�Kc��RUQ�L�b͕{�[7��gQ���h=�:  ��Rp  X��ۍrv*u�5Wǲ(�W��!�2O�Աa7K9�+��R�XS��g�s�\���Z���*���&)��rp9]�k$n�����r�R�1<3U��:  ��Rp  X��������l���:�
e�F)j�bK��^��h�:�:ƚ2���n���S'�{�r���ڝ�z�(f귢7�WL=�:��dln�u`oTe�:ƚ2�  `u�  V�n��Y[�7M�g*�N;u�5S�E�����:�-�G����1�TYÉ'�Y�
\u\��;�[9�n�$wW�����C�[�O�u�:�?z�7R�X3U���t����ӎr�L�k�n   ֛�;  �*�{g�j�R�X3�<�SK�:�?u�5S�1I���&�s��-�G���1Xgu�M����rgu+����ZG֪y�n'Z5*��FU,���:+&�sY�ZѲC"  ��(�  �B�nG��>��y����N�<�T�1\�LF���:���׽kW�}�x�����]�c�e����3�:Ś1���N��v�i�Z��ӵZ   w  �U�ˊ�u[��Sy�N�Y�V��pY��>��9{:�Χ��&��]U�:�׋bf2u�5ѽx!:gO��Au*��ϧ�@u��[���+�LE�i���&�a  ��Sp  X��&������[��:	S�"z��1V�$���\����S�c�����пb�eD���.t����.�Ι�ѽ4�:	�S�N��WUQ�Ǥ)�SK�:t u�5Q��   RK   `ؕӻ����l���>u<u��_��������M���Joq!zK��c�����{dg���ڿ'u��/����j�_�O�#�ȍ�;ѻ~=u�U+����o��u��gSG ��,c���V�nݞ:ʪTe���R� �+��1����c�Z]&�  ���  �J��Ř���:�����v��*K_���`UZ�E���1`�:�Ϻ&f�U�1�л��MV��|.���R�    ��           @��;           �Pp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          �w           ���          @�          Ȃ�;           YPp           
�           dA�          �,(�          ����  �����G����u�l�/_J�50��e���1�uk�(뢷�݅�(N�^Y��3P#����7�����D�8�uo܈���(NM%��{Gv���D��$�ҽ���g�u�l��m���߳�?�s�Jܘ�^ӟ���}���W>c;�ε��t�@t�]M      h w �����#�������`lyꙗ����q�˟��_��Qu����������x�����x2u�4�*����?�����1��k�������~�'��Wlغ-u��'�ƙ_�Ÿ�k_���Ig����C����O�Hl{Û#F��H�8y<�~�_ƙ�.zK����+���Ŷ7�mMfwa>�{�ۢ�0��?w����w�c���w�'F6l����ݸ���'?�����/aB      �i�z� @l|���_���������7ƫ������b���$d%6���x�o|%������r{D��Hly�x�S?o��ߌ7��ߍ���gR�Z��}_���~?�䧕�oc���W�//^���<�:κ�gG<�+�*��{��mozkv����M��"���S��7��-�s��۶����R���Ȇ��O����/�����o}I���������x×�]<���F�]      �����: @�m���xÿ����̳w���oyG��˿��?��X�MO�2��߈M��"u��l}��ⵟ����g?c�ݟ:Ί�x���?��{v��2���[�����ذm{�(5�yK<��_�����Q�e�cO������פ�2�v~�Gn*�gmd$^��;�G�����՟�'~�o>      @(� dcdÆx�!&zd�߳�'���� S�Z#6�3�������Q�v���P����}l}�����e���5�����x�(Ce�k^������1�U?��c�����ctӦ�Q���Ǟ����S�X����K��G����y������}P"      �)� d⡏}bEe��������>�D��?����ץ�1&���g�&���]��,�����h��z���5t�����3���>�:Ɗlz���~$u�������RGX��{v�c?�S+��'~��D���q"      ��Rp ��C��}����]�$��?���#�۶��>�����ק�rW#6ă���1���H<���N�b ��wF�������S���wŶ7�5u��z��Y�Ĝ-O�6�>��'      x��}� P'������X����w�a�Ҷ7�=u���a�=��g?����2�� u����-+?��l���[�~m��_�v~�/��pW�|�{W������5J w'�n    IDAT     pk
�  ����0������q%����������1�h��SGz�<�:�@�al�?XϿ͠=�����Ï��qG��7��#k�      ��� 2021��0:#��k�5Su:Quکc��>�=��mߒ:�m�:�Vmt|��L�LlLa�Fk�;�02>�����qG������7mZ�$       ���  �RUQ�=�:������O�NЗG��V]"      h2w  �k���#�{���c��K`��v�}��c       -w  �s_�|D��:������éS �e���Q�       ����  0@��ƹ_�B�CmǷ�7u��l~���?���1       ���;  ر��ݸ����:�����kSG ������       ���;  X�iǾ���q�����Z����/{y� }��[�Tly��R�       :c����x�x��{#"bd$q �����8��.�����?��q�;���۶��6p6o��^���l��M��Wk�*��ۉ����1Vedt46����1j�}�Bt��V�36=���<���G~�o��    0�^�����#��Ȉ�\�)�h||,���� Rh�=g~���/�B�(���} ^�O����126�*��/���oW��2���x�W���Q;���Oŕ���~ƻ&���ƍk���z裟���3ѹr9u    ��511cv��rn��+'bd��֍ض���-��?��5Fn,�`�#�:�����Η12WO� ����X  �1�iS<��O���RG    ~U�9y���׳������NK�������:���:��V?��KW��Y_
�w�������ڱ�"�?���{��
�@���;�������W�<�~�}��ܙ�>C �����3��Q�۩�     �*�������u�_��/��u������ߊ�W��e���O��>w,�;s��X4�h�     u5�����>�:      ��Pp��g������_w�̦i���	��TD�(���D�aɶ*�=��<��@��( 
"*2�(xPA�i��6M�u����~������|�$�����z�BKj��   PF-'��v      �aC�   �����^��[4      �V
�    e�r�#       
�    e6�E��i�       �x
�    e��fc�1'�      ��)�   ��G٦qi�       �h
�    C �86�zT�1       *��;   �i9�}��fӎ      P��   �����u3fń7��i       F��PB�|Tw����(�a�`��r���9|sO�  ʪ���b֙��LuMQ{Z�_ko��D�     �������=�;?�`U���j���M�}�le�t�/Ҏ� �]���p �
׻�=���Ƙ��C��3nϽc쮯�M�<X�d     �O��6��`��ܲ�ܲ�c0�U�    `�h���~�)%�      0�(�   ЦG���T���o?$j���       �Ȣ�   �@ۢ�E��T�Ĵ;�i       Fw   ������ik-z��cN����$      9�   (����G����y|Ly�a%H      0r(�   $���+"����=-�/��dJ�      `dPp   H��X��k��Ӱ��b����       �Ƞ�   0�/_�����%H      02(�   B��ƺ��,z��׽!��P�D       ß�;   � �X���%�L�����       � �i   ��'L���\�v��djjҎ �[�������1;�/jϔwK����_��D�       �'w  �T��F�O;P+��4���o����>���h����      ���    0����ѿnm�{�w��       �z
�    E�wwG�5W��v�����w�       ���   P�W]�����ls��K�      `�Rp   (R�����7��q�ݢ�U�)A"      ��I�   ��_zQI�����${       �#w   ��|����ޢ�L|��Q?kN	      ?
�   �P��ӎ T��E�ޑ�fc�1'�       ���  0��ץ�@ko�)z�-)z��#���ئ$      ^�  �{�������0�\.V\}Y�{��cc�{���@       Ì�;  � �7w���ݙv������uu�����fK�      `�Pp  �e��FD>�v���o������=u3gǄ7���       ���@����{5��=٪XݱnH�L�����hiڡ�� �A瓏��΍Y�D�Q�
ӶhaL?������h9aA����K�
    ����ksC��鮮�5�uz��1�)Ҏ��v�NT�#�ߐ��})�; uc�N  BU}C4�o4��5Q���:=�j����!��T�B	��ǲ�}3�cc�S�H;
)�����]_�;�<�f͉l�ب�4���ӏ=)&���E��T���g|$�V�GO[kl��S����"ױ����M���b�]�Ǆ�����>1v��cӣ�(     i:bBZ��J�:5�� �
��  )k�v^ls�b���l�ش�T�|>�=�i�xi�B,��Eǃ�9��\�Ϟ�v"���W�ӎ:!&xpT՗��n�������Ioy�?��B.���h��b��\.�d�Kۢ�E�#"�wJ����,A"      �ʧ�  )�6����tL?�������T�ޕ���[���XwǭѴ�kbܫ����S#S�M;VY�Nm�	�v�!5f�c�g��{�6�(C*��F��G����矍��L��ݝiǪx�+��z<��8��=����Xr��ѻ��D�       *��;  ��q����� �g�I;J����_Ҏ0`�\l����x�=iG���~��3�h9����LuM�iRհ�x����k����L�{zҎT�ڮ�a��ҹE����Ĵ�O���}�D�       *�g" `�5�_�|�����q��iG`��d�c��|'�~��������ޘ�uQ=~B�Q*��_\}kV�g�Q'DU}}	      T6w  B�{�6v��G�m�v�ac�]���Q,���߼(�rd�Q*R�+^;_~]T7�O;J����F�5W��f⤘���J�      ��)� ����m�x��QU[�v�a���gc����Ql�Ϝ�����cT�1;Ώ�.�"25^�)�?�,
}}E�i9aAD&S�D       �K�  ���^��6�K;ʰ����E
i�`����#b��'�cXhz�1瓟O;F��]��o�y�{�l�c4���$      �\
�  0�}b��e��c+]�<���&��R5�&��O)��J˱'G�+^�v���v��%��r��      �T
�  PfUuu1���cX)����~<
�}iGa��y�G��y|�1�������O���bu>�Hl����3��o��y;�       @eRp �2����Dͤ)i�V��svt<���c0JU7�����v�ai�k���*�`Ţ�$����N)~      @�Rp �2���Cӎ0������ӎ�(6��wGU}}�1����:<�k��7G���E�����J�      ��(� @U��Fӫ�N;ư�z�y��ٟI;�܄�ߔv�am�kH;B�*�r���ˊ�SU�ӎ<��@       H�  �h̎󣪶6�/��#���i��_�(Ҏ�(7v�=Ҏ0�5l�}T�kN;F�j����m�(z��cO�LuM	      Tw  (��9ۥ�����W?����Xs�/�NQ=�9j&NJ;���D��i��X�M������vZKLz�;J�      ��(� @�L��v��Ի�=�-����x��gD��iG�����49�#B�/آ�E?�����r��K�      ��T�   F������{�-�����Diғ���Mѽ���|�����ӎ�RU}C�;گ�2�7�/A��L=�����ن1%L3�t/y>��涘�Ʒ�g�.�G�+����+Q2      ��)� @9e���I�O<�}�%
lU&S�K/���?[�0���7��}�o�5m�]p��h9a��;      0��/�    Cl�~�O>V���o~[�͜]�D       �A�    +��A�;2�lL?����       Tw   �����[���=ӎ|od�6�       @��   R����/*zOvlSL9��$      H��;   @JV�������g�O�L6[�D       �Rp   HIߚձ��_��n�����%H      �.w   ��-ZX�=-',(�      �4)�   ����Gb�}�/zO�^��Ɨ�R�D       �Qp   H�W�      �J�    eko�%���P���oO�L�Z|       ��(�   �-��?���5����~�	%      �w   �
��ګ"ױ��=ӎ>1���J�      `�)�   T�\�Xy�O��S3qRL~ǡ%H      0��   *D��G!�+zOˉ�Ed2%H      0��   *DO��Xw�E���NѼ�~%H      0��   *Hۢ�%��r�i%�      0��   *��{��'-zτ���m_�D       CG�   ���L&�wj�{       ���;   @�Ys��ѷze�{��oQ=~B	      w   �
����/*zOU}CL=��$      
�    h�՗E����=-�=52�5%H      P~
�    �o��X}��E艹�����$      (?w   �
�v�E�B�{ZN:�i       �O�   �Bu=�dl�������e�hzūK�      ���   *؊EK���%�      PN
�    l흷F����3�-o��iӋ      PF
�    �,��W���5�lu�NUp      *��;   @�[y�Ց�ؘv      ��Sp   �p��M��ӎ      Pv
�    �@ۢ�Q��Ҏ      PV
�    �@��e��[Ҏ      PV
�    �Dۢ�iG       (+w   �ab�}�M�<�v      ��Qp   FV\uI�       �F�   `Y��룷�-�       e��   0������+ӎ      P
�    �L�՗E��;�       %��   0���]����c       �\u�  (��q~r��c�U��;�V����cl�緣���q{��]wk�1�.��=�Kc���5����]iG�_�����;&���Ѵ���z¤��\nSG�;�_rm���J�&=uӷ)j���_�$lI����Î��dҎ      P2
�  #��7�=�Cf�SΈ�5�b�y߈��,J;NYU�k��wK;���s��rȑ1������X}�ui'��ϝ/���Ѹ��iG)�ޕ�E�m)�>�:;ӎ0*t=�dl���y�ץ      �d��   �Q3iJl�ů��_??2�5iǡ�j&O��qA�������8�����F|�=""߽�$���v�m�Ҏ0j�-Z�v      ��Rp `X���c���ɤ����C�r�ii������N�[��ӎ2d��y2��Z��'��-I;ƨ��7����M;      @�(� 0�M9�Ș��CҎA���g�~�ܴc�j3���[Ҏ1�6���#k�)
}}i�=
�Xq�%i�       (w  F�Yg~"��A��&�sR�1F�L6S;:�Cn��קaX[{�MiGuV^wu�oX�v      ��Pp `D���]��a��cP80��֘�G��	i�r��}&6�sW�1��|��Xs��ӎ1��7w�ʟ]�v      ��Pp `�h��C�(����#���%��ZҎ����Q(�c�i��ѷvM�1F�W�0
���c       MK �#�4.��A��&���ӎ1:�e]���\������c�/�M;ưҷfu,��ܴclQ��B__���^��e���[Ҏ      P4w  F��իҎ@�o���޴c�J�+ۇ��b=�_�]�<�v��P��>���߸!�$[Էnmq�k*�ϙ���      �h
�  ��|t>�P�)(����M;¨�����_d!xK6�{O�v�B��3����_ڮ���ΰx=���'=[�劚
�cl�g!      0�)� 0"l���ѻ��_�fpV����#�Z�\.V���2���7��,�K�{�s����D~sW�Q*V��/�%��Z�1d]%����>�֮)a��X��+�      ��� ���ǒo��v
ʠ��Gb�M?O;ƨ���߉��+K���ǋ�{�s%�[��x����o�괣T�B�?^����/|*�PH;΀lz��X���X��o�>P���ѻrE�1       M� �aoɷ���?��X����GN���ӎ2���_O}��wo.�Ύ�����Œ�
��������ӎRzW��'N=:�.�8�(�=��O$�b�օ�Gǟ�X�D�U����/O;      ��)� 0lr�X��/G���ӎB������'1l^��:�s<z�;J����[�S��|OO	���m���G�3;=6?�l�qR������N<x�~ö����O,8&zۖ����.�%��J�S�֊_���c       Ju�   �B!6��w���_�����vJ���-گ�2�.�(r]�i��t>�X<���c�����M��#255�-����?�+-����R�eV(�����7�"���/&��h�{���9;�deӿqCt�����n�5�����iG*Z�c�C�3��hL;�QUW��3��}&�|�˱�nN!aq�׭��7\S�86�(       �e��qZ!�  �]�qlL?�ĴcT�\Wg��\�}�W�g@�f̊�9ۦ��e2Uѳ�56?�������㚷����6��ޕm#�5�lӸ��1+���Gd�i�)�ܦ��m_��miG)���1���}�n���64Dߚձ�ч���'ҎV��Ysb�A�,��M�<���      �w           *BU�            B�          �
��          @EPp          �"(�          P�          �
�           Tw           *��;           A�          ����          @EPp          �"(�          P�          �
�           Tw           *��;           A�          ����          @E�N;�?��u3gGu���j��͑��=�[�oͪ���������]���!�����}&�H�U��c^��Ȏ=˖F�_�J5O��y�mlL5�P�Y�,�׭M��l������z\s*��:c�]w�r7        @)d�k�a�vQ=~|d�6E!��ܦ��[�6z���\.�C"����]v��IS����|�����+�LuM4�k�L���G��G��'�<5'Emˌ��OCnӦ�^�\�1���*�v{U4�kd�k�{���wG��;�d!Ղ{��&��}]L>��1n�}�n��<۷zet<p_���W���[#��9�I�Fͤ�1�S_��o?$2���K����b�W>���7����1�߿<82������gㅯ}1��yk*��}���>�ܝ�g?��Xy�UC~ovlS�����Ï�LM͐��7݋����7��        c��;Ƥ������N/���o��'����kn�e��.�C �����3��᨞0��?����/�(Z�^r�)ܺL�:�y�c��O��cs]��b��Xz��Q���\�zglZ�ɦ    IDAT�����i�p�]���G�#���+�}�Ѱ������֬����X}�u)%��{v�V�K�٘���b�>���$��߰>����h�⇑��U��C��eF�_�������s_�t�_}ِ�J�a���Η�4j&O��
�x�+���E�6XD�|��
�C��y|��g1f��Cz�ҽ��x�
�        ��и�n1����c��|>V�x},=���y��XUU��Wϋ)�:�%���ݝ���ǧR�LuM���˷�k���O.8f�_s�~̉
�)�x���o]�����X���0U��k[�����4���y�*�G��D;������7Ѵ�%N8�2����{�o��GUUl���cܞ{]�255�����t�=""������h��uC�!��׾[�v        ��"���Y�x�z�̓+�GDTU��w����h9�}�LiC�`��?��r{D����s?���	4�?��/Xh��1�?�k�����sc�s���r{DĜ�}f�wm���޸�n������%��c����.ɾ�L9�h|�.[=��fc�G>=�����#�~���؏����1�7�        `بj/��c�?�l��}uu1��_�yg+�j��@.����bƂ�촣O����˜(��	c�{O�٩G���7����̨�o���L&f�����`C�٫q��b���F��	%�[U[/���1�o)�ޡ4��o�٦W�5�&�1��$)6���Q;eZӐ���W        �BU����?���+�������%���������'�`�%7~��GU]݀�f�Y̎��Ӧ��(y�z8��{u����F�����T���^�m_����n2���ffٲV݌Y?��Dݬ9�C*j���        `���s_�q�޻l��zTL?���/�����
|�=Q�2vIv255Q3iJ��LԵ�(_�
7$��v~�Q�ʎi�ι�$ߢc�U��':���W����d�@����#��+�         �C����U�{�~�1f��e��Ԓv3��eJ2xU	��I?f�������Q�_���'xp�'���8טz�1Cr��:{8�         /;�)�|�3CrW��&�~�KCr@��������9��|9�x�Yg}2�c��N b��D��5i�         �h3��H�L�:d�5��ژp����>�b���>�=GF����Ej&M�iG�0�w��M����#�PH;
        @E��4%�sҐ�;��OFd2C~/�`�����fcƩ(��-���ӣ��!��a4[s�/�/�qV�:ӎ        Pq�9%�~c��]c���8���C��1����\}C���?�.?�e���'�f�T�T�k��w�s��l��'zۗG�䩑Әx�fҔ�v���v��u?�7wE��o��jk����|>�7u$�T=�)����t�$V���X�1�����{Fͤ)��f�ޛml����J�        `��L�ӏ>qp��|���EUMM�L�:�3��h���탻�Q������D3����un�B.7��Uu�QUW��^l�o�ν0��c��c���Fӫ^ӏ;%���ɱ��{�4SY
�lu�|�Y���==���_��k��B__d�٘��Cc��5q�}�SΈ��/�|OO����?�~����z��1��o�|O[k���=ez�m��Ysͤ�o��h���%�ټ�~1�����         T���Ucϭ��X|�Go{[DD4�|����ߌƝwK��i�=�y��c�=�M���}g<y��>_�0&�z�Dw<~���|~�G?3����ٸ=��Ͽ$2�5��竛���/�*=������C��,�AO~�{���^(�S:)V\ui����B.�~qm<}橉3�N�S?6�         @)U��ӏ=)��ʟ�8����^n���|��x��#��ui�}�>���3�Ȕ�fc��:�%��SU�;|���d�������3�l�x��ϭ��'���;��ϭ�ݝ����q����6�         @�ls�i�m�h�wU{����F
/����b�9_J��i���y��&�F��}^���نy;ĸW�U�D�O��~��?ؿ)��Ų��♥��zD>�hom�61�=G%�         (�lӸ�vL��ۗ����m�xɟ_s�������8�#�g��g쮯Hv~�=ʔ��J[p������xl���l�[et��Xs�M�w�x�Y�������|�ޞd�{�˔d�
�������)	         �͉�E���D3}kVE�O���B!�]���y���oH_b�2�{��*��
I{�I{�#]��K�&�)ɋ���>�wƘvJ4S������~#�+�u-3bʻO4���Ӻ,��˔d�z�Z�z        ���6����=5���K.�|�歞[��_yŝA�Y��WٳlI��^ϊ�	��U��L&��Hv��+�g21�����O�{�s:����b��7'�c�igE&[�x��c�on�ٞ�ˢ���ʘfp�|�������ʘ        ��i9�}�_I�_�.��h`��Xvѷ�����U�I<���q��ѿqÀϯ���2���w����_e_��eLC)���>�-o�1;�O4S������,=/�+������w�h��e�on�M?0��K�=;�ﱡ�~͕�Ӻt@g[�_��        `�Ȏi���NI<���#׹i�����W�������3����h��;:���[���ʜ(��m�~��:���#Y��_+M�=��'��7^��6�L�3O�7��3>�l6�#D>O�}ѽt���^��X}��C*�|��x��o�-�[{�M���Q*         ����=5�'LL4ӿa}���d��������ф����"�#���.��7\��3��=���YC�(��_�bl��-��]�"�>�Ԋ|���$��o:(w�-�P>��?���}��B�����Ƥ��5��z�/�Gk����uu���m~��x��Sc�7�N)��t=�x<r�A��_��߁ܦ�X��/��~_r��        P�0&ZNX�x������7�o�et=�d��Unq�!���3��`<�ُEϲ%��S�7D��ߍG�}w�oܐR��������e��nh
���_�#�����,եX2�Opkn�aP�L#":�x4���������<㣱��_�
�Q���x�K���_�B�o�}T75EO���i]�v��i]O�qB�Nk����2���Eϊ�������N;        ���r��Q3qR��\��Xq�wa>�}'v8��Dc�tP4��5:dp�2�
��ګb�WE��m�v���߸16?�Lr�i��B_,=��h������D��������?zW�H;�Pt�}�ޒ�[T
�l��-��ܘ�ƷFd2�i��CLz��bͯU������z��c���-��֖v         �AUØh9�����-,���7�"f�����N�dbƂ3���o��2rt/y>��<�v�A�wo���6��@U�f����3kn���rq��ĺ;oM<7�C���*��         x��G�5�&'��uuF�`_o��|>Z/�n�Io}G�y�ˋ����jz��c�n�L6T(D���+�ڿ[z�9�B��1�����         �7Uuu�r��s+��A��[[��kn�yl~�/Ɇ2��qڙE�P*E�g��Ég�����|��b������u����s3?�L�$          ""�uB�N��h&��+�.��$�r�h��ۉ�&��h�v^I2 k���= �^���s��Ĺ%K��z�W����SIs          �WU]]ls���V���[��d9V�x}l~��D3�l6f�vV�2 c���'�}�oo�M�<8�+�����~{⹙���9         ��k��E�D3���h���%�Q�����I<7���E���J�`0Upo��u1��{'��'́X��䯸���U1���%         0zdjj�z{�՗E����Y}�u�{��},y��Up�yF������o���{s�Vu>�p�����s3?��2�         F���u��L4����^T�<�}�}�!GD���eH0p��M�zM��s���^���3I,��W����WG�^�-S"         `��T�ČS?�xn�WFo{[��������^]�w u����d�K6��w��OL<�D�c����M��x�          "b�GE݌Y�f
}}���˔��������&��z�щ_�(�D��W�:���/�%˾���3����$�i��1nϽː         �2�51c��ϭ��Gѳ|Y��U��6�?�h&S]ۜrF�l]����3?�����ޓxn0:��^q�y�GJ         Ѧ���9;�L��/ZpA�����+�G��Zʐ`�\po�}�h�w��,ī��Xv���g���?�vߣi         ��(��ƌ��J<����Fϲ%eH����ѽtq���������)�����2�OT�96����s��x��p�]����         �ӄ7���&�)�rѺ���z�;�������M=���6�+C"�-P��v���x�A��/� �kꥰ���H<3��o���ʐ         iZ�{J�տ�it/~�i�l���$~5>�86�zT���ܧqld�k-���C���;�X�~w��L6ӎ<�L�         ���a�y1n�}�r�X���/���`_q�~�IeH�e*�O|�[/^��o&�)���}=����V�$         �H2�o��dͬ�����³eJ�u+��į����6��8�L� ����k&M�Ɨ�h������uСJ���b���h�a�Q?{ny         #��׽!���K.,C��+����K/J<7�7�!�K�j��y��"����ߵ_{eD�0�P��v���3��C         �jk�i���lz���|��2%�U��$�7nH4�W	��6���1��B!������)�uwޚ�q�N�^�         F��9�EUmm���7^_�4��:c��ܜh�q��#2�2%x����l��D;�|,zW�t�R*������L4��ʔ         ���xf�]��!�଻�׉�g�6E]ˌ2�x�����l�h��4�0�����3/Y�         =���Kt�������eJ�ܦ���*#"t+�!�Ղ{���v=��ÔC�<ٱM���)S         `8�7.����+�Wٻ�=�7�O4S3ab�� ��V�ٱc-�]�j�aʡo���3���2$         ���ئD��V��)��%�VV5&�c����1��:�r���$��         �	{���1�[nSG���	K(�V�\.��Lm�ÔC�?H""
}}eH         wýWQ5&���z���j�=�W�4�t�r��<Oҏ         �{�2"�f��D��*�����{�o�Q?g�A�)��y;&:_��"���Li         ��,i��a�veJ28�㚣f��D3���eJ�b�[;зrE�Ϛ3���;�\T�Rk��k��=�K#
�2���������woN9	        P	zW�':_7knd�4F���L��i�e��3=�Kːؒ�m��B���L���|���Q;eZ��J�9p0�Zp�z��h�c�/��}#SS������D&^��D#]O?Q�0�pQ=�9�9�1���E]ˌ���]����h����߸!�        @Z6?�L��l6��y]����2%J&i�2���z6��o����v�2�#c�!GF�����ʟ��l��Wm�@�O��ƱѼ�����v{U�NoI4��̓eJ�s�Ů��3���r{DD�����ػ��8�;}���Vm�jW]V��;űF��� &r	�B5%$p��K��H �z1�1	�H 	%@B�p	�YV/+i{ߙ�F˻�5��ή��_/�l����E��>���~y=�<��s�ULHDDDDDDDDDDDDDDDDDj��ܮx�����d
DQq�hw'�H8O����[����1��?������,���]�V}�KS
�kS����^�Q)И-X���`lh<�9ƆF,x�����LFDDDDDDDDDDDDDDDDD�"><��@��5��-�Α��x��(Z�^%e���g�p����؇.���}$�>EZ~�)06�L9T.��U�8�ӊ֤BA���<%"�bWs�哚�n�ӄ�/�/@""""""""""""""""""*Fc����Ec�>Q��L^�E�+^3��o󐄈f��K����!�{Ȃ��J��Λ�T�hP�W��)'j/��Ѩh���7!��yJDD��u�9�?���򘄈������������������Wa� j/��9i&�zħ�8�xEk�X�?�!?����	Z�'������ �/?���]g�CYs��u��wW��_T�n��_�!�A��y�;Oj�!������������������������7��)Z�-w���/�S�Ck��&�kF~�R�P��Lall��cj's�؛�E���9M�~`A�A��c�ׯ�j�)���:��ۣ]�1���󔈈����C�L�Kb��d���)�˫�(Ⲭv��c*3A6&�	"���R����O��>�X��	��� R��J��(״�*hk��D��	�:A��f�V� d���{�I�I~�""�-�h�O�u�_�h]�Wc`��B�<%��z�r�W�V�n`�cyHCD3����1'��$lzM��=E�:�<���{:��mJ��ը��?+^7�� I�C"""""""""""""*&wH�}��]m��h�pL��A�ө�(:z�06�l�"�O|���Z���ٳ�pX�DD�s�8�W�1hi��wYYN��7r�lʴZ-a�M`�����*%"""5�|j/��v�ϛ��rT��>tO�ej�V�����6#���yHCD3I��9Lq�'>�3$F<�\�hQ�W����+��hPv�nrlC�<��DDDDDDDDDDDDDDTLDq�o�Rh4��c��Q����c9�4�����}~���j/��%���;�����}��<�!��$��a��Ws���~�F��ѷ�~�p��eͭ��M��]��u*^���O�
�򐈈�������������M�B5�'�.,�Q���u�|t;��Tw""��z�r*�h���Bi����	}�co�>i�h&���o#����q�&شa
S�5���zEk���ʯ@4�Iz�0��'򔈈��������������Ņ܉�ɲ�1�]S^ӑ�UJDDDj�v�)�)�֣V�~t��u���Ȳc	 ȩ���]=���<����	���_�S���ը\w��u}�ދT(��DDDDDDDDDDDDDDT�DQ�ۤ�GZ�6���DT
�/�����THBDDj+�)�S����o󐆈J��!��C���{�)��pޮ�U���g����+��pMz����_�N��&����Mox���"""""""""""""��d0Ԏ@��X2'V�R)܉�$H��q����x��}��Z�]���,��~NѺ�K����y�k]����*^�s���N�c�H�W�v�	���墨��I�?��t���ٗ₻	���b�W�S�:������݈�ޥ�������{݅���=v?���2,��ݞq,�����H9Y�!�2AHӺ�`\�ѭ[TLFDDj��N�֮���|-s|�{�C��%Ӝ�Lo��}��<�!��dI�O�HE��[q� �7>����(�)��W\Q�W�&��b`�c9�BDDDDDD��$p]��xB�(DDEA���F�2�z-��48� �4 �!����J�Q��Д?�
��x\�$DDS�� ,'�Ƃ;�,�����>糊��k��}屰�X�x]�}wpz;�nJ�b��n��������� ���B%�kz�����DD�����1|`�    IDAT�P$�����Z-�&�XoP�aݝ���J�(����,R�͖q�܉��H�Q'3w<�ަR"""RS�}w�u�yE1Ž���	�����MNsM�x�S����(�#�֌Oqϥ����|z�߇�'7�4?�ۉ��K&������0>����<���=DDDT�8Ž8d+�'�q��J��e­����y*�!""��OqW��ҫ�1[r��~t;lˏQ����?$)g9���j�w)F��*^�:{ʚ[�z�	5u�<����?� �~_N2Qiؚ�����ND4�$a���=�8y���KH�����h�,�ܕGhj�Z-G��p8�B"����-'��B""*=��9����)�R�~j��G~�J�2M����Ȣ�#���
��^3>�}�ׯ�Υ uW� A�S�&�c�g�N��DDDDDDT:�Mn��l�+���h��e�$!�L"�#�g�@��H4����x{̈�+��bY����jU;¬WUUQ�8�-�"�J����hj$I��zf^u<F��J���HM�S���|VѺ�K����H��Ӻ����`[~��u=?���ۉ�hL��.E����C�sÿ+Z�:{z��ݻ�|mCm=*����u}?}��ۉ�����f�l�v�ۍ9s樘����ɲ�X,�p8�@ �@ ��v��D���+�v�Ra@�V(pZ"""��1��E1��]*����c�PH�$DDӓ�&qC�<�����V!���;�:�<��W4ǧ��>tϴ�]�����܎���{Z�%"�%�Ч���G�Q�f|��t�Ouz�O�DDDDDDT:Xn'"�A`4�t:��؈ŋc��Ũ����`Ⱥ���å]cx4r���DDDD�BX,�c�jUUU���
I���/�)A���5�!""�E�v�������jh�S�b_�zJ�ۻﻝ�ۉ��L���
���Ӈ�s��eͭS����^�� ���Ü�NDDDDD4K��ND�[����X�x1���`��2�I$x�{��&�T!#�R��OC�a4�p8&�$�w"*Y٦���;Q�$DDT,z�rJ�+��Sܧ������ځ�߼4�k�����8������ˡsVLz����_�N����M���` ���NDDDDD4+��N�DQ��d �t���i���v��"f�9}~*�B4M�<
�ߜ�F��BH$��OT��V+�V+B�������c��,����Q��aS�	f�݉���x9�N���f-%R~555A'�c�����J�$I�h4�[me5�C*�"""5E�v����ý�|E�j/��6 
*Z�8�x�>�|z{�}wpz;���S���xs��uE�\g�C�w#�{פ�j������ ��*^GDDDDDD�ek���7���r�Xn�t:�n7G�\k��'|o����Z�e�\H$�B�o�p�`�Pccc�z��x<��|���C2�Y�43��f̝;>���݈��w�����~ZcAe��*�N���j���W;ʬ��Ғq��DT�$I��z�(�r©�>��z���HU=��י�@�L��9>Ž��{]k*�ۣ{:0��#"ʷ��`���Q{��Ж;'�f*S�믹Q���O
�DDDDDD4�qr{i�j�p�\���Beee����jTUU���� �:���c�k�^/�^/�����ߏ��������CCCH�RyLL��7����app0}��K}��uf؊��/Q6N������lp:'���J�*�PIDTl��b9�D܉�f�螎�Lqw�� 법��u��v�|����P�
��%���M�:%S܍s�������ArlT�Q������o[�(�� )N�#""""�����ҡ��0g�455�����ͨ��CEEE�'�˲���^������rY�3���}�w���.�� �F3���������%�I���}}}سgv�ލ��.D�Q��"R�(������fCgg'� �
��"��1���;���rtww���jmm�8����C��J�$I�h4���́�߫R*""R[!���_�Ź�]�1�������W���X �^��|��J���6��7>������>�	fJ���_�UE_�@����Ӈ�)�T4��|}M]��L���A�R�&�)�F��^�*++'�QWW��F�dH��D"�d2�T*�d29�ǩTj�����o�]��@��N��V��^��F��^��V�=��y�V������`ٲe>߁��޽�w�Fgg':;;'L�&*F6�����Ν;��}�k$��:~�6������(�(�p:�V;ʬ �bւ��ؘ
i��rO��	�	-,'�
�O�������Ӂ�W^���u��Mv���N�����{�(�B�	+:�Pd�J@y&�*��!��T0�����w�&��>Oq����"1:�x]!%�X�<i��/�'>�c��h4*Z��)�6��^<��ڰp�B̟?��χ�b��zY��H$�ŐH$�����?��6Y����-����h4B��e-������Z�����c�M�z�ؾ};�n݊m۶a�Ν��NEG��c���صk�~? `Ϩ�3��-knwj """ʅ��jx<N/���6�{o���#�����(��Mq��>�w"�Y��'���s ( 4�)��oT�'��	�˿R����>e�J��c��ّ���HQ��}�jEkO�����܁�Mq�����QC����GO�|�ɧ�z�
��/yL59�N�9_���5R4���@��l����r:�X�p!,X����eR��%IB,C4E4E$I��g��i�ي� @���`0�K�eee0���"�����+�b�
 @*�Bgg'�mۆm۶a˖-)��iv������o�
��j�����JD*�z��-P;FI��R�>��
��Q��v�	�a���~N*)1;
�Gڽ����Agg��1f-�^����K�(��?~�q���L���^vħ �̐9���h֊���ȯ_��,eC~5Ž|�I�~��<=���v �v�Qt�h,C�57���o�)�25�^]�Kњ螎<�!*=9/������!4\���ֹ�^���Dhۇ�~���9 ``�$F�����G[��>?������G�C�cg��*�V��7�󢥊���(�����������^xN�Gu�.]������k��x��>^h��㜊�Y���������e�������`�F���V�����3� ����o����[�lA0x��K��EE���`ǎ�H�R��� �m����I"�9��
5?y\�%m�֭���x�E�U���G.K�t*;Ք�_� �'�|7ި|��NMMFGG�|%�Z[[3v�
�ܕ��fY�'��'��������S�ں��Z�����?�5�c�^�97}Kq�hW'</=�x]���� �@�]p��_Fd�v>�1���b��h��&�����<�!*Myy)=��f��A�A�]a�U_Bd���q��8��G}Q�No��p��5j��及���UX������[1�̓H�._A���h�雰�)��}｝�PDDDDD4�lM���&��].��9��h�`�,[�˖-CSSӄ7��'I��0B���0��0R�T�<������ ��ja2�PVV���ɔ1齮�uuu8묳 Iv�܉>� |�>��=-���(��;w.�oߎp8�`8����p�]��}DDDD�f08�=�DQĢE�2�{<�?���H�lS�-�Ob���h�����ˮEt�n�����7 �ق��������}�� ��aD:v��u��	Z��#X�Z��{oG�[����WV���P}�%��� ��1�ÃyJFTz�RpO���A�S܍M�8��? ������Odَ�P~�Ӓ�� ��[ٽeͭ��i,V4���1��o"��c$�cyJ��� Ü&�݇��w #�<��DT�̋�½�|������7���rE��k����&�@�(����H=�ܞ_��/Ɗ+�b�
�����H$҅�P(�h4��CQ��h��j��j�? A&�x����h2J��,O(�˲���J��J� I��d�ǩT�`�{2������O>F�&�	&�	�:�.}�(�hkkC[[>�� ��>��͛��{����$7�n�;lݺ�d�.���Q��������ͺy�x����^��HD�DDD���u��e+���"�Y���;Oqt:̽��]q=B[�@�`[y����b=]~����2��K�����׹��,��|��]�B���u���
e-s��C���9ET��p���ˡ�;�4�V��ֵ�X��=0��(���~�9_�Ɣ֊z=���8Q~�7�i~�Y����/T}����E��EKU�@DDDD�������Ԅ��v�\�MMM</�H  "
d
� �j�0��t�����x�]��@��dL1/��{<G2�D"���>�H�(#�2"�"�HzҤ^���j��b��l�V����C��+��~�!�����3r��h_z�MMMعs'����M��
ݡ�N�Cmm-���Վ2�X,����T
CCC*%""ʯ�a	�VMfX�=�7�b2""R[d����E��<W�ڲ��{�����]���s����O�����/cS+�M��AN$0���ՎATT�VpO��a4\{S�.q@�On(��~�j/�vJwU�����T;��ܛ���uj� """����s������8����А�Y�
�����F�e��������E���?a�X��Q'LO�&�L"�#�#�!������x<����tὬ�V�f�f�9}3�F��ҥK�t�R|��_Fgg'�}�]���[����I�}��vTVVbhh�^춻Ь-���DDD4{��n��� �e�X�|yzW�qCCC��OD3�$I_�,ǟʂ;��;�:��@����{1��/z��vub�7/�u�9jGɫ��F��O�DE%ow��)�_�L��鐢�>z_���+��=�݁��W�(y3��_���?���|�I,�QްܞUUUX�r%��۱`����Oi����B9-� �ј��P��f|��d��X2�D4��&IҴ�9>��[ķZ���l�Z���755���	_����Յw�y���:Kk� ���:x�^��q|ߟ�cμ�DIDDD�� �3g>��cȲ�v����؈���	���0�^�J���
#ۿ!�������KDD�ٵ�W����
z����\��ys�����I�A4��%/R� �����1��N^�=J����h���y�	��	Oine7��Q��<�%G�%��1����T;�Q��������f��I��^߄r���b�}�\.�?�xw�qhii�zN4���������Ev��P2��բ�ja�X`�X&���D"�F�����S��@�$�|>�|>� �������^�>oΜ9������~�!�z�-�������DQDCCv�څ�c>Ĝ.���ٌ��Z������Y,�X�b±T*��>N&$��O�eȲ<��0�jE�����*&#"�b����y��e��p�!�k���EA��k��t��64��M���E����Ѐ�1��N��#>�����zħ�})���W����ɩ$��p9�>�[hmv��䌜Ja�]�-4f8���jG """���ۧFE,Y�k֬�1���2��������z���w�L&�f3�f3ô��A��C���n����X�P(]x���	�,#
!
������#�{8��iɒ%���+��{��7��_���iO�����p�f����������y������W��(�hoo�x~��ߏD	N�$"���� `9�T܉��~t��V4��w
r��~r*Y�k�C�c�þ�X8�;Q�(95���0���ՎAT��^p�S)l��_���W����߅$	;��z�¡�]� b=]�x�EX��SgH`�����~�v���N�+��,��թ��$��JDDD�W�ܮ�����իq�Yg��re|<�������MkR�����B��d�V���h?��N���)��p�P�`�H$�V���088���A������:���|Z����hoo����|�M���+*���H]������x3�W�3skY"""*}����裏XȞ�#�<2������J���
O�$��8�e�?aH ����������.=
����u6m�����z���$l��
,z�9�.Q;MN��{߾I��%)ߍXNμne1S��-��� �>Ǉ���a��OAkw��]w������.4������A�]C4��{���|�Q;I�%�����S�D{����U;F�$�>���BDDD�/[��zNn��N���>��v�.]�1*�H`ll^�wZ�v����
��
�ɔ���O�Ѥ������{ P<�?� ����f��v�=}3CEE֭[�s�9��>^}�UNu'E�f3�V+<� BU&���ODDD�G�բ��;v���uhllĂ&�BV)�:dYΘ�)�@ّ�B�6�������,c�� ]����r�����=�~'/�]h�` [/�<�s��/R;δ���>��RH��Q�J�Ő�����}�'�v1iz�C����S�L�����E�0��M9���������Or��j{�w���Ϡ�G�wW�G1)��o|���S;JA��R4
�h�������s��{�5ؖ�v����;�#�X,�ONUU�:�,�x≰�l>&�2�~?FGG�<O���l6�f��j��'xS��h4��l�?�D�`~��`)���B!�B!����f���t����+V���+044�W^y���o
��.{T���رc��M�e"""���X,hii��]��4UVVbժ��X,�����Ѭ�� ,ǟƂ; R��^����ʏ?%����}l��BH
���g~�\��� �'�gJ��ߺqƗ����{��5�s#�v(.\��x����O�$x�~3oY�����;��X�3��矆�m����~<)Ş[���Vn���gP�:eM�jǙ�ж����O3c��dȉ�V�G-?乩�;��H�H�Nx�V���,4f��Q�N�Ǳ㦫�U;
ь�5	\��Pnw�\hllT1Uqimm�%�\�k��.��`H,���񠻻����+|aL�ף��UUU���Cyy9��ʠ�hr�i�
4����p8�v��7.$�IEe�X,�׋��Q�R)����ٌ#�8����QWW���^�|�|}J4��� ��bmw� *6��ۺԎQ�<OzⳐJ�d�bE�E�p�3''T�g˖-x��T�Po1#Vf�pL���9��j�����zՎRԜN'N:���O���]]]��w{w�(//�pL���J�̶�n�ڊ
x�ڨR""*6r2	�?����1�A��l��_b�W 
� aq��1x^��X�#W@�l��~������
y=?��v�j݅�~7�e��� ��GHE㒣#0�e��y����`��'�j��܁���=/?���]�,Z�h�<���W_����~���ED���y�W}�e�mл*Վt@��At��Ct|�F$�ՎSp��߃}�*j�x��Jb�W ���
��0�D���kΆ�7zA��SI�������jG!"""�q4�����o�-_�W]u.��b477���e>�}}}���C(RTJ*++���B}}=���`�Za02�J��"�z=,\.l6t:$IB2���cH��P(���D"���^A��h��܌3�8�-B0D___�?+*U�d���٦W;
���c���`����L&�0坲f:�łSN9eةT
]]]H$*&#�R5�
���[*����Hz�TJDDD�(���`������eM-Sz��Ώ������=�g���e�����W����BY�<bqQ��	?��_�/�o���q
.>8 )����=o�WO��������{�m8OZ]���>ڂ�_�r�p;��>�`    IDAT.�c~�8��>�h4�PSw�;i��{0��M����b��H�fτ���]|j#��@�����f�� E���6z�߾�|���o9���硵�a^�8�N�h�.l��2��U��C���a���AYs+�����몔��}�_�
co�V�(DDDD3΁��s��Q1���z=N=�T�x�8묳P]]��X<������166�hZ��hDEEPYY	�����,���`�XPQQ���rh4�R�I��ǧ����A�e��AP]]�իWcժU�����,�y�����t:��2���~Xp�>�I	�K��j�V����W;JQq88��QV����%�Ituu)�]��h�L*���1PB
��G�Q�J�z�y�9���*�D��zhL惮I���������B�cG�Ҫ/��b����y�9��>h��9]j�dyoGv����0��3H�Cj�RM�o�������H�?�{~�=���B�F�y�Y��+`:l���E�DOn����C*�aᏇUşA���m>L��Ck�C,3AN&�
���F�����x�Z����}]=�V]a�\�>ć��؉��-���T��
�cW�P� )Fh��7�95�b�L����y�"���sZ���܅H�N���H[��5�>D���1��5�'���v�y�8��3a�M,AE"x<x�^E%a�^�Á���	��&����)��B8��n��	����/�K����.��̷e��bN9�ٝ#**���ozQ�%m�֭��B<���:��gԃ�#��*�2�}VѓO>�o�Q�GW��+�X��t��t*%*^###سgo�PYY�իWOx���������D4-�--�ז������J��Nh�����D�g�����J����EK��pCk���d ��w�m!ڵ��i�
���8�Z�b�	K���QD�t"�u��Y��G����0�F#�{:�}��Y5��i�X�\m��Q�����:7�M��������fNn��b�����9��i�m~�����&g�N�Cyy9GFɘH�p8��ҞJ�&��j���r�j�N8><<�����*b�|��i��ݸĦ�:�CTTXp�>�I	�K���CGGǬ����������D"tww+z�@D��L*�����/���,��KDDDD4Y�C�BDDDDDD�{,����l�ڵk3��$all��Ê�g[�V8�N�l�������d2�d2���~������\`0PYY	��A�v�q�e��������?�W^y�}vr���j�b ��"""*-v�mmm���P��m�X�x1�.]
q���}>fu韈�@$I��5 ,'��Q܉����2��NDDDDDD�5	\��Pnw�\���n4q�g���χ�bIO&����Ȥ'h�t:8�N8�NNW��E���x���KO�=�X,���n����������Kp�y��W��^|��C>�<&�	~ o�!""��b6��p�B�ٳcccj�)�^�c�9�c�$app^/��'":����0��OTJDDDDDT�Xp'"""""��ږ�[n��3���r���Q�T����p�I'��/Dyyy�x2������Դ;A��ڭV+��S���zTWW���
�@ ###]����Ӄ��A��n8�N���ݎ�/�g�q~��_��^���Y�h4"���;�"�F���x<tuuA�e�#���B{{����c�z{{��&v""ʔ��Ck�u�H����������x��NDDDDDD�5	���"�Ǜ�n�{�Ln�j�8����}nB�=�J���Tꐏ��hPQQ���
Nk�� l6l6��(<�^�A�D}}}�����(��������q�g`�ƍؼys?R�(��h� xS�.���ٌ��.�A���V�őG�y�楧K����Q�����T"�Iʘ�.���cQ/Qb��������
b��ۏ:�(|��_������`xxxR�v�^�Ӊ��
h4�|�%�2�ш��z���`ll���H$<?�Lb`` �gBѽ����ַ��bÆ����Y�,: N�$""��VVV��;###���=���KECC�/_�ɔ>
�000�x<�b2"�ғm����D܉�����Â;�ݶpM�oB���r͊r{mm-���/���=}l����x�L&�&�	n�6�� �3.Q�h4�\.TTT������ ������(���һ,Z�?�я��������p�>*0ݾ숈��J\EE�����xJr¹��G������X,���߯b2"��%IR��
��Eк�Hz���8܉�����(�����=>D���1�˅��FS��l�g>��]�:���	M###��h=�f���v�l6�;.Q�� ���Á`0���!�������ݍ��aTWW�o�hoo��������g���0i"܉��h��h4hhh@MM���0444�ݻ��r��hѢ	;��b1������g�>LDD�'I�}�,'����*�"""""*.,�Q�lM�{�&����=�]E���K�p8���~?������zo�����������KTP���P������F���	�ٌ��j��f\x�8��S�q�F����LO��ӈ@�6%""":$�V���ZTVVbhh���n�EuuuX�`*++��C�FGGz�*)��F!s��,��w""""""ʋm)��^߄r������%K����/GSSS�X,C���o����a��f<���ٌh4���ax��N��Bصkl6������r�p�7��O�C=������������l��^[[�`0�������:ս�����hii��d��yl ���C<W-�L%I4̈́ce�	�́�߫R*""""��;�ܶ��ǇH4�>�r���بb��1�͸��q�i�A�V4S�122r������`0
��h�F444��vcpp>�����~�A��n��n����?w�}7^x�lڴ��`���F�z����k��Z-�nw�ho��!�2"�<�� "�H^3��)��#����|��������������DDDDDD�S��ܾb�
\}�ը��HC?���A��l6TUU���,�1����hDcc#��0��'I1::���j���C��bݺuX�j��>���/pz""""��EN�N� �����
��F�F���`�m��`��Q^^���JTTT �L"�#�����H�$���""�C�6�ݲ�$܉����>��;��l*�;�N\q�X�jU�X0D__��|�ٰ�N���dBss3� 892�H���ccc�����hDMM�����w��<p�i�DDDDD�J����r��r���R)D�Q��q�R)H��� t:�Z-�z=�Z-t:�Vkz����� FGG���_�����Lf��J��������DDDDDD����.֬Y��.�f� �L&��ߏ�����5�L�����d*DT��e�Za�Z���000�X,���`0�;v���n��(���K�,���>�7�x��ɉ����rO���l6���NF8F8�c*""�.Y�!B��� �q' ���*�"""""*,�Ѵ͖r{MM֯_��?<}��󡯯�D��t:���Q^^^��D3��n��f���(�L&3Αe���C}}=,�v;��կb��ո�{022�Bz"""""""��6�ݲ�܉������;M�l(����s�=_�����  �D������]�r��v�3ެ"��p8���0dY�8/����v�uuu�j�X�l�����x��UHODDDDDDD�]��7L�:�逃� """"�Xp'"""""�)�����r\��X�lY�����J���n����6]�'���h4���������
�PSS���rX�V���+V�Z�����7��,ːe� ���&3,�V#���TLFDDDD�>Q� DDDDDDT�fC�}ժU���{����	ѽ��,����������,���`@ss3���a0���L&��ݍݻw#��ĳ��v�{�X�re!��$I�,ǟ�B""""���	�DDDDDD��L/�������/��'��>644�����[{�K�����t*&Ѭf�Z��ֆ��!g}C8`ǎ���������7�����x����THNDDDDDDD�W���G��r2�B"""""���	�DDDDDD��L/�ϛ7w�uW�ܞH$��с�����m6���Xn'*0APUU���6X�֬�$�ItuuaϞ=H~���i�������ͅ�KDDDDDDD4�,��9�V+ʖq:""""��Xp'"""""�I���vQ�v�Z�z뭨�� �|>�ر�`0��N���F455A��2.�C�ף������j�oX����}�v��~ @}}=n��v�]���Q��������&�6T�r�i*$!""""*���#""""""��L.�;�N�t�MX�x1  �J���ccc\SQQ���jh4�B�$�C���0��������7�L����x.��d�e�]�E��{�9��,DDDDDDDD�"IDq�|J˪�� ;J�t��NDDDDDD�4���,��wޙ.���a�ر��v�����V��ձ�NT��Z-���|��v�؁'�x۷o �Z�
w�u�Ν[ȨDDDDDDDD�e9c���Y��ÏR)��Xp'"""""������5k���o���,�Į]���3�����7o�f�
i�H	�Պ��68�άE���:~��_C�eTUU��[o�ڵk���������f��� `9a�
I�������DDDDDDt@3�ܮ��p���c����j�H$������`�7�Ƨ�WWWglLD�K�Ѡ��MMMY�������nlذ^�:��]v��կ�`0����������f#I�2�Y�W��������8�]y""""""�j����n7n���|�� �P(��;w"
e=�����̓�d*dL"�!�͆��6���g�x2�ēO>�?� p�	'��[oEUUU!c�,�m膶����������H},�Q��Zn_�l~��c޼y ���Qttt �Hd���h0g�444pj;���h��Ѐ��Fh4���k�Z���;x�� ---���;�t��BG%""""""�Y(���OW!	���j(u�퍈�f���m�y�0�L��b>dAP;F^�%#h�v����J�L,����}�s��� �"$IBOO�^o��V+�����
�����n�#�J���--->&�����c��.��j�w��]<��x��WUJLDDDDDDD��$I�6�Ǯ����TJD���hB�`S;����
����'Q�Ѥ��H�E�λ�X`R��>MO.�<�;�#o����JI�c�ŭ+�
I���X}]��;�S;��]I�{�3�ܮ�jq�u��N  ��qtvv"���8NTVV�����1�����86n܈�+W�SNɘ�L&�q�F�~��hhh�5�\��s���D2��I�������(�d9s��~N3�M��w�R!�¯��>�_�v*q����j� "�)��qD����h��{8��ϓ:wf��������H�]I�ϰr��b�����t����cǎY������c��h��e��������K/���� �Y�����a�X
��������fI�2�YO^�B"""""u��NDDDDDD3��^UU�[o�K�, ����T*�\�Áy���h4:&����>� �nݚ�1�V�͛7㥗^ q���;PSSS�DDDDDDD4d��nn?A�$DDDDD�b�������h�������6�v�mhhh�,�������`�y� ���s�́(�)2�l�D��SOᥗ^ʸ	FE���cӦMH$����-�܂�s�%0�V�	��à��S!�z��=�,6���sn��f8�R)�޽^�7�<�V���fTVV�������ￏ'�x�@ �c�P�>�(FGGQ^^���X�b�
)�������h&�(�l'�Q'�JXp'"""""����yx\�����9U�*I�ݒ-/�,������`l����n����,�$4	!M��<7�����y���Nr!@H�z�!���\v� �lY���/��?�(���RU��z=r�~��|$�W}�{��L,�_}��z�����z��t��Q�Q����j������0�544��������4j�4M���jll����O<�M�69�     d*۶G��\|�I    �Pp   �)(���a����}��'�4
�t��1E��Q����J�ǁ� ������~�im߾}Ԟ��і-[�w�^����~��ڼy�)    @&5�]���%r�Ls    �
�    0�dZ��4M=������%S�����G7{�l͞=[�a8@I&���o�-[�(�L�����һﾫ>�@�t�-���_��L���     ����)��%����   R�W�    `
��r��?��/�\���٩���QS�<����U\\�DL il���z�gG���������+��/~�z�G�v���	     2�XS�s/Y�@   ��   `�ȴr����������.�$�8qB�������|�?����S@�hllԏ�cutt�X7C���z��%I�^z����o+++ˉ�      C�Up�^�R���    �G�    ��L+�{�^}�{�Ӆ^(۶��ܬ���Q���婺�Z�ǁ� 2Ioo�~򓟨��vĺa���ճ�>+˲�f������|>�CI    @&�m{�m��V�J   �w    �p�Vn���֓O>�s�=w�����3���bUVV��r9�@&�F�z��cǎQ{�pXO?����-[����\9     ������/��  ����;    d�L+����������/_.۶��Р���Q�M�>]�gϖa���,��+����^{m�$�D"��{N�hTg�}�����+''ǡ�      ��Up�Y�FF6�5    �Qp   ��i����<��?ТE�dY����5000��0TQQ��ӧ;��T����_V2������3�(
iѢE������:�     ���|s����:��    �C�    2P���?��^YY9\nq���VUU�
J	`�ٳg��{�9E��g��~���)Pr     �m�)��K68�   H-
�    �a2����z���~W���W2�T]]����c<����(�H��Ǐ�?��7ݘ���{NZ�p��z�)egg;�     �����.I9k.�<�    �C�    2H����n����okɒ%J$:v�B�Јc<�������J	`�����O�S���X7MS?�����߯E�驧��g     8e�m�*��9����   �A�    2D���W�Z�d2��Ǐ+�g_�44�}������r(% �����O?�����i����u�9��'���)k     �Y�5j-w��$   R��;    d�L+����G}Tk֬�eY���W8q���UUUEQ �����~򓟨��yĺa��/~�`0�+V�����r(%     H'9�]�r?w��ہ4   @jPp   �4�����zHk׮�m�jhhP0qLvv����)��t�ᰞ}�Y555�X�m[�=����>������a�     �¶�Q%wW~��W�q(   0�(�   @˴r�$���Z�~�p�}ppp�~nn�����fB�I*���g�U}}��u�0��s�)�jݺu�뮻�     ��XS�����I   �Ԡ�    i*���r����Jٶ���&������7o�\.�C	���b1���?����G�۶����������u�u�9�     �˲F��/�T��p  ��>�    IDAT �P�    eb�}�ڵ��[$I�������������J�&���b��^x�Q�����yY����[6lp&      H�m����*���+J   L,Z    �f2�ܾd�=��2C---���������s�Rn�vb�����Q%���������j�ʕ�     i�/���$   &�     H#�Xn�={��x�	��n������{�~vv6�����'�744�X��ڲe��n��q͛7ϡ�     `��,kԚ��KS   H�    �&2�ܞ����}�{������S{{��}�ϧy����r9� �G<�/��'N�Xokk�믿���l=��S*))q(!     ��ƚ��1K޳9�   �X�    db�=++KO>��������4j޼yr��%���D��sϩ��c�z]]�v�ء��b=����|%     ��XS��6\�@   `bQp   �I.��i����-Z�h4�����<������xL	 �/
��g�Uww���]�v���V���z��d�<m     F���{�%$   &��   �$���vI���u�*�H����J&��{��d���A=��3���^3MS[�nU{{�V�^�;����     `2��!!˪�V��*�    ��;    LR�Zn���?�k��V�e���^�Xlx��v���JYYY&��700��^�pxx��v��_V8���_�68�     LFcMq�[��    ��t     �h�Zn���ԃ>(IjllT(�3C�z�N�������/�K�v�mr����3MS�?����n}�k_SCC�jkkN
`�J�6������|��$ٶb�p�3lu��KE�=�1\Sץ@rt9�I�x��   �5�=��u���:�   ��   `���r����w��y�^���j```���9s���J Ψ��ׯ�k��_��Ð44��W���n��&}����#�<���~����l[v$������[Q�#8"
)4�
�   �²,�\�k���^�D{�C�   ��e:     �'�Zn7MS�>�������ק����3f�Paa�C� �YЫ��:b���O[�nUii����Ox     ���x��i*�΄   & w    �$2��.I7�t�V�^�H$����{���*++s( L۷o�|0|�0;vL�9眣��˹p     `R�m{�Z�ŗ9�   ��~   �I ���k֬��7߬d2����Ӆ�~�f͚�`: �<~��ߩ��P�-�4t����~[3f��5�\����w�u8%     p�eYr�\#ּ�,���Dɞn�R �$ۖm%d'��?��JJVR�e}�-�Vb��d��5CÔ㏿�����uS��=�a����6����n    pر�2��>}�t}��_�i����W,���|�;w��T  ٶ��^zIw�u���Ћ/��{�G?���������pR     �4۶G<�j�\��+��􂃩  �ȶ��caY���xTV"&;���N��f�.�,�n�w��W�;K��+��.�H?gTpO�<�U�v�����DX��K�"�|%�>���/}B�F_�
 2A��uV,��X��4�+/Զy\�0��ɨV52Q�g�J���r����w��]��婽�]�{�G���5e ��x<�_�������'�O%�͛7���7��M��ξh      �5���e�(� N�mˊ�eEC�baY�X���'.��£�Ð�������G�̬l.�I|VgTp{r�㋾1^Y�^VY�ܹEN�W8  R���U��N�W{\�t�)'/:@��˔r�$�s�=���������ۇ�M�Tee�<�<���^��w�=��rppPo���֭[���O�����pJ     0���t @��Q%���B{48Tf�-�c�۶�,�.�\�\�>�\^�Lo�d��P`�9��;    `�dR�}͚5��+�����<bo֬Y���v( ��'Nh˖-��$M�9t��͛�+��B����[o��pJ       @���Y����A%Ã�z2�D��	%B�R�_����fV�P������pQ����N    `Ȥr{aa�|�Aٶ��Ǐ+�H���(��| e�޽z����o�\.���k�D"��׾��ӧ;�       0�ٖ��ź�nګp�~E���L�r�Xl�V2T��]��c
7�Q��A�z[dEN��,
�    �r�7c��a衇Raa�Z[[�D��rrr4s�L�@�ٺu��=:|�4M��W�Rnn���o����       �?����v��>R��V�Y����҆m۲�!���n=�P�E;��`%��L�    �ve�?ͮ��*�^�Z���^�x<�;w��p0 �˲��_�Z}}}�k�`Po����>�l�t�M�       8͎G�P���BM{�iV2<(۶����d\�@����n�Q����n���˜    �Q���;�H$���2�n��̙#���`: H_�PH���/�H$$�\=t�u�M7iѢE'       ����+�߮p����)�ݤd$�t��g۶�~E;�nܣhG��^ɶ��d
�    �3��x��o}KYYYjnnV<�+//���w0 ����V���k÷].�^}�UY��G}T����       L8�R"УH[����n��N���l�R"ثhG�B�{�j�:��    g쮻�Ree����4000�^XX�iӦ9� 2�Ν;USS3|�0mٲE�����L       �(V<�Xo�BM{�<�dx@�m;ƶ��v)|�����o��L8Hk�    gdٲe�ꪫ�D���6���z5{�l�@�y�W���9|���K������-_���d       �qc�C��[��(L�+Q��Eᦽ�v�3�8M�    �-++K<��$���Q�eI�*\QQ!�䟝 0�b��^|�E��qIC?o�~�m�B!=��C���v8!       �t�VR����Mk�����dۖ��'*薘��2�    ��v뭷���\����D"��3f̠d	 ���C�����m�4���/���L��s���        �ÎG����n���9	�Ȋ��W�e���m9	��(�    NKUU����uuu���~���:� 2��ݻ����ۡPH۷o�ƍ�|�r�       N��(�y|����&�J:	ȊG�nR�i��'��>w    �g�r�����4M����X�3g��� `���o~�����ۻv�R �C=$���`2       �'�baE;�i9�D�G�m;	)d'���M��m�����;    �3���k5�|���+��Ϟ=[���d 0u��a�����/|�\.mٲEeee���N       �KV<�hG��-�tSl��l+�x_�����o�l��H��A�    �L�>]7�|�"��:;;�׋��UPP�`2 �z���������ڵk����ZUUU9�       �1;W��ahb{���8�d�dB�����)>�A�w    �g`�|�Ay�^555O����Ryy��� `j���������۷oW4�< ���?       p�m%�mQ�i��]Ll�'��qź��&��FLq��    8e6l������եp8,i��^QQ!���p: ���ɤ����]�dR��r�����F,ЦM�N       SS"Эp�~���d3����*�Q�H�Y���q GPp    ��߯��K�x\����륥����q0 ���Mo�������^9rD��~����L       S�)r␢����q�� �%Ã
����$
�    �Sr�-�(??_��Ͳ��)YYY*++s8 @��z�-�8qB���5�|�My�^�q�'      ��g'�v�+�rP�h��8� �W�p:
�2�    �j���ڴi�zzz4888b�4��% L�ei˖-J&���J����~�z-\���t       ���^�[�+�v:
2�m%�nR��!Y���q�	G    ���^��������b��~S �R[[��~��������W��ސ       �̎Gi�U��Nv2�tL�hP��m�l��8��q;     0��w�yZ�j�N�8�Db�9�ǣ��r�� ����ok���*--�i�z��t����.�믿�t<       ���N%�Nǘ�q%B�J��t)�S"�+3T�˔ǎ�cHv"*+��c�0L%�,%�Iٶ�H,&Ó#۝����Ζ�������/��p���i�1��ض�x_���>y�͕�c(2w    �I��n}�K_R,Sw��.�8k�,�\.� N&�L�7�����.��p8������;��{ｧP(�tD       �YE�dE�JFNGI	+R���b=�r�:��T��wŕ�%���P�*((Pnn��8��E"*�V������/�Ԡ�Ѡ����P��9�Γ��R�'{���͊Gn=,O�te͒��{L6�    'u�Wj��٪�����K�(??��d �O��Р�>�H�{�$�w��}�ݧo�Q?���N       �0�-�R���d��4�*�תp�!��AE�W�P�߭Y3g��
���'<�����Sii�'��۫��mj������g)��.όE��^"��x³:)�߮ddP��y2=>�� も;    `L~�_7�t�500tiE�˥�3g:� p*~���묳�Rnn���o��k��V����:;;��       �py�+�R�������c[��U��Fy�fMwjδ|U/�Vy��3�
EEE***�ҥK��,�Rkk��{F��}jO�ș����䛱@2L�?+R�堲�g˝��o �w    ��n��6��~9rdx���\���T �S�����N�_�$��ѣ:���y�f���?t8       d�痧x�b�MNG9e��
}_y����ւ�
-\�P��UNG�ij֬Y�5k�.��Z0���o�n��TK̯��J�T���h��Yǋm[�v7*�WִJ.*�H_��    �2}�tmܸQ��݊F�����l9� �Y�ٳG+W�Tee�L��k���n�A������:��      @���Ɋ��:elVB���J6��,uj�"-[�L���O��\.��n��n�<���_~�,K�e�/�Lʲ,%�I%	%	��q%��3Δ����+Wj�ʡ���yQ�vw��=[�y({�Ҵ���+�r@޲yr���
�    �Q6o�,I���^+//��� �����V_��Wd�������ѡ;�CO=����        �xK+e�²����-��(z�m�I6i�9����r�\g���G999��Ζ������UVV��^�Ls|K�e)�)�)�*�����]�E~~�֮]���l��ѣ��ݗUΕ=�|�\ �����v2�h[�<E��)��t�3��    a֬Y���K��ڪD"!I*((���w8 �tttth�ΝZ�f�L��֭[u��kٲeڳg���        s��ӫ9qH�u��O�m+���B�_Wi�^�_v�λq�<�O��L�TNN��~��Gvv���T1MS>�O>�o��d2�`0�P(�`0�@ �@ 0b:�'1C,Ђ$I���ڵ�t$Z,ͿL����kI۶�i�	(��R�y�ol R��;    `�[o�U�dR===���,�9s�é  g��7�Ԓ%K����P(�Ç��n�c�=�t4       �(�ǧ�is�K�y��oU��~]0�\+6_����>��dee)??_���*((PnnnZ\���r���m�
����������N��***TQQ!۶u������쭒ٕr��'�˘�P�����U���`���    VQQ��.�H---�m[�TZZ*�'=/� ���o��+��az�w��/}I+V��G}�t<       �(��"Y��o��ٖ��+��U-ʋ���׫����n�[���*,,TQQ�I'��#�0��Η��Kz����o���+Z�c,^�X�/V0���D5�R|�_)�by*��qa��8$o�<�r
��|*
�    �a��z������$I�G���� ��]�v������ӕL&�{�n�q����~S       `|d͒)�O�Էo�|�~���+u�����Vegg���D%%%���K�	��%;;[���*//�m�Pww�zzz�?񾹹�ڰ�2m�t��>�����5o��o���J�pl+�h�1y�g˓_�t�Qp    H����u����i��8c����p2 �x�,K[�n�m��&Iڹs���~�Z�J;w�t8       dÐ�t��-e'���@�v����}��5���;N�����*--UII�rrr�%O�3C*((PUU�B��:;;�����e�E�iѢE�����o�'5��_y�\��)Jzl�V��Iv<�����zs�w    �$i��͊F���۳��UTT�p* �x:z���;���jIC%�͛7k׮]Lq      �qf�<�U)�v䌞�M�����gT�ݾ�*+[uJ��z�*--UYY�rssO��SENN��Ν��s�*���S��b'�OYY�6�p����������fȷ���R����t�N��-�'<��C�    �h���jll^�9s���  e�֭����aڵk���~�\�R�v�r:       d�痧x�b�M����`��?xA���u��Ԍ�?�|����b�������t"C�����Wee�zzz��֦��ޓ�Q�����+7�x\o��S}Б%������8��K��d�8$���2�YN�F��    ��7߬h4���~IR~~>S  C���iϞ=Z�|��жm�t�7Rp      �	��/�*�9���]�}�g�?��W^����}�}|>�f̘�3f���id��a*))QII��Ѩ�����ڪx<>���G��]��"���iOh�r��"ӗ���Ɗ�i=,ߌ�dx�N��Qp   �)n֬Y:��FLo/++s0 `����Z�x��n�jjjt�����������       �;m��XXV,|�q��|I�{���+�Jee��������5k�JKKe�8&�_�z��;w�***��٩��f��1���|�z�F����E��y*<�f�5��|`%b
����,���q I��t     �����:E�QH�ޞ���p* �D����Ν;%M�ٱc�n��F�S      @3L�ʪe��1���R�>�[βt}�@�iӦiŊ:��sUVVF�=��PYY�V�\��K����������ƫ��k����?jp��)Lz��d\��dE�.��F�    ����B�[�N����k3f�p0  U�y��K����h��ժ��r8       d.�㕷�r�Z��ڞ��V����ޫ�~�ck�ʕ:�쳕��7�iq*
�l�2-_�\���'=���D_��j�4�K��_�κ�<5��T��VV$�t��;    Le�6m�m����

��q�9 �
��v��!I�m[������_�p*       �l��By
gȎG���լ�?֓_�E_��d�'�t���iժUZ�x�rssS��"??_�/֊+TXXx��,X�Gnݤ�/k��N�R���}\rOF���)��;    LQYYY���+���)i�RzLo���w�Q4�$�رC_|��M��p*       �l���
����_;K��v�rrrNzlaa�V�\��~�q����t�R-]�T~��c�кu�����~��<�=�)?�m[����GQp   �)jÆ���Q__���'Ǽ^�é  �
������q;vL�6mr8       d�x_����F������p�������d�-]����i���P�{�.\x��碢"}����[�����dx �)O�㒻	8Sw    ��L��UW]���nY�%�0TVV�t, ��{�=E�Q��+2B�    IDAT��_W\q�'��       ��zw�Z�_��/I@��H�x|�qn�[���Z�b�������qTVV�U�Vi�ܹ2ͱ+��V��#׮V�{?P���'<9۶i?*+r:
� 
�    0�Y�F3g�Tww���� Lo��)
i׮]��H$�`0�K/���P       �!��A����:���t��kllԳ�>;|���L�w�fΜ)�0R�4MUTThժU*..󘜜�y��"��_���H�S�Ͷ����ʊ����)��;    LA�\s�z{{�H$$I���' 8���S"��az뭷t�UW��	       ���m���Ju��?Nz̶m�t���{�Z�p�<O
"�|>�/^�s�9GYYYcs�z�������Iq±���P�}���15Pp   �)fΜ9Z�d����$I���Lo�).���F���ե��R-[���T       ��l['������H���'=��ri�ƍZ�hQ
��i%%%:��4cƌ1�

��;nв�_k`�R�nlv2�h�Q�ɸ�Q0E��     H��7j``@�hT�� C�y��{�r�\z��u�W��   �L����	  d�dx@�t�zw����UUU�;�Pyy�$����Z�bE�Op�m[�XL�ht��m�J$ß%��C�4e�C�].�<�����VVV��^��1���ri��*--Umm�"������/�Yǎ����r/{X�'ۡ�C�xT����._(��{�ɉ�;    L!n�[�^z���������:�
 0������Z�d����t�����X===NG   ��~������  0�B���Q��c'=�4M]~���k�r���#��>�ŋ�0�T�=#�XL�`P�`P�@@�Hd��>Q���������������\������M�9'Zaa�V�\���:����گ���Cee��O*z���[:ρ�bEC�v��[V-���S�/
�    0�\p���|
��� ��w�Ւ%Kd��jjj�~�z���N�   �.\(�߯��F���:  `�u�������X���L�6M��s���������Ucc��Ν;Q1OK"�P������N\�'�)�i```ĺ��Rnn��~����UPP������;]Os/**Rmm��m^^���o�Җ�U۳^���8�tH"�/��EYų́�F�    ���7O��x<���w8 `2immU}}�*++�w�^]q�z饗dY���    �9�0��  2�m��������>���i����z��x\cc����T\\<�)?�d2���������O�`P�m;���|�w``@'N��$�|>��竨�HEEE�x<��tӦM�����Ç�,���uWk��z��\p�C)����e����/s42w    �"f̘�%K����Ò������ ��m�6UVV*��4M�X�B�w�v:   �4��ޮp8���N��   �+���q�z���I�q�ݺ�t�e����>|X+V�Pvv�x�<%�x\]]]���R��.���H$�H$���I���Wqq��������p����|Z�l�������<j��՚VW����?+o��%ӹp��Y��+WN�c��(�   ��q�����\.9	 0	:tH���***�{ｧ�7Rp   pƚ��TXX���\�A��   ��D�[��r���9�1����򗿬�����؉�<�+V�4�3Lzr�x\������Toooڗ�?I P Pcc��^��M��iӦM�+^��y��������V�dr�~UU��ZP�o����?&��w$�mۊv�o�"��#��&�'    `�p�\������-I*))���r8 `2�m[۷o�$�8qB�V����l    ��D"����B!��   ��ȉC:���O,��s�9z��'?s��c�`P�������l�Vww���ۧ>�@�VOOOF���R4UKK�jjj�s�N577+�;k���R-_�\>���xII���r����J��9�n�m%�l˱�L�   `
8������d�JJJ�� ��v�ޭh4*�˥={�h�ڵNG   ��/_���?_�f�r:
  �	����x����Oz�ڵk��(''����ѡ���3z��E�Q544h���:p��z{{��q�]8���ǵm�6<xp�}_rssu�窠�`�^NN��v�u*����8�@�!V,�hW�c�Gf��    S�������#I��˓��q8 `2�F�ڳg�$i���Z�n�É    �����4�j	{����￯��f��  ����:��Jt��o��n��f�v�m�v5庺:��������~m߾]�����b�+�ض���.�۷O;w�Tkk�,krL%w��Z�t��������m���?U���$=�t8v~d
�    ��>~W������N H;w�4Tv�1cS   |&����F�÷�Ќ3��   H[����������������˲t��A����t���n}��Gڻw�� ,��p8��G�j۶mjhh�����`�.\����1�n��z�=��M{H7$�Ӭd��ߌ�9
�    ��.����a��qy<���9	 �������,�0�m�6}��w:   �4�v��H$��^.Y�D���L  i�o������'-��������-Z4!�F�:t�l���c{zz�����g4�R"�Pcc��o߮���IQt�;w��ϟ?���7^�s��C���)N5ĶmE;��N&9?2w    �p_|��T���"��p" @�صk�$���Q�֭�!    NY"�Q ڳg��9B�
  ����^����od'�c�O�6M��ַ4gΜ���ק�����wuui�Νڿ����f�j,�R[[�v�ء��%�����u�9��4GW��޴QK�^S��C�Iv2�XW�#�Ff��    ���kɒ%�/;� �N��ۧp8,˲�FO:       2���7t�7�N�}�9s����WYYYJ�477���{����jjjt��A���䘪�ɤ�c������D��RRRrҒ�U�6jQ�oi9�@2)�Sb�ˑs#sPp   �v�E)
ɶm���)++��H �4�ǵw�^��]�v��/v:       �D�����kd�#c�WTT�GQ^^^Js>|X�PH�hT����裏400��S]"�P]]�v�ڥ�.��EEEZ�d�\.ר��ޤʺ_(�zādR���w�SA�    2�ڵk���/��� ����C�1���Ѕ^(�0N       +�X���$+s�ܹ��׿����'�"�w�^�ܹSmmm)??�$����ڿ�"g��Z�x�%��n�F3>�Xg}�sٶ�h�q��)�Ho�    C�������n���� HC���joo�i��������       &�~L�p���1�����裏:Rn�X,�eY��#���h���jii��@��㒻i���v�u*��oJv�<�)�w"��Ef��    ꢋ.R �m�***b�. ��ٳG��o�>]t�E�      �������R������g��< �ϗ�d��ɤ���TSS�`0����n�����y��ʎ�R�+��&+����w    �P]t����%IEEE� ��={�Ȳ,uww��/t:       �;;ӱ��׊�s���z�ᇕ����dH'��������ؘ�i�Z�hѨ�gn�[���E��/�����ѮɁ��Ho�    ���kѢE
�z�L�  ����A?~\�i���ONG      ��c�:��{5p��1���#�(???����l�VCC���ۧh4��s������z�zNN���|��QJ�H�+>О��"�Qp   ��r�Jʶm: �jjj$I���Ӛ5kN       �����g�����҆TSS��۷+�L�8�U__�v�ޭ�����\s���^RR��V�hp�R�G��'d�#)?/�w    �@+W�T�$�����4 �Lp��!��quww����w:       ����[t���1�L���_���b�����r��w��o��`0��HG�DB����e�v��[QQ����Q���պ��S�c�,�44�>�Ր�s"�Qp   �c���-[�`0(��'���t$ @��b����i�r��\!      @ڋ�ժ���C:I���K.ѬY�F���檠�@555ںu�zzzRi���Y{��U<O�9�:�1��?��5:�c�)�"I�H@��Δ�鋂;    d���j�\.ٶ��v ��:p����U�V9�       N����N�P����w��:묓�������XG����ut��,����߯?�P�@ %�3C�-Rvv���뾸Q�����L]�^�b�-�����鉂;    d�U�VippP��� W�V,S{{�V�^�t       8m���Wn�?����ޝ��u�w��a
��6�Vq'K�H����"%y���v����ĉ��q�8�v;Q�y�NғN&��Y��N2r�I<��v����II����*����ګ���~��"(�E�(��y�98��ZP��s��ի�y�曚��r)�z�400Pʘ�1�tZǎ���dE�\.mذA��q�á���Ǖ<���q���);3RњX�hp   ��e���qy�^y<��  jH6�ջﾫ|>�e˖�n��E       ��讯k���E������G]�v�]---���Ү]�t���ۍ����t��)W����Ӛ5k
���>yw��'vU$�Fl\�l��5��p
    jHcc��-[�l6��� ��8y�l6�����j�*��       ��$�Nj�/��p8���z�`�녰�ljnn�aڽ{�>�\.w��6����g�Vl����Vuvv��^�Z����NW��^z�g&/V�'�   ���s�=���D�; �,���e�u��w[       n��Mk�?�|&Yp��r�'����.Y���&9��?СC�dF��Fmҙ3gd�f�k�X�B�`�`��;?$ߛ�U2�e�pE.Snn�b�����    5d�֭����x<%�� �+��Ο?�d2�����8       p���e�]<Z�ڣ�>�H$R���@@N�S�����ۧD"Q�:X����*��n�ٴ~�z9�΂��|�����ֿVf�T��~,N4�   @ٸq���抮� �T���d���r���x��       7;��.?��E�mڴI+W�,{�߯P(���~[�w����t�kbq�ɓ'�����x�v�ڂ�p8��KbJ�,k��g�2b��Ņw    ����r�\2MS���V� ԰3g�H�Ξ=�6X�       �/77��?��d�����i۶m���z��Ԥ3g��^���HE�:MMMU�ɽ��YK�.-߶u���?'�������H��K�w    �����F����4� �jvvV�����      @���_Vfj�`��vkǎ�ۭi�t�\jii�����٣���[��cjjJ�O�.{��ʕ+��z�?��#J��We��Af.�,����   �F���*����Q6���8 ���ק\.�իW[       �8{Xc{��赇~X�@�
��vE"MNNj׮]:z��Ց`���	��������кu�
���=���@Y�P�]�Q�    P#֬Y�l6[� j_�l6�2���N��q       ���3t����ͳ�ׯתU�,Hu}���2C�w���Ç��嬎���j`��M��`P�[�lV��_V�����F�*R��    P�~���$�� ����A��i��;      ��t�~Ss�.����-Ht󚚚�p8���/�СC2��H����!��������z�?�s�������?(;;*3�b��   ����*�J�����v[ P���Ο?���imذ��8       p���Y�ݯ��l6=��r�\�Z�`0(�өW_}U���S<�:*h``@SSSe���ph͚5�HD��2���Afΐ�H-,4�   @���U"�P0�:
 ���0�]���(       p�K���g��6lPGG��nOCC�B���;�ݻw�����4M�>}����ZZZ
�?������սVvvL2����F�;    Ԁ���+�J�����( �:200 ��.��iu       x_��K�>�\�xcc��o�nA���x<jjjR__�^x�[	e���t��Ie�ٲ�X�zu�g�v�]YR�r��~����HLW���    ��9�Nutt�f����[ PG����F566���V��       �d�u��_,z����;\.�ZZZ444�ݻw����VGB��i�>}Z�i�e~�˥������שi���f1ٙ����F�;    ,r+V�P.�����Οy ��:w���ǵf���       �&<�Ĺ#�˗/WOO����n����I���ڵk��=ju$����LY2ttt����`�G�S���e��A�lJ��ي�Bu��    �U�V)�H�{; �/^T:�֪U���      ���3s��W
ƝN�x�UVss��О={t��!�r9�#��599Y��m6��/_^0��ڪձCR�2_O��hE꠺��Y n��M+��T>W.�P.U.9�|:�|&U�$�MΆ����9�9|Aٽ�r�����T�  P����577�����  ��ŋe���=      �r�/|]������[���$�F$�$����r�\ھ}��n�ũP*}}}ڼy�<O��nnnV8����U�O=�E�8�[�;?\���%c�g�dw�&��A�;Prs3J]�Wj�O��}�L\PvvT��Ae��2��%�isz�
���3�&wS��KV˳t��K��ӺB6'o�   J���S�|^>���( �:411�D"!��]LӴ8      �z�O'4����744h�ƍ$�^0�$:tH�ij�֭jh�ix�3CgΜ)����+��[o]5��بu����)���zl�&�n�.{T/܁b�J^:���74w��Wz�O��X�ie&/)3y��u��!wK�|]��s���#�=r��T8)  ����ڪD"!��eu @2MS�.]Rww����4:�ѡ       *ol��ھ}����n�������o+�Hh˖-jjj�8n������U���Ң����Ɵzx����ny6|��5�e�&�t�fw���S}�����%�N�W��%�h��;2��ձn���)=6��؀f�������&5�ܣƵ*��5����F   ����U�C~���( �:v��%��Ϊ���w       �����?�V�xss�֬YcA����x��x��߯���u�]���:nх�D�r�����������������|�4��%��������"��R�䋊�گ��J���:R��)EO�U��^I����V�?�@�c
�Tv���   �cŊJ&��D"VG Ա�/*�Nkٲe:|���q       ԙ��\t��-[��f�Y���9�N���hhhH��V�^�U�VY�����߯M�6��뼡�A����j|�[u����%�W��������T���	ͼ���y�����"�f�k�l6�|>��������L&#�0��f��f˖��e�U��W5��ߐ��S�����l�����e�  �,_�\�T��c ���Ȉ$��
      @��3I]����`���Y˗/�|�E�n����E333ڳg�:;;���ku,,@,���:;;K>wwwwA����S��Ԁ��l�����\:�|&Ɇ�u�w�ʘ���'�j捿�̛�Wfj�ds766���E����D"
��
�D"
��|�z��x<��0���)�LjnnN�hT��Ӛ���������5>>���)��٠��$=�G��{t�ٟWC�F���������u��
  ԟ��.I���8	 ������1uw�      @eMxV����7o� ���D477�={�(j�֭�������8�����K~ϸ��A---����j���u0���    IDAT�W�Y�PI�c�&�n^V�:�>4�U"9xB�����Q��B�B!uvv���K������Pkk�|��dr:�
�
��}�a��ؘ���588���A�����3�B�]<����4�ܯ��y�"�~J-��<KV��|   �͒%K��> ��V6����P.��:      �:1��cMMMZ�b�i�+'u�߿_n�[۷o���8�'����ٳڰaC�����*hp��eU��=1%wS�d����2��4y�YM���çni�ǣ���\�R+W�Ԋ+n�hn�ө��v���kӦM�g�Y]�tI�Ν����Ξ=����ϟ:���~M�����<���~ZM��3���|   U��r)���� �*022�X,���v��D:       ���;�4w�X��{�pkB��$����2C[�nUcc�ũ0���)MOO��@�T��B��fgg�tc������t�Y�z�2s�rɨ���A����@�����MyNf�X�s].�V�\����k���Z�|��?
��kZ�r�v��!I�����ӧu��i�:uJ3337?�i*�wP񾃺��ϫ����?������
   ���٩l6[� �exxX�TJ4�      ���~�`���i�ʕ��MWN�>~��R��6m�T�&j�����6o�\�Һ��
ܗ.]����+s��$�i���@��QM��/4���>���F"mܸQ�6m�ڵk�r�ʔ�z��a�w�}���$��܉'t��1���+����<�dT�����}�T�������O����  X���ڔJ����fu  4::�L&���v��  �Y����\.��7�9s���y�r9�c    ����ܧ٣�_����p8,HT�\.�\.�����F��۫��N�c����422���������$�ϧd2y����^�c|R���ֻVnnF2�mqo����O-�
�Nk�K�/��S�~ޒ%K�m�6mܸQ���%_U�ش�����];w�T"��������o�w�Q6���9���(���<���|�ߩ������/sr  ��Y�d�2��<��Q  P.����V�^mu �Mrv���ٿ�:�%�[��o�����hu    X4�v����^?��p���עD���p(�hddD�O�VOO�W�.hɒ%%_�t�R�;w���za�K��+i�k���rɨ��Au��(���9]�����K&�H��s�ᰶl٢-[�h�ʕu��>�߯{�W��{��٬�;��^{M'N����m���u��/h����m����'��\Av=  �OSS��n7� Ucll��G       ��42�|�;�+W���� Q���l
�Ú��ծ]���֦����Xu�0������.]�T.\P>������1M������4�u�w��Rç5�_��ߖ�3n�x�á�7��Voo��v��X������X,�C������s�������t���Ւ'���~�Kr66U 5  @i455���Z �����Y      @�~�ȈM��[�΂4hnnV.�Ӌ/�(�߯-[��|qܼ��!utt��r�lN�ө����� �s���y[��{JV��\bFj�K6�+��@�d��5���4��������V=��Cz��+����ܹS;w��ٳgu�������f��}^>����C����%O|^�?�K��  �B8�� PU���d��N��Ɵ�       ����������W>�w������o\�v�-NUr������|������^���$zT3*o��i�KF��#4��ꙹ�l�ҭ$*�\2��������*�����{zz���k�����^F�V�ҪU���OZ����v�ڥ����>'��k������T�?�Z���.��S��   
�hp T���1%�I������j       �PٙE��U0�n�:�l6�Z~�_�t��a���[������T�exxX���%��=���*�J]5~w�]�Rqٽ��7��������fħ��� o�:��Vǹ���jl�k��~UFt������ڼy��x≒�����|>=���z�G��oh��ݺt��u�c�'u�;_�ؾ?Q�����[~�Bi  n^cc��|>��Q  x�����       �f���2s�'H�Y�Ƃ4��+�2�y�%	�s�=jnn�8U}��rQwwwI�]�d�.\�p��]z���k���Y�Z����J|���Q��kn?/�4�=+oG�l������~Y���J���l6�6oެ��ђ%K*��8�N�{ｺ��{u��)}�{�����u��=����Q�x\�����[vW��  �X[[���|IW� p�L���Ą�����      �FM�V�X[[���ip3�n��n�Ξ=���zK�ׯWWW�ձj��А:;;�p8J6g�w�ݮ��E��Jqy#�|6%��S��Aut�0bJO�����Qz���KVK#��ե�����$�漏�����{�я~TmmmL����۫��^�>}Z�������^��ѓ�t�+�ն����ԯ����0  ��ҥK9b P�&''�t�R�c       �A���J^z�`|�ʕ��B9E"]�|Y}}}���ѪU���U����ؘ���K6���Q0T4�j�Υ^]JF��KV���ܬ�!���:Ft\�ɋ�dTٙ�"�e�5q�[���_����C{{{��O}J���
�[�~�z�_�^�N�������ҥK�>��}��5u�����o(��G+�  �PKKKIW� P*SSS�z�p      @�M��7EǗ/_^� �-6�M�PH333ڻw�ZZZ�q�F6�*�����6�K�ݫ���}��5z��k��'KZ�Z�dT�В��@u��U%;;�����33#�{�r4�*�)5|Z�J�=t��-_�\���'�f͚
%C������_��:��}�{���CvzX���'���g���'g���I  �I0���:  ����t�#      �қ>�\�XKK�������	��2C{��U0�֭[e�ۭ�U3�ɤfff�K6gKK������1�5�gi�S1��K6�Fjw�P5���u�ۯH�����W6����LS���@�������z�駵m�6V�-b6�M��w��l٢^xA/���2�̼��<��5��.u���W���K�  ������ �JSSS|F      ��2S�J�^0���mA�Z$�$8p@v�]۶m��S��:122R�w�ǣ@ �X,v����]����n(Y�k���\*.��E-��%�
F|J�ɋ7�X3�Sj��{�p�$3qAg~}�.>���6���v�رC_��״}�vn���˥�����_�U�w�}��w5���Ə���?-#1]��   �����:  ���d���1       Ԙ���F*���e�,H�r�����|z������/+�HXiћ��R6�-����ckV�R��[%�SL>/{X�wX.77����='�I*=q�,y&^�sf��'����5k��+_��>��O����%���S?�S��������>v��wu�+[��B�   ����  �(�Hhnn��       j��[�P0��x���fA������ױcǴo�>MLLXi����+�MMMc�CK27����ȥip�4��R�tB鱁[��ˈOɈ��.K6����չo��r�h�Ǹ�n�؏����������,YmT���^}��_�����p�����9���G4��_���U0!  �W�� �Z333,�      P2�lJ��]]]��l$B���n�B!�={V/������(]�|��������V4$KZ��|*Q�4��a�|&���~�f����L]*�q���:�l����e��\it~ꩧxSTg\.�>���~����5��̜�������Ne��]�  p�@ ��R @՚��R0�:      ��E�La�lGG�i`�ө��]�|Y{��U__�Ց��������D
��X�L��ֹ�i��p�l����0�i�.���Nצi*=~Nfθ�9�_�[���}J/z����3������/������`�����3�<�'�|��d�S�u�˛��
�  ��n����[ �y�����      �d���ooo�pX�f�)+�i�޽:z��Lv�)���%��X�{SS���'KZ��\	6FFusZ ����;{[M��72J�Ȼd���,͜����w����}LGG�>��ϱ��s:�z��u�=������46V|����������'���G?[�  ��9��9 �^�hTmmmV�      @�˥b���*��+�����w>/3oHfN�9ew�$�Sv�_O@v_@NX6;�Z��=c
���A���2C���W0��w�-��au��5>>������7��_�cFJV��|:Q�
���QY��������܎\2�����M]7���Y����5�ή��m6�v�ءO|�4���+W��_���}�Y9r��c�ٔ����V��u�����tW8%  (���dʻm���R<sӏ|0 �j�hTz�*s�ʔ�Jɽ�{�     ���畍�*;3�llR����2�_����a�MΆ���6�#��{�Y*+77��so�/]�Ԃ4�FWN=x��v��m�&��cq��L&�H$JvZ�����W"qu�y�?�f^��KR��k�����Ԡ��ٲ̝�����_x����ϩ��>��P�c0�~�>�����;�,GL��׫�}�sZ�f������0��J0�珔>��?��r4�j ��&��)�~s)oU�/������e[��E  TZ4]��P�R}�L���I�; �R�lVccc���joo�:   �h�S	�����idoBӔ�����V��9�Mr7����L��9 3�+��׺Ҹ}��a���[�*X���LNN���]�B�PA��ڕ�z��y�[W��ε�FFfΐ�At�*���FlB��XYkd��+�M�{=���N��������ե_��_����c������:�c�'_ԩ_yH�ɋL  jUCC;� �Z,�T<  �0C��������   (��)q�MEO�Wz�Bi�ۯeJF|Js�R��>e&.J�Y�:�e�����_�W����A�`PǏ׾}�4>>nu��1==]�����w�ݒ�)&�M���C�;*"��V���4�J��-�bo굿�����y��mۦ/}�Kjii)wLԠ��n}�+_�ƍ�}Lr��N}��]<V�d  �y<� U-�H��      n���)9|J�3/+;3,�2�LRs��)zz���DEj��g���v577[�����V(ҹs�o�>Y�r�XL�a�l�P(Tt��,���|��ZF�;��42J���Y����lJ���W�������32�t��m6��~�i�����<OE2�6y�^�����v��9�c2�C:��+z|O� �Z�p8� PՒ�$��      pK�ظ�'���ɥE;��S	�Ͼ���Ǌn��
2M%�)njj�~n���P(��Ȉ��ݫ��>�#Y�4͒���v���]�{{5Kͤ�����e��5��J���fs3�ώ�Z���������Gy<}�����w�]�|�]v�]��ԧ�l�2=��EW��Q���Ǵ����"[?aAJ  �^�[fCCYk�����n�� ������ c���P�߹-     P�LSJ_�S�r�*�c�u�Rf�r�)5,�"�/`u�����'#>U0���6�M�pX�XL�w�V[[�6n�Xw'�NOO����d�566*����}y[Po��{�%�s-vp�mtD��2S�ʥ���N����']~���^�B���?����
'C=�����֦o|����L#���)�����?cAB  p���len�s8v����`W\ @�[p���2��V      �-0���P66nu��T\���,g���8u'1�z��H$R�$�5MMM2C/����e˖���FK:_ ����Uc]]]2����kcIk}�ma]��ie�c�7M���o���!�������z�ghnGY�\�R_���]1j�s:�͟��+߮p2  �ع\.���9 �n���      �13�U��CU��~��7�x]�KVG�;s�.:�+��*
��p����z�W
v"�E�dR�l�d�566�95$/��F1�������zEG��̦���`Y��=_�����s�N�����U+�zzz��/~�U|����v}�K_RGGG��f�й?���x�U8  X��n��  ��T*eu      T9��*����Ĵ�Qn�4M%/Ufz��(u%9|��8�_(5��/�ǣ#G�h���%��ڔ�������s�d5�ϱ�N����g����YR~b��+����%I�V��'>�	IҚ5k���EW�����ojǎjk+~L����ܟ~N��U�t  `�r:�VG  ��hp     ������+��Y���܅�2f�w��Z�*lpw:���l�^���N�<�}��i|�6��K���v����nv$KVc>��^��@�e���O�YR{b��ɞ�����Ɵx�	9�N=��Cr�\�dC}���z��d��B��$�����y���>���ܟ���n�"۞�pZ  �ذ�; `1��c\     p��.�%#1eu��3M%�Q`�C��V��i�LR��PH6�͂D�'.�K�PH�ϟ�ѣG�n�:-[���X%��vqQCCCA��Ҁ]�KZ��i��{�bw�T>Wv�H�nL����pwV?�p��H$�g�y��Fc��N�:��^zI�G^���q�ۭ�}�c���(�<3�����b��W()  X�hp ,��5��     ���'�+;=bu�[f�s��?"����*5rF2��HĂ4�Wv�]�HD���ڻw������T�D����|����%��%�KZ�Zy��vj�(3���yKJϼ�?t_ð|���k�HDw�q�\.��㎢Ga �011�={�hnnN�`��c�N�>��������|6����a%�)gT  ��y<�#  pC�aX      U(7Ur��1n[>�Pr��1jZr�T��p8\�$�d����F�o�>���;2M��X��0�������P0���$cf�d5�a��E�;J&3yI�l�W����7��>���\���n��������v��JGD�K&�z��500pS+D�N��z�)�����K����Q�r_�� ���M �b��f��      ��cjn�)_�+�b���$#6au���(:N�;�
���d��~>|xўhZ�]܋m��p8�MO��F1V���2hpGI�Qe-x��>�����'����k�@@����7�_���<����B��y���z��7�p8n���CO<�/_^���P�o~�?�  @Q6���  �P&î)      �Zz�r�i�c�T-5�W���`��;�S�X�M6`�+=cԁJ�#z%��������%�Q���J&?�k�mf�Pz�|��f���{������M����;�m8^�|�B�P%b�F�={V���4�/����ڹs�����^O�����1�Q  ð:  7��+      |��7�9cu��˧�L^�:FM�L^*:�b�
=��cڸq��ɤR�T��W�����|:r���߯X,fu���L&K6׼��\�j���q?����ۖ�zoL�3sJ��k�ܿ��M�n�[w�y��N�Ϸ�l���-z,p=���ڳg����K�H�J�{GGG��3?Ѕ?��m�  ���(  ��      ����Ś��/5�.;�A���>���Fچ�=��Cھ}�r����x�#W�z�
:q���ۧ��	�#]W)��\����%)�̕��|�<�#j�-�tB�X������}�S�������]w�uS��.�K���E���d2ڿ�����Dd��J6���ԓO>���֢�����.��o��  X�r��         P2��RcV�(�|6��Ԑ�1jNf�p�H$R0�r��}�v=��#r:��F������r)
�ܹsڳg�.]*~����tI�s��c!_��3���6�ً[g�J[p���Ч�[������m6�֭[������+hŊ���s��Q:tH�@@.��,5�n�>�̻+���|I���K�m{    IDATR  ,>�<;�  ��
      ��L���l�v
�F��VG�)�LRFb�`�X��6�M�6m�c�=&�ۭ���rFn�n�+�httT{��U__�Ց��N�e�f��+����,�����6q�	�,S>=Wњ����@��뮂k�V�RSSӂ����В%KJ5�ҥKڻw��X�[��z���|��dI����?��2Ӭ�  �a�: ����     �+�S�VG(��܌�ɘ�1j����4��>�f�鮻�ғO>���&MOO���X(�ͦp8�X,��{���ѣU���i�%����t�5�m�Y��j�^��˄[b��ΌT�fvzH����|�k;�/��ի���o'j�����٣��Q��������?\����ٯ�3��lE3 ��C�; `1��      ��722��VǨ�4�L.9[t|�=^+V��Ν;��٩��Y�r�R�nY8�az饗t��a�ݳ���������W.U��?y��kw�pK2��dV�B>�̾�я�G.�A�\�򶦷�����-�T�������k��ԩS�D"��l��hmm��?^�~������  Մw �b`���      �.Fl�nv�6b���_	���4�_��ޮ�\�W�V,+iS/p+����8���t'��(��B���@  #>U�Ř9��"ܱ`�TLFb��5�_��~�c���\5�v����[��>�O�֭��y�8�8qB/���\.�\.��q�|�rmٲ�����[�>�\� �jR/ 7�      IF|������42VǨ	��L��[mp����I�=��6nܨd2�T*u[���������ȑ#ڿ�b�2�v~�R6�;��1��/[&Y��Tt�fT�X���`E�͝{SZ�Tww�U�6�M�֭+z�ŭjjjҲe�J6������٣T*�`0hu��l޼�����s��lſ @����:        ��e�'��PAf�w*�������J2CC�z�!m۶M�tZ�x�$�����*�ĉڷo���+s"D)O/��n���T�wX7�^�hpǂ�)��s��KF9�=���zzz�K^s���D"%��%�k߾}���G}TMMM㹹���g%vo �.��C  ʥ�Q�      �3f^f:au��ʥ*��r��%�E�K���x�=��#r:��F��*��r)
����ڳg�.^�X�z���]���2�lA]M��7�4���h����տ����B!uuu���u���x�6?�c��>��G�*
�n���.�KO>�d�7���5��O-H  ���p�% ����     �\*Qw}��T}5���i����\��Գ�lڴi�>�����Q333e��,�ݮH$���1�ݻWgΜ)K�R�>_����_4u��;;QU��1���8�C�����m=��8�N�[�N6��l�].��-[V��a���>���Kr8�z�Vǹi�`P?�p�k���}�  �/6�]�2�'���4���ܩJ  ܪ�7���wn�/t     �5�t������k.3W�D�r5�кu�c�555izzZf���@U��l
�Ê��ڷo��=ZҦ�R�5�g���'��f�^��(ᦘ�����+V/��ՊɃ�k�'
��^��컫'	�?��5P9���:z��"�����qnɪU�488X�/�Nh�O~R��l��+�  �����(��8��R�F���l|� �jm&����_�n�J��      >���ߩ��Q��,�iX�D��+V�Њ+444��'O*
ͻC5P	�PH�a襗^���ז-[n�k�"��s����}�ĖE�)����+���XO����������Z���dRǏ�aT���<R����߯��E"��ܶ|P�p�`<�wP�{�ȂD  �*���VG  ��X�      3��:B���k.��zլ8����SO<�V�^�X,�l��ͺ��A9<xPP*u�[��r��8e���~DM��7d����K����{�|>�U�.�K+W�,k�T*�cǎ)�a%�bf���~�m����
�p$zur:�z��ǋ�Q��/+;=lA*  `�h4�� ����d�       ����gDf���R0���U�w>MMMz�Ǵq�F%���j*J�������7�������<G%��\��`��ZD�;nȈ�������̜��_Нw�Ypm���e=b�0?~���E��ٳڷo�r����Sr---ڴiS�x.ե��  +d�Y���Y �y��n%�I�c      �j�:lO�٬NPL��o���A=���o߮\.�x<nu$�9�׫@ �'Nh߾}���V�T�<�����1���+����׾��>�X�xSS�ZZZ�V�4M�:u�����̌�z�-��a��Ֆ-[t��%MLL\5>�ʷ���gܰâd  �&sjBf�Ι����f����jll,S"  n���]��,�����
ww     �G6���g��w��zas��h���)�r��}�v���cǎirrR�P��X�c.�K�PH.\бcǴv�Zuww_�9�.ʙ��3W��[[=.��4�㺲�1�����҃-q�����֬YS��}}}���)k�G6�ի��*��]�S��v�y�=��so
.�����_G6�Ǣt  Ԟ�W�X�y�ƛ_�i��D p{�^�r�����pNџ��2%     �l��kO���\vO����c%�l6mڴI�t��	�����T�gv�]�HDccc���WWW�֭[7�cK%?�&3�r�K�䌚Ĳ���+;{�GU�.����c�<\0���-��]��/^\Б�G�ի��*��/���V�����;�(O]����ǂD  ����欎  ���^�d     �~��^�#T��Y�����l6[�$�a�=��jjj���tU�8��c����ǵg�>|���R��>o�{�o��{m�_�2b�2s�yC0w�>���`5PCC�:;;�VwffF/^,��(���!�ݻW�a��/�f�l۶M��UG����ΎZ�  T;� ����M<      HO��*�᭿�\vW����t��ܚ+Vh�Ν������ð:�\$�������u�����&K���|',�e_��wg���^�L�|N�C��v�ڂK�V�*�
�J�R:u����h4��{�jxxX�p��8�s�ݺ��
�s��F��Y�  TR2��:  �jll�3      ����fwX����ycwn�(-��+�.]��\�֭S,���Q�B��|>�^y�8p�����7��.���2���Z4���\rVy#S�Z�w��G�R0���R�&�|>�S�N�2n����z��t��	��ᒮ[�V�^��K�����#�Gߵ   ��X,fu  �U�'�     ��lr��V��(��MKa�������p8��{Lw�u�����欎�:������444�����|o��4MSyG�wp��OX��WEQ��Xe
��˞Tkk�U�6�M===e+;00�x<^��Q:'N���/�,��%��mu��Tlw3���w�bA  P)���e;� �������      �*��X�blv��4���|_7��1�����Gս�ޫ\.G,���(�ǣ��Y���X�
2����ۉxC�7�M4����M+���n�sG�^O>��`|�ҥjh(~��횞����HY�F�kϞ=J�R
VǩjmmmZ�bE��ԡ�V���,H  *att�?� U�n����X      U������7%�
����p�ۭ�۷�G������ՑP��|�o����z�H$488�h4�๊��>33#����gy�%hpG�J��nmt�W0x�1D�C���e���f���W��Qsssڻw��D���hl߾]v�5?�MS����5�  @�[ �����     ����7��t[�"ܡv�#Ԍ��o�鶚�l6mڴI�?��533cu$ԙk7���l�z�J��Z��d���\R6WyO}��ip�E4��jf^F|�"�2�|_;�^0���.��<oj�����d�27n�i�:|���z�-��a9�#-*�PHk׮-�=���X�  �[,��*  ����+�N[      ��f�3�au������^*6�G��P�x-�[�n�v�ء��&MOO+��[	u�����l�x<2CCCC�i�ם�Xof4]��c;��$�q#6)3��@���r��q8���*K���QMMM�enܞw�}W/�����^��q��ﾻpwI#��O�  �J�x �J~���o2     `�<M���&���.�cԔb�����ŬX�B;w�TWW�����������u�[�G6�M###�|��/�m~�4��s��k��d�΃��������{��0���@HJ  b@*��M�N�u*�nb{׵)WvSq���J�ɺ,��ql�,�֎dY�#��+ْ)��^ H"������=}_ϳ�v��y���~��T%�����0����>��I9�Ԑ:��O��c�kև��o�	�v��e]�|��}qw���u��q�R)uu��q����٩�۷׬'N��gκ�  8�P(��x ��'���  ������А�Q   ���F��u���Q��mnGh9�����v 5<<�'�|RJ��u�cw#������|>�477w�g�r�n�{�
�u�O���D�;n0Ky����,K��)��ᛖ=�FGG)��{�\.;�7n_�T�/��K�.�����8-e߾}2��E�ҵo�_�  �1MS�D��  ������cJ hW>�O������s;
   �p��{܎�_�O�z`���Z�����7�ǭ���q9rD{��m��?�s�����
ZYY��쬊�b��풔�8�|����w�Pɬ4�N��	=q������!�߭�������L��ǳ,Ko���^}�UE"G����x<�͛7׬���G*.q�  ��w @3��b4�     ��/�ߚM����v���?e�1}n�&�����z�GT�V��fݎ��N�?��z�J����P�1�*�qghp��lc�c�f�Rggg���Ȉ�,���Ԕ����]�|Y�>���ժ"���qZ����_�fU+Z<�[.�  NZXX�=�  �|>~�     ���W�}��������-)4���z�6�������z�������J�܎�*�۲���Q�R�{-��-5�cɠ��
IR���Y)9^�8���쫽����O�p��z����ⲵ�5=��3ZYYQWW��q���Ȉz{{k֗��O2K�{  ���������: @�`z;      >�7ҥ@��c������v��������'iN�ah�޽:z��B��VWWݎ���۾S5J���S�4��V��tt��NH����|s�[~M���5룣���*�˚���}_ܚJ��'N�ܹs���b�h��w�}5k�̪V_�#�   ���ͩ\.� �b��
���1      ��B#��Eݎa����2��N'ng���ܯ]���$����ӓO>���^%	���v$49�ǣX,f�~�b�f-�L��eo���hpoU4�C�LU�	�˘���ԮG�Quvv�^����_��8��7�ԋ/��p8,���v���c��������B  ��\.Ǆ
 @S��b�f�n�      @3<>E�엱�O���)г��-��9(o������mٲEǎ��ؘR��sXWgg��^�m�՛ྒ-K��6;1��um�W	�E%��eV�/4���>P;Uzxx��R�|^�7;;��Ǐ�Z�*m�;m7*�ϧ;vԬ箼�̻/��  8�P(hyy��  ���T�6�}&      lh�pL�$��$w��+��~�c�>ø�u�4����!=zTJ��u����zzzl۫R���l`)g[�u1��u��UsɆԹ�7'�G��z���﷽�իWeY�����t:�g�yFsss���v;����D���g��'  N)
Z\\�al�w -�w      ܪ@ϘBC�{��'QǶ2<�M>��"�{k�r�������mt�x\G��޽{��f���ݎ�&100`�^�b���B�g[��0��u����,K����e�so���լ�z̅t���⢭{�>˲t��I���[��ꪹ�����Wooo�z��"�Ԁ��  ��,�ҕ+Whp 4�p8�P(��      ܲ��=
��5+O ��G��܎�6�5�K����E":tHP�ZU&�q;\f�`��NX����X�[ݨm�,feU+��^{K�x�f}hh��ZW�\�}O�z���������*�D�ڹsg�Z��V��?s!  p¥K�hp 4���.��     p�£�*<�[j�;����;?#O �v���L�����8�C����)�J�	.����m�z�M�T�c�m5�c���U����*��bV�����H$�h��;t������m�7[^^����U(��܎�O�}���o+'~߅4  �	KKKJ��n�  @�x��m     pG����+y�����������7�/�_A�;�ah�޽:z��:::hto3����Q��ྰ��:�mp�����ZVs�"@�Ts�c�\}C{v�S�>00`{������u�|^�=���������vܢH$���������S95�B"  `�l6���E�c  ���.�     pǂ=c��<(O���(2���VEw<*��w;M[�;��f����o|��k�.=zT���J$2M��Hp��Аm{Y��B�P�>��o>�D��F�{��E���'�m*��@�����~[��e{`��^�u�:uJ�XL^���H�M۷o�Y������   �e�Y����  uuu�R��      �7ܩخ�����T^O�C��)<z�]�8X�����gd6۲e��;���1�R)��ma###��U*���q����z<A�[��� pO%߀cE*%��c�,wvv*��	�ڵk�=f�w�yG������T$�7��j�֭z饗dY7�[\}�5���R*  `�J����Y=��ü �&�(� 6��Ҽ����w;�+~y6�\�}�ZXXp;   ��O��=
��+7sV�\���=^��Q���a~l3�������5����y�����!)�H�̙3
�u�bc�F����m��Nv�V���z����hpocf~����i��Ў����>{�X��]�f��lyyY?�����e�73�#�h``��Ñ̥WT^[��s��d  �.���<M�  �twwKR��� ��f�*�y���8yiI�*?C   ���Wl�*�e�]T5�p����)�7�������p{�;k'�K4�;���[G�Q>��o�!I��E��9�]�������WN�"�	�� 7���ƪŬ�56U���׬����ZgeeE�R��=�Q�\�ɓ'��z����v�h��͵�,S���V���N(  `�˗/+��19 �����E�c      ��b}���Tɬ���Q9qMV�l���t�߳I��^�=��V��-
􎩴2}�����R������|F�RIo�������Ѩ۱p�FGGm�/��լM�'��豵�G^?��-�3TڔY�ɪV�����鼣���;����mݯ�9sF���B���~��[��x�&��x��kp  ��L&ÉF  W����}      ��/ڣ��u=��(8�M�p�������w+<��:�=����(ط�F�&��������R)Ҵ�@ ��СC�x<J&�nG�m
�m�J�Rw0�L�����`��p��T��q�Fe�=ݻcSͺ��ۋ�"�,���˗555�x<�H�'�V��ӣX,�t:}���[O�,��	�w �F��d4==��[��4M��  ڌ��W4����Q      ��|��u\��i�,�T-�e�
�̊,�"Y��W�����	v\��/�n~ܑ���i���|ӚeY:w�{�1�R�'�0�o�>I�ŋ533�x<�r*܊��1y�^��[o�͂Ǿ&�����.&��)��}�w�Nj������yY�e��`mmM�<�VVVx��&�/c��Z;�}�   ;�r9]�|Y��EEu    IDAT�( �===2C�j��(      hG�<����a�*4t��#��W��	��+�3&_G��X��S�q�o���i����	MNN���G�d�>�&�y�f[�����/����jk�z����5�.��T����ݥ-��>�OѨ�O,KKK����*��N�8�s�Ω���&�6222Rw}���N  �p���� \��ݭj��       �+2�@���o��gdM`�֭�����ؘR��*��ۑ��`PCC�NV�f�5kg��[�|�a�hpou4��!�\�Uu��U�i�Hg�z<���:��(��۶_�;{��N�8�p8,���v4�z����56  p���܎ hC����?      �q]{�z�Z.������0�kppPG��Ν;����R��v$��-[��㱯e�T*�����	�Vc=F ,��u���s; �,d��[�����5���ݶ�az�����Յ����܎�D"uuu)�Jݴ��~K���|�>���Y�*����5�Ŭ���T)ʬVd�U������I����������<{o4 4���5���hpp�	� ����|���J$nG      ����5]��j��|�Mm۶ͅDXOww��x�	��y����,K���S���o�n�~�Lm�i�Z���:�xC�@��ېYr~�VeARm�{<��������t:��'O*���g��idd���]��������r'n�U)���S9��jfU���I�$��બ-޸fx��E����?>,��i �*2���^��O}�S�V�n� ����>��r��v       -.��3�ut���y��믿���ɟt)>N8���U.�u��i�r9�����W===���fk֮,$U�}��:�����;o �Y�9^c4P{wN P(��F6�U�P�m�VbY�N�<��������z9�׍���]_;�\c���U2��^~M��Ǖ�>�����6��ZU9�����z�{�^>�jf���  ����.�z�  ����O�eqz       �^����V���򲦧�]H�[���u��>|X>��v@'�c�[��V�u�/eö�Y�'mH��	�m��	�V���}�OT�����Y]]�u�Vq��y��ϫ����v�X��=}����'*�T�W�\ҹ"��rr^��|���?V{� `㘛�S"�P4�� �����W�P��      @C�<�w����Ԭ���s!n�aڻw�$��ŋ���Q<w9Uk���ڲe��{f2���\�l��N=�`D����v�h�6c���̪�5����Y���Y���:~��r����h�p�����9��ړ�xf1��{�*;�����Qɬ*{�z�F�� p��ښ�{�=�� "
�����       4L�}����w��)ql0���TOO���L�t;RK��{���m�smm�f�ʵ%e:6�Z�o���vA�C��6�i��Z�a5�v6]W*��i��������}�YMMM�����8hr+++ڶm[��T�ʛ��Y�
��i��s��-���ZP���*-�/� l8�t�w @�H�J���I       ���S�C�f}qqQ�/_v!��֭[u��1���+�J�R���e����	[�4MS�l�f��U�T�o�n�p��5��zh3����ﭝ��x�Fm��L&���;�4����ԩS����˱X�7�<��S����>&��덌�aU��^~M�����ݨ�YUn欲U)� pJ��Ν;�j��S�  ��7�[��T       ���߭���+�48	�488��G�j׮]J��W���-[���a��t��w�4MM�v�Z���'h��͋�6c�����~��D�Nu�S�Tʶ�6���{O�>������z�Ţ��>��Ok�����͛���L���Ŭ�_P9��v�����P��;  �YZZ������� �(�׫��~�r�S       ��yߤ��5믽�ӿ[@WW��9�|P�|����aڽ{���&�ɚ���5bc���(o��!S��hpo3f����V��M�����hmm���6���?~\�DB�x��8hb�e)�Hh���:r����k###���5�Mn�T##BR%�R���r�Ɲ2Ye.�P5מϻ �%	����x�q ����^y�^
ξ�       5����k�s���|�M�	�pXԣ�>�J��t:�v�ettT===��Y.���pp>ט^Fo��!u��xh'�%��������}��Fk���T�ZU6��m���T*�ĉz�w����4N|�D"���n;vL���5׽^�FGGk���4u�u���Rʾ���J��(�Ȫ�����B��( �[�J�hp 8nppP���      �}���d�~���ϻ�N���z�Gt��!�|>�R)�#5=�0�g����7��P*�jp��>�0yÝ��A�㡍Xղ,�r�F��\w��	��t���G39}��^y���ᛦp���T�V599��۷�c�5�[fU�k�8?�,�y�,s�4�Xղҗ^�& � L����T�7  ������L�t;
      �6�ߢ��&k��y���͹�N�x<ڻw��=�h4�D"�v��566f��v˲�~�ƕ5U1[k��	�dx���A����4bJp������pضkkk���̦��u��q��i�h=�JE�dR?��8pK������ipw�U-+��+�6�����ʅ�j̯� �	������� pDWW�B������Q       ���'~���~��'A�MLL�رc���S"�`ˏpjz{:��{��yk��Z��"��A�ۡ�X�4�j���^���ǳ٬m{5���5=��3ZXXPww��q��VVV�e�MNN�֍$���uי����[2�w
�Y�(���1  � �H�ҥK�z�� `���IR�Tr9	      �vֽ�o��5X����/�P�?��e���:v���ǕL&�6`��;v(��|uu�f��|R��	�k}�a�v�K�nhpo#����]������R�6�����_~YgϞUWW�-M�F�J�R����SO=�����d�w&�;����J��V)1����1  #������L*  8bhhH�e�A       W����G5�BA/��������AMNNj׮]J��*��lF~�ߑ��B�g��R���N^��u�\hpo#�Op�L�t�k�#��m%��jK��[o���W P0t;�X>�W�\�O<�]�v��>�����k��2��9V�����c�&?��
���-..�ҥK�x�� `���.utt(��˲,��       hs���<�����Ǐ3��uuu�ȑ#ڷo����r��ۑ��} �$���Ԭ�s�t�g{�z��ކ�As�ӡ�X7"VӋ��="
�V�վ��������*�J���t;��i�J�Rڷo�}�ѻ��o���k��޽�}����۲���U-�T�> ��D"�s������ �BFFF$�%       �x|��~��׬'�I�:uʅDh�pX�c�=�j��t:�v$��b1MLLؾo�T����򬥪��a���+_���:h>4���t��2T\��<l��*��|^�=��fff�6?juuUCCC:z��::j�8�S���w�U2�2��j�J6�rr���+�L��_s; `�dR�ϟg2 �V��Ò�r��r       �n����Q�
���Ose���|:p��:$�׫d2�v$�8p���g���5����	첽V=�H��o�>��ۈӓ���?�+��.�Bac7�Z���'O�7�P,c�&>V*����דO>���1����驻^N^��V�k������� X�i�Z\\ԥK�x�	 �EWW�"����"
      h��	���x����N�>�B"4�ǣ|P����F�-��m۶j�T*���V;��+9U�}�׫����@�{��,Yf���b�uܯ�t钞}�Yy�^�B!�㠉�J%��y>|X{��q�N�	��v���T^[t;�c��9����1  �XZZҹs���� ��mڴIR뜰      �u����J2���o}�[��M&&&499���~%	���v����C9�w����JUC{��Q_@�P�!��|�rhV��c�ê��l�Q,֯�����}O�TJ]]]n�A3MS���ڽ{�<������ip�Wi����?'Y�TZ��v �:VWWu��y����<  hm�ahddD���      ��tlݯ���Y����믿�B"4���q;vL���J�R�T*nG�#���wd�n�PP*��Y?5[T1�o{�z|�����D�{��L�|�����糭�F��^(��/hjjJ===n�A�K$����g?�Y���Ԍ����F���,S���)WL̊���9�����%���< hm
�*�~�      ��4���M�)�����y_��ѣG�k�.���5�wllL۶msd���Ś�r����]���(�0��5���mª:��6jk�|>u^4ܩ�2!�̙3z���D���ݎ�&��dT�Tt��1mٲ�����h��rj��9ZY9� ���s�rA�̲�1  �XZZ��o�M�; �lڴI����\N       �E�<�����Y�v�^|�Ea#���ґ#G�o�>����?<���Gud�L&�l6[���Ԛ��LU�v����7\�m����^;��W*YM>"xjjJ����U�T�D܎�&V*��N���c��Gq%�zܫ�t����rz��SY��k ���.^��b�h�ͧ �����400 i�       ОF�_ם��g�g*
��'����z��T�V�N7_/�az�Gm�۲�����Œ�챽�z���i�G���]�U�KDC����lp/��w
r"���O?���U��q�㠉Y��d2���	9rD�@��,�Mp���E�FUY[q;B�T�Lp�fe�����t��E�� ���証^���"��      hj�-�����Ԭ��i=���.$�F���t��:tH>�O�T��H7�ڵK����콺��b�X������D��Q�`D�`GCj�y���&,9?��#TۨkgM�����U�Tt��	]�pA���L���J$������zzz܎��|&�0���ڣzZU5��Um�� ��---��7ߤ� pG���%��q�       �l6�w_�'�Y�����D"�B"ld�G{���ѣG�F�L&]���ק|Б��岖�k�\�ez�c�#5��w6��͍�va9���3����K��&��={V/����ᰫS������J���=��;w����[�ɭ�����w���j!�v �:�ɤ������d�kt @������$�J%��       �'�l�Џ����R��?��?q!Z��Ą&''5<<�T*�j�����PH�vl����|ݓ\������Q��/_GwCj�����.,珏���d�i���gvvV����U,���1X_�R���z�!=��cM�LVo�{����Qͷ_�w��~�g �(L����
S� ����\NV(       �����M�ޱ���_]gϞu!Z��Ȉ�=�;v(�˩R�8^�0=���
�Î�N������\^H�J�>Gj�������C��U�.�� �Z��c�,���[�ΠFJ��z�g477�x<�j4���m޼YO>��"��#��E���Rޅ$��,fݎ�p&�������̙3�,K�Q�� ����|�t�t2       �(<��F��Խ��o|C�r���Њzzz�������W>�w���~X�����]�V5??_�n���Y�e���Q��+_��!���hpo��mp��j�FY;gܚf��^|�E���[���j�)�hkkk�D"zꩧ444�v�O��5��G;��%�#4�U�? hfkkkZ^^�ŋ�� �%�6m���i�*���g       [��S��O׬/..�����Ъ:::t��A=������u'�ߍ]�vibb��=���|�)�����L���~��s@��ϲq��������M2n4�������~�P(�`0����8>�����ڽ{��qn�[�c�U�#4���qK ������7�x�w �-�$�߈      ��0<���+�W�����r����B��<�C����imm������mHW_:���3�/�����~�ax��hX=4?�ۆ���!ǛdLǛ�?477��Ǐ�P((�5�.6�4�J��������n��wwNKh5V�����6�=�F������)%��� �X������$
��       ��	�������u�4���}M�j0����޽{u��utt(�N��>===:t�cCL�岮]�V����}*�z�[���_��װzh~t4��<��1u�n��y=��s���Qww��q��VWW544��G�*��ͦ��s"  4�r����e�>}Z>o  ַm�6IR�X�       ������]�>33��|�;.$B�0C�v�ґ#G�ǕH$n��2��'�p�s]˲477W�3�sW��~�Îԭ�0<�w6�6�ۆ�M��%�?�tr¤i�z��W���+�9>�[&����דO>���1�����cxگi���ݎ  ����:s�,�b�; ����\?4�ɸ�       ��j�?�R�a����w4==�B*���۷�رc������[F"MNN*;�gyyY�\�f=�/���d4�d_׀/}G�����&VC�����T#�K���s����9�_�TR&��g>��ٳ��8�(��5k�ؘ�v<2���  ��ɤ���t��En� Եe���j��R��v       �k�݇5p��Y�T*�򗿬B��B*����1=��Sڱc���lM�V(��䤢Ѩc�٬����^�J][��Q��+'��Q��6a8}7�ׯR�FY;����ྼ���Ǐ+�J����ֽ�ZL���ʊv�ޭÇ;v��5�{Cν8j'�?�v��3�$ ��^z�%y<Nt �����8�,�ͺ�       �3�����Y_\\�������G�Ҟ={�����%I�����3V*���սv~&��Îծ�n�A��d4����VC�:_Nv6�{<�|��J%����t钺��m��+�H���_O=�����qlWo��w[xCnGh8o��~� �Q-,,hvvV333Lq �d||�ƍ���       ���i�/~M�/Ps��_�k���B*��H$���GQ�Z����u��GjY����YU*��k�\A?��/9=L�Gx|�;�V��SM�����vL�>s�^y�E"��~R�U��iU�UMNNj˖-n�qL�	���m�	�ߍ��{���T*iyyY/��2� �<��m�&�zs�i�.'       {E����O��׾����ڵk���߯�СC:s挮\�b{����r��׾}%�Bx�����=�Іzl,|e��<	��|��,�SSS�����J����w��r��L&�O��:p�����r�\�Y�K��-��ζzfx�m9� 6���]�xQ+++��L
 ��6mڤP($I�f�.�       g���خC5�BA_�җT(\H\g���٣r��J��R�d˾�DB�D���ޞ�B�l�s�<��|ў�����>�wmΐ�M��B�$�zӡ�ԝL\_[[�3�<���U��q۲��X����Um߾]�V P{Q�Y�Y�	��0<^�:��y��i��~ h�LF�dR'O�d�; @�ah��풮��a�{:       �L�W���Ǉk�-,,�_��,�r!�r����+�X,���e&����B�kWV����w��z�^�h����D�\�vZ{�R����4�W*�8qB�ΝSWWWKO���K�R��bz��'����v��Y����mp������a|����@+���ՙ3g���ir�67<<|�ԻL&�r       p��kH���ʨ�Ww��i?~܅T�����t��e�b1���*��P(�VOf�X���l���P,黙{d;���|�yC�����C�{�����n�j���J�b��^����Ϟ=�'N(���w%�A    IDAT��|>�R��#G�hbb��8�^�{��Sqg��!�#4L��}~� �JVWW�J���k��� mnǎ�$�4U,]N       ΋�>�ѿ�+u�}��ԙ3g��5;;���%IRGG�6mڤ��N��e�����m�R���t�Ǚ��?{ߧ|l���ex�
�ljhMlL4��	�Ӏw+Pw��#�����fggu��q�E�b�݃�U*���i���z�����S��]4*���7���G��nyBn�  �˲477�S�N�Z��� mjhhH��ק������       g��Y��vͺeY���������|Ļﾫ\.w���`P������Q�R�;��4MMOO�ۿ��I�wʱ���w���2���=�:ې�q�Q�h�ꮗJ%�j�kpO��:~��������m[-��d2�͛7�'�P8v;����d�u&������w��� 6���%	���[����1 �|v��y��
�       @������*<���R�Tҗ��%%	��V�:w��M�>�OCCC�eY7��-���������޼.tq:vO ,���u�1���&��*E�~����Z�B6�[���'O�?������v
7nM*�R ��䤆��P.I���u��q�|���ܐ�`�>�=�n�  ��4u��5�8qB�i2� �����M��-�r9       4�7ܩ{~�/�����L&����iz6��|>��/ֽ��x��߯��!Y����ye2����YJ���%���6K���ؘ�n�G���_wƪ?����_4��;wN�?���^�MM��G�E��y>|X<���q�JݻK�������O���n�pLp`�O�6�@��v�VVV��o2� ڈa��{$]$�4       �U�����ߖ'��633�/~�z���ʊfffֽn��٬��d���\A��Gf�۩���w���hx]l\4���'g=Ѻ�v6���e?~\�|^�X̶}�zL������~<x�I�uԛ���$Å��Z]p`[K6����}[܎ �A�\��⢞�yU*^;@������l���       �Z�և��O�3HvjjJ_�җT�T\H|������J�z������^+���/s}*Dǜ�W����{��u�����F�nZ�{U5k?��εj����9��euw7��!l,�dR���z��'o|P�Z��CC�����y|A��w��v��ݎ�< h���i�������Lq�6`�v������      ��}�ok������Ο?����ߓi�N��5}�����r�J��W�U��O�ΉFī��"�Ð5��ۈ�:��ex���֬���;�Ӳ������%uww�0�����N�%I���w9Ms+�u��	�p!M{�o�7�:7\x#]
�nr; �F�bQ:q�S�����)�~_6�U�Z��       ������?�{��ɓ��W�J�;\U�Tt���'����jjj��c-�ҟ���B�Í�x��s@�P̕���hpo#�/�x��b��R�tGG�����ڵk�tc����U,ƓnV,�J�t��A�߿��8���bݣ���Ð"��dx6��^��Ud�>I�p ���իJ�R:u�S���y�^ML|8�%�ɸ�       �����u���^{��W�����4��U�tZSSS���Y��]��s.�١'��CH��QWjc���]v�e���%)Q��]��c���fggU,�6�www�q>��4����ݻw��ѣ4a݆�����4�;��)4z��1�Zxl�����1  (�J���׋/��R���+ hQ۷oW0x�}�l6ˇ0       �Q��-��K�y�g�^>u����/����?��u�?�^Z��k`���`�ɠMw���6҈	����5n���4M���kmmM�`P�Q2p<���h�dR}}}zꩧ���������q���
����pg% ����i��i���k�z��. lL�`P۶m���l6�b       hb�G�~���'�^~��W��/Y�J�����,��7��M}�[��׿�u]�z��1�]Xљ�!�]���'��Z}l|4����Lp��O���K������ ��'���,����86�L&�j���G�j�֭n�ٰ���k�<��B�4�7Bx|��]CnǸm���B��� �r��k׮饗^R�P`�; ���;w�xn��gl       @}�ׯ��������^?}��~�7~C�B���ЮL�������駟�t������߾�G��K	��>&˥���`��Wj�u���F_���k�aI�52�L��g2���J��~�-����c�d�T*J&�:p��8���]����#�K[#�ٲO�����2�O[��z �fff��f��/���|�M� ��!�i||�Ư��       �����g���Oս��;������t:��dh7�bQ_����/޴�����|�+�,K/��ԩ��K��ק��6�d��E�B;1���%
FH��U���ddY���e���)��+����>�O==�)woyyY[�n������q6�B������������}��;�?>�v�O��c��^� �\.kvvV����VWW�� -��{�q���ښL�t9       l�/������^�r�>����ڵk����L&�k��k:w�\��o����������o��}(ؿ��>U�:�ڌ��|s�\����4M�r9Y�������*������w@*�R4�g?�Y��e\�z��N>ټυ4m��Qd�C
�mv;I}�ئ���in�64;;�b���Ǐ�0y��	 �{���7�O��}       ��3<^m������~�����e}���ٳg��nzzZ_��t�ʕu3��\է�Oy"�&�Y >,o�ӵ�h-t��O����R��������������[[>�W�Rё#G411�v��������`��c�c��2��3������£�J��  hG�JE��Ӻx�._��w ���^�v��}��kkkuo|       |�������~��ֽ\(�[��[z���ԩS��������0m��_զ���d
�o�ǅ	��pL��p��u���f�4��Wcu�3���~�-5��������j*����z�!=��#�;�ҥK5k�/���]H���C��|\�h��Q��+����#nG �lnnN�|^��)�4ir�j���D"������]N       �ah�g�om�����0�j�������?�U*������_��~�w~G�r��c_@������O��׼>��07������&5�&Zݣm�ܗ�u���٬m5�~����l��K&�ױc�n|�gLMMլul{Xȅ4�Q�P��;U��}2�����Աu��;���/  ��4MMMMiiiI�O����m�! ���D�}���^[[s1       ���#?�{����{�?�����/hee��ɰѥ�i��o�����{"�/ڣ���z�l�5O�C��1�cJ�ã����7{ w��6��e������sf�z�\^�N�;1::j�^pO2������䤆�9��i���u�b���u��=��oR���t��O ����y�Q�
 �X]]U"��3�<�|>�w �`x�y�^IR�XT�Xt9       ������yB�����W�^կ���N���w�ѿ���V�ϟ_�1������^Rl��=_��~���ND�I�o�<�������nCF��)�ә�M/�\ζ###���+�*
:r�����v��q�ҥ��]�78	>��Q�g�:wQ����w�{���#|H�V�ޣ
�o��
 �qMMM)���^����(	 hn�������k��      ���ch��zI[�{=�N�?����?��?U�Zmp:l�i�����~��]�Tj���vѽ�ǫ
O|���qG�k�G��8�?���ڐ7�Y��Ѽ�y�G�R�z.�SWW�-5����ŔN�m��a���ɤ8`��n]��A�W���������?>,�RRemI���*�eUK����萯�W�h����2�~�B ZM.�ӵk�t��)�߿_���2Ms���  ���|ڽ{��_g2U*      @�
�l��yB����i�/��eY��w�������~��488�BJ4���}�+_ѻﾻ��C�O����޿���ã��v���˪�����[����{?��6�	vH�eGk,F%cE�ֳ̛٬�u6oެ�g�ں'��L&�c�}�S�r;J[�,���5����f��������gT�dU+2�Y����JQ�Y�̪dI�zex|2�!y���2�� �W�\Q�����\�������T.�ݎ Xǽ�ޫP��)~�i*�ɸ�       Z��j�gC[����e�j��^�rE��+�����֧?�i��BR4��^zI���7T(�}�7Ӗ_�]�<�wn{�P����l`�	F��b�^�zhpoC�P����W��G݁�������~{������d2E�QMNN�������=����c.���O�H7(  �R���ի���:s����+��#�4?�? 4TOO����o�:�Jq�       4H���Ux����?������bQ_������/�s���\H	�%�I����Μ9�Oh�?����Z�p���a�sw��<��B��H���>_am����:o�{���\�iw���G]]4v6�R��t:���w��q����?g��A�$@Tv��5�(�P���N|�I6�o|oֱo6�����f��}�M�$N�Ď7��Rl�H�X��H�)KT�D���	�`ш�3��s�!A3`����~==��3���"A`�s�G�7oֺu뜎3�?~<�zŚ�8	  ������F�c�������U @�U�VM|�H$�;�       �{%mwk������8�9]]]��?�#���K)�Cl��[o����?����u|Zw�ѻwTn��S9O�;�i�5,*H���>G���Oq�h�˺�Fs�OkkkN�wζm-]�T<���^�ӑ �ȑ#kn��7;�  �D�m�̙3��bڱc�$���� �N�,Y"����}FF��@        �+��Z?�=u����.��zN"�г�>�����POOO���.]��?��?דO>y��4fI�:>������*�]��[�.��w[�5\��ɸ��������/zS0d�E�H$�W�-\�P�a���pg���UQQ�GyDUUٿ1C�E"�={6c�b����  ܒp8���~?~\�O��i�r��� ����*���O|�D�J�L       ���K��O�l釦<�̙3��?�c}���� Y8ollLO?�����/d�p�_��mZ�ţ����9�a�L��;e����a�T԰P.oq�3S��0G��Ҽ�Hۺ53������s�OII����>-�366�t:��~X�-r:>�СC�,+c�b�GH  f�s��)�k�����Lq�i�4M�Y�fb@:�V$q8       @����Z��_S�/��w�	ضm�?�����@�w���Y8ò,��������}���Y�[׸��j���ZK��K�V5�-��[,om�M�o�|����9��+��pn��Xy��\���p�>n^*�R(Һu�q�F��OS�X3L�*V>�@  0ӥ�i�9sF�HD����à� [�d�JK�h
�x�       ��ej���w���Q��xx���᰾��o����o߾&D.�8qB�'�'�xB����=�b����ώ�~ۿ�
пs���)���y�a�[�.�8{�'s�a�U�Wz<��m.X�d�2������Q����l���f�t2<n,h͚59��܋�b:q�D�z�][��W;�  ���������l�2���˲��N  �GMM����'>W2�t0       `*���Z�_whh������R�CY�����?��?h�ҥ��'>��֛���;wN�>�����nx���AͿ�%�n�T�M�^ +1�t,��b�0�m�����ɀ���>��%y�c4e�b��XO$��b9���ri���9{>\��ȈJKK��#�Pn���ߟ��P}ϯ9�  �&gϞU2�ԏ�c�R)y<�� ��x�f͚����m+3�       �3�P�OişU��_��'O����}��_�������ܹs����}�_�q��p��Ok��;Rn������C���r��1���ILp����J�R��9�Qki_�z8VQQQ��Y�x��;�T*����d�&�?��r��>f�سgOƚ�S�����@  0�$	uww��v��_և?�a��n�@�\�R����B!�       3���A������.����H�O�<�ĉ:q�V�\��|�#���	�>}Z/���N�8qS�vnR�����/ڜ�d7f��w(�zbpεr�YR�p:�u��0���㓕��u�F��J���GGGs:���󩣣C�O���s�*˲4::�M�6�����8��P(�߉�5?W��8  �ٯ��_uuuڷo�-Z���4M��i�����`�͟?������1       P��?�e��K��<������W�Oy�#Gt��-]�T[�n�ʕ+��r�Y�������_���ޚj��?V�.M��_�"�<UMJ��K���^�
�s�Y\!+9��=ƒ�.�����k"������)cwjٲe����6�9�r�J͛7��(�{���:���g~Ł4  `�:s���n=�������-���ʲ,�/�<*--�]w�5�m�q0       ����7��*����_���~�%Y�Ȕ��<yR'O�TCC�z�!m޼Y>�����h4�ݻw���_W ��Ǹ�՚�����G>/�3=��x*d%��.��YT�t@�9�,.W2�߂�$�թ՛�&���HN�eeejiiхr��sU$Qee�y�����ڵ+c�]Z�ʻ?�@  0[������[.���?�_��_���Q"�p: �J.�Kk׮����K{�P��       `pyK4�㿧���V/���_*=�������?����ymܸQ[�lт
�x�;{��v�ܩ}��)�L��c̢2�o�m����YR��w�W��t`
�s�Y\&�pɶ3'<���d��"y��S�GFFT__/�˕��V�^��/��mJ$J$��{��x���;p��i���e��l�u�����  @����TUU%Iz��w�~�z��n�R)����|�rUT�w{���q�b��<       0Ӹ�j��?Pöw����W���N�cccz�7��o���U[�lцr:�v.	�Bڻw�v�ޭ��ޛ~��ȯ�m�S�G��ܥUyL�n��:�%��B�h0��$Җ��k]��7[-�����7e�Tyy����u�ܹ�=�\`Y����6nܨ����nl�ΝY���L��  �����Keeeڱc�ZZZT__/˲dY��� �y�橭�m��t:������        �l�/����e���u��t��]�pAO=��V�X�6hժU�z�J=3�������ڳg�N�:uKCv=���U������cJ`n����Uy/�K�I�k�;*;���>22�ӂ�$�\�R�ϟ�Hs�����x�bmذ��(ȑH$�d���lQq�
 �� �L����Z�b��{�9}�ӟ���Q"��K ����Z�z���P(��X       ��e�j������?����U�����cR��<�����iժUZ�f���.&���p8<�{t�ԩ[�CuQ�"�o�����\^~O�\���K*�p���t^�7��/U�1���F�����r�WYY�:;;��Օ�眍FGGURR�m۶99��of�f����:�  �%�`P�/_�$���kڶm�D� p�\.�֮]+�����FGG��
       s��ȯ��>��S��/h����W�C���ڻw����+�4�h�"�Z�J+V�PCCC��;ϲ,uww����:~�����o}���R��mj�������J�����F���YR�Td8�[�5��8sZ|0TcccN�Z�z�.\���Y$	E�­    IDAT��q�s�=�vfJ�Rz�72���Um���  s����UYY�={����M�-���Q2�t: �X+W��t�d2�H$�`"       ���*���*����{��ʛ_����dx��M��:y�N�<���~Z���Z�d�į���|�aY�.]��3gΨ��K'O�����m=���Y�����o�k�mP �Pp�$�]ZU����h��+-S�5:i}ddDuuu2M3g{i�ʕڷo_Ξs��m[�`Pk֬Q]]��q�'{��Q8�X����  (˲t��I�Y�F�>��>��O���V�i*�� `6jkkӂ&>�m[���       037ߥ�O~E~�9���v~S���e�on U(Ҟ={�g�IRyy������ޮ��v������$��BNض�@ ��/�ҥK���ֹs���o�9�W��N���*V��W�:� �F��$��B�˔m�l��l������w˲
�TSS����,Y�����e߹&���M�ׯw:
�ȶm���+�.O��}΁D  �f�LS�a���鈴��1�?^���z����OZ>�O�m˲,����Q]]��˗OZ�|-       d0L�*���*���R�+
����}ENﺥn`8��Çu��ት��J͟?�W}}�jkkUYY)�0���Lɲ,ippP���P__�zzzn{:��n��W<�ꍿ����YR��� nw\e2K*���թt��xG�JL����𰪫�s�����Һu������9g���q����zH.���8ȳC����7c��O�S��@"  p3\����2���Ϊ�{oo�***$I۷o�'>�	y<%�Y�y@�kݺu�~��F�w4i       07�����������*��y�>����d���|�PH�PHǏ���ۭ����Ԩ��\~�_*++SII�|>���������xT\\����x\�tZ�x\�TJ���D"�F��F��D"
�
�BV8�� ��Xe�T��_T序�]Z���pk(�c���� ����C�
�]4���J�
�TU�������֦�����y��T*�p8�-[�d�� ��/���hj���X�0  ��x��YYr?}�����u��1555iӦM%w �Ԯ]����&���FFF
>	       0�y��U��gT��g��ȡk���
}E���;z�T*����(m�5.R���b��U��~����邂;&���ry�e%��7r4լ�����%�@ ��[��_�^}}}sf�Y ЪU�����t��Çu���ʵ?����H  n�l,���i�<yRk֬�+���y�橥�En�[�T��x 0m�^�Z�����Զm�B!��       �;b�T�z�z�H�b�]
}E�c�h�ě��_}��o���/H��N�#�wL���(1ܓ�}��R:VT�����d2����Io��BQQ�֭[�ݻw��y��P(���z=��#NG��oߞ�h������a  �m��%���1�>}Z˖-�3�<��|�3*++�m�J��N��ig���jjj��6<<��L       @�5.RQ�"�?�o%]-�GϾ��w=���.���9��֙%*Y�J%mk�_|�ʖl��r�ӱ �$
���Q2�+۶�׻c�: #5����!UTT�|"YGG�.\��˗/��y����S�|�A�\.���	����3֫�}\��  ܒ-Ɉ��E��RI���>44���577�g�ѧ>�)��W$��	 �?�/^<imddD�D¡D       ���Z���OJ��tR�=��=����4�{R����N:�V2���a�J�Tq�j��������h � wLb�n���JE��W0f��X�Vx�&�'�I���&�{n޼Y?�я�ͼ+ʲ�,K�PH�6mRyy��q�˲����g0\���?(x  p�����|嬾\�9�K��ϟWi����^��>�1��nٶ-���E� 0�UWWk͚5�����'.l       ��ӣ��5*i�����N*1tQ��e%��Q2ث���J��(5Rz,$+q�s�[n���u���S� wY�<�ֶ�Wߡ��N���r���F(�#���� wI�o���1ٱ�I�@@���2M3���{��믿>�KB���Z�t�6l��t8l�Ν����X���WUҲʁD  �v\+��Em��R���Wr�m[�N���w߭����J[�l���Q"���# ܮ���_�~ҝ�R��FFF��       �v�#_C�|�7<�N%�ɊE&���J�"2��2L�̒
.SfIe�b�!\7>s�YT&��� {��S:4V���N������hѢ�<w!��a��nm۶M,p:�ǵ}���u�ej��ρD  �N�mK�3tNv��v����p0Y�$�I;vL�tZo��9"I�x<��s�[��z�q�Fy�މ5۶(�       f<�핧�^���I���-Qi�:�["_}����� $Qp�<�ko�N�⪌���a����n�:UUe�9�%	E"�w�}Z�z��q0Ml߾]�p8c���GE�8�  ܩ�Pr�F�:s�l���Cuww�0y<��@���nmڴI~��z �eY�         �C�Y�K��r{o|bDbI�m�X�m[���y��4M�����|yy�\�,K�@@K�.����/���t$L���z��W3�ݥUj�W�@"  �+s��>88�.(�N�g�Q ��`�q�\Z�n�***&��A%�I�R         ΢���C��mw T���yk�����өs���k˖-Ӻ U[[�Gyd�M�G�=��SJ�R�����]V�@"  �Ks��~��E(��;����Ѩ\.u�3V�Z���ɯ�D�Q�b1�         Σ��)���d��#��l�=�&�̜�800�t:��}�͛�U�V���D$�az������tLC�ѣG3֋���~�o9�  ��\(�wuu)
)
����R��LӤ�`ֻ뮻���<im||<o�         3wL�p��}f��%5d��R)�m�+V���#o�+R��FGG�y�f�]���8�������SOe=���_�z�  ��f{�ݶm�8qB�hT���z��d�6%w ��ҥK3.hO$��         Qp�x*
V��%�,�Q\�q,
)�d>(�ЦM�T__���Y���joo�< ���hLo����3֫6�+U�zԁD   �&J�c���J�t��Q��q�8qB?�я$I�i�4M��@n-Z�H.���N�eY�C�     �l`��NG    r��;��p{���l�+�	�36?뱾�>����k����~�������gddD~�_۶ms�d����ɓڽ{wƺYR��O�/ �B�ۖ~���-�'	?~\�tZ��/�,Ir�ݔ��mmmZ�dɤ5˲444D�     ��+��3��OH   ��{�y��+�m�ֽ�R-n�UEjh�z*�R��������C=��^zI���y��������z��d����x<�'�xB�mgk��W����  0}\+��E]�����J�Y�O�I"��N�<��˗�?���^���~��Wt��� P---Z�bE�:�v әYߠ�/���1f��K�����c�dR��w0u�9Q����}��i��q�󉔬i�#��������N�   3���ɤ�o��P    �(���#wY�����열l�i�/W�ˎG'��*--Ueee^��6I}ǎ��by�#�JittT��s�JJJ�f���zJCCC���T�~ÁD  �	���><<�ӧOk���ڹs��n���^��nٶM	����Ң�+Wf�q��i�p{��\�t��J��N&%IF".���5��������m[�T��D���� Y<x��  `��6Do�лJG��   r��Ѹ)��FF����F�#�֬�����V>����rmݺU^�7��
���ڪ�~�r;nɁ�k׮�u��Dm��G�W� ���Z���L�]+�pj�L488�s��I�^{�5���Wo���x������U�V��������#     ����:id�k$   �f n�az�.�+螻����dN��m[���y��XUU�|Pnwnnr022"�׫�[����1'ω�#
�'��zl��~Q���'  ��l/������ٳ��W^yE�D�����Ң+Vd��A%	    �������"���P    �h�y*e�̂�K���p���g���������uuuڶm�|>�m?����b��x����"nĲ,=���F��*V������  �t1J�/^�m�ھ}��?.�j��4��	 ܎�&��B��ޙ     �n��ďQ:t    ��q��-Oea������3�,e)��a���_SS��[�����gY�����j�*�{�L��m��~�S�Ne�{*��[���w  �-���~��]�|Y�m�瞛����vSr0muvvf��}ddD���$     �E��}#;_s 	   �?�nqK<�ryn���x'�W�k^�c����D"Y��Juu��mۦ����:?
���A۶mSyyy^�av;|��^|1�m�Cm���<���  ���^r?w�����N����}O��t���v�N �uvvjٲe룣���    ���gY����}e   `���[c�T5tK˲��H�ҥuY����*�H�5CEE�y�UTTLy���$i�֭jii�k�~�@@���7e�vƱ�����\�R ��l���Ϟ=���Aٶ����z��w%I�iRr0m�u�]Y���pX�H$��x      7+����]'��s    �?� p�ܥUJ�+=.؞���^
���1Y��c�tZ/^T[[[^�-~�_�>���|�ML�'	�R)�s�=�z�y�sG,�����*�f�/�-��?u   �	������CF�_�{%����]��m[�O��a���Ӌ/��t:�M�6�4MIR*�r8%���0�Y�FMM�C�����H     f�l�L"��t 	 dgţ�e9�,fx�d�=N�@Pp�m�V7+�{������w}�Z�:��P2�ԥK���ښ���\�z�z衇�g��={V�PH�֭SUUU����b۶�q���d�T4���ߓ��9�  ��J�_��JJ%]�>���\�pxƗ�O�:%˲��Р;v(�h�֭2MS�a(�L:�c��֭[�����c###��    @�d�CD^}с$ �]�{��c��
`�)^�R��V�c� ��Ƭ����)�����c6g=����ۛ�i�Z�v��l٢m۶QnGN=��:t�Pƺaz�����[���?  ���mK���Yi�;�x<���g��3�\��~��eI��ݻ��+�H������� 
���jӦM��    @�e{m7�}V��H   �w�6OU����˲��y+����������*��$577kÆZ�r��^o���ܲk�.�ر#뱖_���K�8  ��fs�]�Ν;7qכ���'z�d۶\.��^��Lo���ڲe����3��B!��      ��No��F�    @���0ݎL�����`�TZ����Ȉr��eY��㪫�Sm�{�VTTh͚5*++��~�{>�'�|2�������'  ��l/�www���[��o�>���?�eY2��;�����ҽ�ޫ����c###w      �Ͳ�_}��$   @�Qp�q���.�,��}�^w�UT�����\����b��������$�43��|>�^�Z���9�sϹs����}M�ee+[���~�1R ��b���{zzt��YIҡC����|G�x\���z��� wb޼yڼys��l������    @�e{-7�wY�S�   �w�qǼ�-2\���|�
��V�S�ۛ����������n����U\\|�s�PKK�V�\��7p=���������7ߥE��?���H  f��^r���UWW�l�Vww���ohddD���3ۅ� p;:;;�v�ڬ�%�IR    ��.����^s 	   P�q��#oU�#{�;���C�b*��Аo�9S��,�Ҽy�TYyk��+++�n�:������07�_�j��~ު&-��e:p�  0;���{�N�>-˲t��=������$��n��n���L��ڵk�lٲ���׾�Pn     ���5��k/9�   (
��	wy��"�#{�>�ץ��$#��@ ����>�eY��㪭�U}}�m�|�n��-[�e˖1�S�W��ɢ�g�i���H��f� ��l���u��Q�R)E"}���VWW����T���pB 3QQQ�6oެ���gK�Ӻr�R���     �\`F�뷩�AŎr(   �ܑ3��6.���Z��](R_��)�V�����JKK��Ԕ�Ɏ���Z�~�����n��kppP_��
�2����Z���WI�� ���Z�ݎF&�fS�}ddD�R,S2��SO=��{�J�z_��;+>O �QYY�-[�d��["�Е+WdY��     �\��rG��7%�v    Pܑ3��'o�G�N�-��r��ES����'�}?�%	�����&����<�i����ЪU���;3��g��W(��W����n������T��A� ���o[�/�s���>66��jddD�m��_Ԏ;d۶Ð����� �_ss�6oެ����c�XL��Ó^c      ȇl�َ��Á$   @���>r���_��ޱdZ��Ұ�y�sB��z{{�N��L&��ب����g�����w߭%K�����}?dr��joo׺u���٩��Ƃg����W�����c�۫�����\��  sS�5�K��dRG�U �$�ٳGO?���񸤫�k���`vq�\Z�z�֬Y#�̼S]$Q0��     ��0���k�����q(   Pܑsޚ��Δ��i��&��uLyN8��А
>����^�ׯWss3#��r���Y6lPss����������ե/}�K�'��Lu�ַUy�G�  @��%w˲t��q]�pA�t��i}�k_��ࠤ�w\�z���s���ź�{�`A�;��AE"���      r-�k���;%�r    P84l�s�˔��ͱ�#����k�h��%���a9rD�d��ɮ2MS���ڰa��ϟO�=O�PCC�֯_������.�K˖-+���Ç���4>>������s�Q�����   �f���%��ŋ:{��l��������СC��~�H��t�����O����,���Аb���    @�d�D�xŁ$   @aѬE^�Ee�T6:�x,��{�*[8�9�<��t\^�W���Z�~�)��������a�-^�X>�o�s����t�Ҽ�y뭷��c�)�Hd3�>u���T���  �F�Bɽ��WǎS*�R:��~�m߾]ֿL:�z�2M�� �`��-[��7��ͼ#]*�ҕ+W�H     �]�ad�>k�E��C�   �¡Q���V5�,.wl�H,��.Vk�tє��b1:tH###L6���ӢE��q�F���d��ld������a�uvv^���~UUUjmm�y۶���O��'��(M���ȯſ�#U��?r�7  ��%�`0�(��9�߿_����'>v���x<���pc%%%���{��ٙ�x<���P֟�      �)��c{vI\�  �9��;��W�.�����K��lO��K�HF�?��dRG�U___��M��x��Ң�7���C��Ŏ�)������1���m�ލ������:g���{�1���Y���j������lO  �\�%�k����K�.]����TOO���w�z��a	�u�}����2����Q˶�'     P��(G�|Ł$   @��=��0��յ;Z��'-�sO�.���az��cY�Μ9���.�߸�6�|���Z�j����(�|���R]]�V�Z���׫���'�/Y�DEEEw�mppP�g�C�e=�i���۩��uw�  @>̅��eY���ҙ3gdY�"�����ok�޽�x<Lu3�    IDAT��b���Z�~�<���	l�������      ����c�xL�]�;�   (,ޭG޹|��ֶ*~�c)Kϝ�衖��2}LV<�����~���i�ҥ����<MEE�***�J�488�+W�(;�1~�_uuujhh�ZB�n�[˗/���o�����?�X,��xI��Z��~ ou�D  Ȼk%�?W��R���J��p��Bs���O���Z�|�|>�^|�E�:uJ������e��\.����������r��v���<��d2�������      �������q�    ��Xh��_#OY��,��+��ڙ^)��z����8�`0X�t��v�5�|�^�Z7nT{{��~�ӱ
������M�ׯ��w߭��朗ۯ)--�o�q�e���c�=6e��j�/j��M�  �sa��$E"<xP###����n��������$]����ze���1������kX4U ��     ���>���$   ��w���EV2�t��[|��M*\�X�� ;ܗ��d2��G�j��jmm�V�ϧ��f577+�+N�J��Nǻc.�Keee���Vmm����
�CC�FGG�ח���}��_�ٳg��`����S�'�@�F�   nF�e��՗�!��L���H$t��������Yccczꩧ�~�z=���r��r��r�\J�R����kSۯ�l����%	'�     d�`G�N�4��5��    �G��c��w*�wJV2���B�J�R�x}��Bg�<�ҥK
�BZ�d��������|>566���Q�m+kddD�pX�pxF�].��~�*++UYY�����W�Rgg�"��FGG�{ށ��O(�f=���7���Ϳ���   Qd��ݡs���n۶����x�b�|>�ݻW�����'>����\.y�^�R��6��S�����=��s�t钤�e�`0��v     0md{�<vx�ң#�   �A�e�n5,�x�I�锣YB1}{�Fm)SS���T�Im���ڿ�:::4o޼��y�a���B��t�����F�F566�Tʹ�w�˥��������T~�_~�R�`:0C˖-Ӂ�L&3��b1=���ڵkה�Q4o�~�{*^�2�Q  
b���%)
i���Z�p����444������{��}H�aLf����܁��S����x���'?��{�F5::��c     0�d+�����I    �PpG���*�wZ��섴�xJ�?kj����Tҥ�X(�y�e�̙3
Z�h�|>_���:�0&�����566�X,�X,�x<>��T*u�S�^��^�|>�|>��^����TZZ����[�MW>�OK�.�ѣG'��;�'�xB�`p�����kj�7/W��Q  
b.��S��N�<�P(���I�Ν;u��%}�cSEE�Ð��U:�v�"R �>8����W�=������e���^��a�"     L����"��p(   �
�p��W*o]��眎"˲����`�*�\]�t�k�s����}�]������iƔ���Z�|*�
:�Tjbz�m�J���\.�\.��)�0d��\.��^��=�Jee�Z[[u��y���������~��)�[�ۧ��E5<�
�  �0�R�]����
��d�������[�w�|P6l���p..pg\.�<��ǖe魷���o�=��3����w*&     ���Mo�?��p��4   �s(��1��*���J�8E��5�7Fk�sͥ�=)+�z�eY�����А-Z�1!}�3MS�iΈ)���`����;�򗿬P(��I*nZ����J��0  @�͵�{,��Ç�`����(�H襗^ҡC����}L���2C�G�eM\$
�pÐ���pOO��o߮��AIW��p�._�<�N    ��#�@��ۯ9�   pV楟@y*䭜�t�	᱄��2���V����=wttTPWW%�Yj||\G�Uyy������d�{�Z�G{)� �9�Z�݈�N�]+�Ϧ;�\c۶.^��Ç+�z!l��q���w;r�\��|2M�ɸ���v���z'���x\;v��7��͉r����{zz(�    �i-c��e)�ʏ�	   8��;穚/Oe��1&X��nO\�4ԡh�r��ot`۶����o�>����F�,�N�u��y�߿_�`PEEE��g?�1��W׮���������[�PZ   g\+���H�]������7Q�M��ڽ{�{�1�?~�k����� L.�K^�w�%]]]����;�ٳG�m˶m]�pA���ؘ�i     n,��.)~�R}�   �E�ӂ��I��:�cL�׷ϖ�p���Su�i��dRgΜс��f۶�������ҥK�,k�XSS�>��O^��_������T��C�  p^�m�̱��eY���ց4:z���z��'�}�v��qIWo%��z��xf����0��x&�݊D"z�g���~W�pxb�����x�"�    �!��ѷ_w 	   ༩GS�i�mYJENG��HYz�ܸNV-��6�W��QY�ؔ�G�Q=zTjooWYYY��N�?��S�6mڤ�PB���*�kk�  L_�J��Y�W���Vr�ó�X�Fu��!͛7Ommm2MS�����ӧ�u�V�Z�J�{S���R��é����vO��nY���٣�;w*�HHz�\�e     �4�&�����I    �QpǴ�m�lK��������#��5�ז�Y���=ddDTMM�ZZZ����lxxX/^���9�t�t�F�{~G��J  03�Ւ�m����U0�UYY�H$��^��}�Q-X�@�d��\.�R�Ԥ;�1�4�vO~	���[/����\�2�t�̙��;     �L�mz{��Y%.�s    �<
�^C��v�pM�I�dY��^׹�&=�ڬ��J����@ �@ ���r�������@iq#�PH�ϟ�a�]���=�_��D����D�����0=�
  0C�Ւ�$����ȑ#jhhPGG��n������o}K˖-�֭[UYY)�0��xd�6Ew�&d+�kǎ���X���:{�����:     ���6�=��M�    �wL?�!_]��y���1=uTj�[��jU9�%+1~�Ǆ�a9rDjnnVuuu����l�֕+Wt��eE"��s��P�N$dY���tR�*��D�r%=  �\5�K�400�`0���V544H��?���.mذA��w��^�D�ݲ,��i����\.���I�����~�m�ٳG�tZ�dY�z{{u��ŉ5     ��([�}��H   L�1myk�p�J�����Յ+}+�՚����ኌ�Ӳө�>fddD###***Ҽy���ؘ1���N�500����������ux�Z?i�X<-)����G�fA  �\s��H$��ե˗/���CUUUJ&�ڽ{��;��~X˗/�t�M+��%˲�J�f��p#ي�e��w��[o�������P(��g�NZ     ���,C�R��?}ҁ4   ��@�Ӛ�j�dJ{����e��)��e�����.�S���l��E�X,���n]�tI���jllTiii�R�������ו+Wnj�����X�L��5MI��c��A�|�r���  �~s��.Iccc:z��jkk��ޮ��"����������٣x@��풮�z�^/Ew�Y.�K�iN�Tf۶�9�7�|S�Phb}llL�ΝS0t"*     @�e��y���   �
��<��$��D���Q�4O�SA���L��h]�e����l뺏K�R���Uoo��~�U__/�4�|�I�R�r�����Fo�1�ǧ�cezg�MC㶤�_��~��ry����fb  ���Z��Kv�l���Wr����!���Qmmm2MS===z��'�`�=��jkk�D�sO�����ݭ�_~Yk�TJ�.]Roo�,��?k     �$�&����c�    �w���z��^��eߠ4XRo�M�@I�~fA�V(5xFv:y��F"�9sF�ΝSee����TSSC��&X��P(�+W�hhh����D'��z7ڢ@4-��D�m)>xNE��p��
  ���l[��֟sw��t�����^���M��K�.�'�P{{�z�!͟?_��{:��̋Yg�b{OO�^{��g�΂��<��ʺ�'I��HJ-��n�h���8�{&�a�g<��n�\�����eG8�Ox�}�����}p8���iu�n��P�($q�+�@��H$������ �U��%P$P����+X[[��<�l�������&"""""""�'�$��G�0>���DDDDDD��w�J8	}�<�����'l��ֲ�Eo����ܯ��<�_�g���X��P*�P*��(
��4FFF�N�Yv���(��(�(�p]�����8>m'��
M��ۍg��N�}��"Nr��eYXZZ���&N�:�t:`gZ�~��?_��W;xY�!�2�p�Ew�{��@Q�}m�����o`ee��N�\.���u�q�Q�'�,�����������,���5~�0D�M������a����� 4u��uxv��n�-��d�--���|_) R_��(���"��#��C�e$	��� �L"
s��c�&J���"���!>��>l��Qq��	�:�lN������<�m��I�σ%w`��M�|�	��8fgg122 XZZµk�p������:��� �Lq�4B��{��;��&IRgb��nܸ����'�d2{�W*,//��l�TL��.�NDDDDDD4Ⱥ�n��#��ܩ�HZ����p�u���e�xg���d�N?�˓&������.��y��2��2  "�L"�L"�H �_��m�R�t���'�d�8>��p��q�G�]ބ�@�cǲ}"""�~�[r��Y��(��.�@�VÕ+W��q��i$	!�駟��ի8}�4���/�G�s�KUU���)��׍��$I���w�v��x�lnn�Y_�հ���j�zR1�ǰ�NDDDDDD�D��}��Z�w�S""����S���1�h����tBXp��$�
�G`U6aW�~�90���f	����4�����"�u8����e�&������`����������	z��V�Z�Z�z�v��6&�PS���'�8�K����t)���[Fh�"$����I�uq/`�%��Z��?��T
�N�B,�+++XYY���4�}�Y\�x�s�k�8�y\�=�Ս���,�Pe��=��'�|���z�\n�m�j�L�sB7�~ڏADDDDDD�����������C"��������h@��N�K�H�@�tX�u�_��J���K&~"Kxd�I<>-�^����^8��L�D>�G>�YQ>
!� �"
u�;�'I�0`��&��&Z�Z��C�r�pkV�����h�6��O}�u`斡O=
p��>!��s�xA,���\��%��WlJ��8u��ѝ� 677����H&�x�����Ow��$�2dY��3՝��kZ�i�������Zm�m�r������p�e�7�?������h�t;n�|��>$!""""�=,�S�S�#�!��ex��w�C�<�ō27������S�0n��V��܄�|�	v�v�v����|0�����E�4���g9(�q:��q`Y,˂m�0M�i�0��y��%	Zb[VW�i\��7�8�R��\�	��A`d��DDDD�J߿5ɝ%��J�J���8fgg122 �T*x����o����x��g��|�$I��ϩ�tR�6��y��W�»�۶��V,��dP��O**�EQ�x�ѝ<���,��~o���,�PU�� v�F�QD�Q�޹���n���7��$I�7��k5���>%"""""�-,��@�a�S`�W��w�i��d��O �a<2��N�8j@n�`3�}����yn�j��.IdY�3rwR�I�djb�V����$�- @��r܏]�CF�FG��BDDDԓXr��Z��+W� �`ff���$	�i���~��_�ҥKxꩧ0?��ɕwNu�<�_O:2���.���7������{^w��P( �ɠ�j�dd���"�gW�#""":j���l�^���h�4MX��P�TU�x�T
���@$�eY0M�V�f󡟇����r; �~�`?|�����h��NCRT蓏��l��l�}��m9�p��Ȳ���<;�3�2��6�jv� ���_�q��9�F���q��4V�Ad�n���h[�B{7Var 9�;
QO�-�?/-@DXr��f����%���bffSSSP��⣏>�G}�t:����x��'�D |6����~D��{���(]�6|��x��wQ.�
�m��f����da��I�4���������/�i�T*uJ�G�^�q�Ε�nܸ �F�������,��� �2�A��D��@���U����Y�+�5^ɇ$DDDDD��w8Zr
J(3��>���^�y�R�R?�Øys�L)eLim�fN� �2���P�`jl-9��V���s&��֭���#�����!����N����2^��~?�eaee��똘����,��  �T*��_�+���ӧO㩧��ŋ;e�ݩ��N�(J�s'!VWW�����ի��/�v����f�,�Ё������i�뺨T*(�J��N��čF׮]õk�p��)�>}H$�<�F�j�f��͉����C�e���>�!""""�=,��@����a3pE����acq��ō�?k����#���Q�Ę\�h��h��4+p��k�Y�N@	%`kQlAd����*����%_c>,�6a�W�8�w"""���;����~��bss[[[���$��$$I�+++XYYA2���˗q��e�b���Yv�{�W� ��2�{�=|��h4{nB�\.csss�$w�{�4p�zm��3�l�R�g��Z��)�'�I\�t	�O�F<G<�m�(�J�T*<y���t���z��i���������Ṁ���(>{O!�ێMI$���GIn���d�dH�
I����R��D48Xp��%�
�c���Ⰺ�{(����א�6�C����0�|c�$�BLn"����g��YMx��lB���f�r09��@h:j�����"B({�
�6m�֎ܓ�Rr�VreZr��(DDDD=k���< Xr?!
�
�t]���&&&:S�+�
^{�5����8}�4{�1\�p�P���new����"�$u^w+�7\�r�1666��n�&��������n:�`0����u�n�����S��n*�
�z�-�����x�"Ο?M�011���Q��e�E݉�R�}0�7^�!	�!�mB8歏��玵Sh?����H�I� �Hj���!���u��q�"�/,���S�i(zfan��w��zr�r��gy���$� º�pL�.{zm�U@�=H���, 	��A� ��x��$��
�S`
�+��drM[B�t�(�h�6�M��p �o-�îlAF���~G!"""�Y�x���������M,��aX[[���:R�&''�N��Mu����;����ҥKx����;۸��,��Sx��r{����a�2MKKK�r�
�_���u �@�TB6�E�\�Oz`�$!`�Ω�DDD4x��͛7Q�V��r(�V��>��\�|P���H�R(�=_�'"�ew����k,�Q�<ۀg��Ym�����d{! p, �}�K�)��� >[$E;��D�@Xp�� ����4�������~��Pk�P;�%�T ;��]�g�����Wy� ��˛,�݇.�+��i'��n�T*!`rr�u�s{&�A&��K/���g��ҥK8�|g�;���OQ(��I�����2��)�_�v�Sjw���w'Onooòzkg6��@  Y���}	DD�1ϊ    IDATD48<�C6����v_�4l~������x�g�N��(
��ǑL&��f�l6��ID�W��i��z�EDDB��2�لg���M�=ǂ�f���')*�@J0
9��G!ɊO)��^Xp���FG���JpE��А�$	jl���Q������.�_\��X�`���Y����ud2�b1���att�@  �.������EQp��9<��8{�,���m�m���ߏt{�]���Ni�J��y���w-����B��|>�z�%d:Z�p���I��'���j��L&�4��rd
�����.\��O>	M�0??�j��\.�q�!""�Zpo��I��h(	�Sd7��:\�1t�b���m��?;�!BP��»�B҂����i�H����i����z�]>��#8z
r �w"""������x^����\�%�#�@�VC�V���2��x��i;�at]���X\\�$Iǹs�p��9����9�v�t�ݒ;'���0�v!���������%�r���s�B�\�����(��p�ĝ�DDD����y��]�W�^�͛7��/��� �D"�h4���Ns'":�;���E��}JCDD�@�&�vn�:�����6<�  �� �PJ(%��_������R�	��%ؕ-8��ӑ���4����Q������.�+��i'�	!��*��*nܸ�d2���Q���BU��}������������4���8�<.\��x<�g�����K��=�;ѿ�0����m�ם*�
2���ױ���F���~��T*!�ϣR��{G�.�  �m�|NBDDD�p,�����P��~���'���? P���(�J��x̍��n���1>�N��C""XB�5p[U��*<��;Q��l���]�C�d�zt��N@�t���i�I��@zZlVyN��w$ jt��,$���=,]|�����K�GI�r��r���ׯ#�J!�N#�N#��ҋ�mcee+++x��1>>�3g�`vv���F����[���n�}�������~������ξ��lbmm���XYYA�R��}�@�XD�X�):Q�P����,�#��IDDDD��R�`uu�;<S=���ￏr��_��_�\l�����&��9%Q��_���+>$!"��#<�	�Y��,C��߉�ޭ	�5�t��C���D�,�3�/� HZ�����b�g��QB1�s�!��]<WX�������p�܏��R	����p8�T*�T*�D"����������_� �L&177�Y��ƺ��6������2ln/��^f?!
�666��d����B�pׯ��z�R	�b�V�(�*D"�2��0 �L%^ܕ����U>������1|����z��������bG$��S���d`Y��	��z˾�cB����	CDD�5�p�E��
�7<'��ɳX�-��9�IA��!i��?���w��(�8B3�`��+[.�K��Ɂ�(��Q�����.�+��i^��܏[��B�����dYF2��Lx�--�T*�T*�裏  ��cvv��LNN"�~���;�^x�s�7���\�0lll`cc7o������'i������R�p�"�.�B�$�����(������d�Ylll��w�R	?���o|�����@ �)����
Ѱ��˼�g�?K���p<ۀ�(�m��9<��O�Նe�a�7!�Т�P�iH��w4����;ѝ$	Z|Zlv-���nԕ��%��FG�(����B���坒{�%���y^g���7
��L&�����������q����:]�166���i���b||���Pջ_|�������|̃�=����>޹�A!P�V��籹��B��|>���,��Sh7M�s�p8�@   �/��<�����(
~G��F/��"��o �J TU���<n޼�+G��~�曯���������4�pjy�f��4ԅg�`��J7�DR�b����߱���Dw#���P���k�p�9���H�-9	-6�b;�	Ӆ���xAp��_��6��6��� �L��-�'	D"�}��@&�A&��S�t��㘘������$����|7GQ"��i�\.wN"(����r��r��.�@��B�VC�VC��`y�z��i��  ײ����ω������������c|��D"�s�[EQ077�L&��)D4��Mp���C�Q?�lN-�Q��>!��Q��(B���F�FG8՝���Nt��"����`�}��j jbZl��� """���;��yq"����,�B�P�<dY��c�"����ǹ��|>�|>�O>�d�m��#�Ht
��d�T
�d�D�3��4�M4�M��u4T*���N���%˲�h4P��Q��P���ܩM�OQ�b�Ο�-�D��ۉ����lll��~�e��_Ʒ���Ή��,cvvkkk���n��eX�7|HCDD��m�`W��k~G���YmX�����(��8$m�13"�w����>���]�C����G�Oւ��Pc���NDDD�#t!�\i/��"���K<�C�RA�R�SU�p��D�QD�Q(J�i�a�0loow�]�4�B!�B�=۽}��窪v
�AQH�Եtߍ�8�I�m�0���Y������f�F�Z�f��结���vg��V�a<����$�2�DgZ�Z���&�Q����f�~��y�V/�����ov�w)����y���¶m���n�ۛo��C""�iB�i�`W��Ym���]���堆�����߱�z�D�$)��4����/�,<��A$����P#iۉ���z�.�_X�b^�%�^�8j�j��
��$A�u��aD"�B!�]��;�ݶmض�g{JQh��g�i�'���-ͷ�m��m��f��v��ӭi �Yn�l��r��TDDDD�S.�����w��Q������7~�7>;�QU177���U��!��ӭ��x�|HBDD=Ix�ky��m�'�:�U�ӪBѣ�P�I�#�,܉�$A��@���*p��pͦߩ�!I�%�������������C�/.�yq"��{�BtJ��bq�m�,w�#����B��p]����ߏ�e�[n/��N�'D���)��̭a��랈����i�X[[�;F���rx�����SOu��ALMMacc��dDD'K�2H��ބ���i����v� ��e�}�F�рAKNA����D�sXp'zX�5��I��Zp�E8��˃��DR4��h�1H꽧EQoх�s���,�����Xr�o���j��ju�]�$h�UU��*4M�,���(��Ή��`�<��{q]������q���q�,�E�ۋ�m��GC+ ��Rw6��d7|LEDDDt8B,//�I���ʕ+������Lg]<G��D�R�1���:����N>�����nMlg�l�yVfnN0-5%�;Q�`���Ɂ0#a�3p%8����0I����Pc�PB	����DDDD�t!��7��I������Ga��.�`q����a���=�Ɗ��/Zy�=�L&s�o�`~�ӟ�7�7�F;�&&&`��1���6����>$!""�	�Q�U���v��5�p�נ#��3P��ߑ�|��TQ"zx�56
}�B3����!)�ߩ�9B =�����8%�d�����h �NrW��M�-�w;�D����v"zp�� �H�+�G+%���-�R=�j��|�'�=,˲��l�:Y�1==���D4�$I���[*����>%"""�8�2�W`�Xn�{r�&��%�����<)��'�39B`d��,\��Y��,�3'LVP")��ȁ��q������Nr�;��܉�N�$I�B�B��'��W՛>%#����*(�/���1�Z�Ղ���*{��ʜ����۝?ׁ�n������؄�����+W���n�<�L��c{{���XXX��A�P�1����3'o�p%����b�Ѹ���n㴪p�5��h�H
��4|��':)�E�A�c������{�²�1���N�=����DDDD4t!���
^��Ew.�ǒ;�ѓ$	��#
u=h?���w�9��Q�u����w����Zvy~�@��>�߮�Qw{�;B�"���4M�c�w�}333��u###��j�,��dDDǧە*���C"":i�u`W����<.EL�^�Ӫ@KNA���܉� IPBq(�8b�لۮ�iW�-���-I� ��[_�'�1]|���'�5Y���:t]�Zlw]�n���V͇tDDDD�4Mloo�c���>� �<�Lg�,˘���|"H�$�+���*���§DDDt"��]��.oBx��ih@ׁU������G��Dt"Xp'�ۭR��G���!\n��Y8���d-E�A�u$+���I���K�DDE�e�Ah�v�;�����*f=����L&��t�㰴��Gy�T��.�"���h������u����ś��*�j�*��5�~G��Ym���FGH�BRX����W8Q��jtjt ��<��h�3���$���P�(d=%����:=]<WZ��$w"���e��@Q��
MӠ(�>��u]����V�;����o�Z-T�U�c��?�_��W��e���N�+�5^��I����	v%���q':N��]C`dj$u��)o"�q��C�t��Q �pmxfs��n��Ymw0��I�%��G �Nh'"""�C��$�T*ũ|DD��x�v	�{B R-㻵M�z�BGDDD�mkk��ommO<��Dg](B8F���1������k5�x�u��q�J7a��~��+��@��֏K����v%\fnn$������@b����H�%��Nv�	ׁg�:�w�nC�&������$E�)�B�n}��/�BDDDDGF�mi�S�I�,w��DDD�'�@�^��նpڱ��CDDD���@�R�;�P�r�
�}��=�FGG����S""��������?��\GD4���v�m���,#"	 
 T���0LDe�EH����*A6��w��p<�����,-W�)�`(a�	���J�D�e�a��i�Y�5�}j4�w�#��(� �J(%߳^x.�cB8<{�pLx������o�$CRTH����Hj ���y�Sى����D��o�;�h�p�Q�o����v""" ��~rVVV���#�u�E"�B!��m��nC5o��C"":	�� 8~��Ձ�@�5��B�����m�4	Ղg�w���Mx�6p���q�� Dn-{֫(�0�0�P�A�VQq�(yQ�.��6
�6wp���3��]E`d�]<,�0IV �@ �����N�ݻUx�\@��/;S� >��	��M�$)�,��p����@Q������z�.�cɝ���\�E���L��g�.�,��q�r��C��<�����'�س>�J��ND��	��2��ɫ>�!"�� B���̯��Hh���TSq�r3AI��qn���l��aJ�GA8�Z��	 �Z��z���si� ��������+M��8��'�i����@֣~�!zh,�;Iޙ����I�����N�n��_�shk�=��H�z.Tσ*<$3Vg]���DDD4���2�ܒC/�~�:��=S�c�dY��ǔE"Lݦ����%D��C"":Ijt�ل]��������(fB6f�ft�uN���z�E��XF(�!���Z��8�0�#�M/�L�@�X�e�~G>R�c��.AKLBKNw�xG�Ox|���������.��ʺ�1��������E�#�V��|>�����:Y��FQ��|LFD�p�����C""�C =�l�5{�Ħd,�������q��)��������J��&�R(e0`\V��8��	l�Q�0����#WmcN}B��l�m�_��r��'܉������������h(���f���'�huuuO� ��$�D�פ;��
�A�|JCDD'N�_@{�S��;�>c�M���"am��fp�q<�,�P��@U�κ�O
B�uw&�{��q�ng�Q���	����g� ���4N'q�J�j�E�P���w��5�ho~���(���q��w"""""""""""""J�R��Ckee_���[��0E9�"�q�6����{pk��_$5�����5�Az4�����F�:�vh�CnW�$�A��Y���EU�}'�����mX�˲`�&,˂ah��0㡿Ξm��-CpA���$��Y\7Ӹ�w����m�]���5h�IR3~�!:܉������������h(qZ��A�P���xg�$I�D"��Q_�V�k���I���o�����U�������y�8�p�5��4R]��D��D�D
���~�$A�4h��p8��>B���V��f��Y����߅�]�*[8+I���1>�+�(>�2P���o������NC����DDDDDDDDDDDDD4t<�C���;�P��r{
���w܉��9�]�.��Ч4DD�7-1	�h�i�̕<$I�l\�cj�F�J튢 �!�#�!�AӴc�|$I�L�O�ӝ����h�V��^��V�����m\��,�j��|a�4��ޯDp�f�����x9�
�ͫN����~�!�/܇�k�Ѽ�K�cр�?�5@�9>"""""""""""?5����==���-<���{��m2#Q/��� ��O��>�!"�^;o�Sx�ylϡ5\7p9R@�-@�����{�d2�T*�D"q��O�,ˈ����u�a�R��\.�R��q��o�sa�n ���P_b��x�f��q�����[%wE����Xpf��g��%3��� ��{/�z��w������.E��PU�pe""�u+6�|Ň$DD�K$YAp�,�ͫ�h�}��t<�e�x��(�NE� 4M�����4�������똜����$������"J�����k����$+���Ӹ�M�휊L�?�c
υ�����)������DDDDDDDDDDDDD4t�ͦ����y(��ݳ>�V��������Mp�W~�O""�)r ���)���#��dT�3��8,óZ����A���addd�T�a�F�Fq��)���R��|>�j�z�ܚ�>�8;2���9����V���WB�̯B�&�Դ�q��b�����������������a��e�Y�V�Wp>�!":�n���Kp6n�����z�M�3��k��ƈ.𴶂K��c³𼪊t:���1�R��?�hG0������`Y
�����O���Ha�M�O���JI|t����Ve�m 8v���ޟ�$��NDDDDDDDDDDDDDC�u]ض�w�FXp'�~�oz;�ƛ������zY =�l�5w%�������7 ρp���h4���)���w�9E�0==���i��md�Yloo�=��(!�(����t?�$qu��^�;�2�� 8~������w"""""""""""""*���;���u,�Q?�Zp�E�QO�$'΢�q½K},��K��J�x����i������$B����P(�3g�����(
�f��T*�}�۪"�zߎ���cg�F!��������m�af�!8q��Z1���������������h����w��w"�g�$�[ggVa-_�!�:I�_���!����5OV��D����خ�:fff099�i��H�$���all�v[[[��ڂ�����YF��+�'�1d..���Z��R�k6al-B�:I���CĂ;˲��@��Z�}�E�,��-���������C""������U�س^�%�����Da��{o'�H`vv�t��R7�P������666�8�>���1�<���i\I�o    IDAT�N�Օ6���'��4�6`l-A�|����_,��Pq]��t��8�<o_I�w"��&�7^��Q?����&�V 0����u���O��S<�����=@�4���cff����d2�=��.��y�����,>�4�}��vJ��'�C҂~ǡ!Ƃ;�{�m��'�ME&"�%�$�+�;�-W?�)����iD�KxF��Ej޽�y'�I���#�H�PB:(EQ0==���Id����=J����ң��
���> ϱ��ZDh�Q���7�+@DDDDDDDDDDDDDC��{K�(>$!":�n'�4�|݇$DDԏ�ob��g�q�r{8�ŋ��}���'�2����/|gΜ���{��g61V~�xr_9�"�2���k��.A8��JOt\Xp'""""""""""""���	�Ŷ�}�LD�k��?�x�E�Q?q�5�������W��������+!��/����x��1::�CRzP��`vv_��133s߫S��<m���Qө�	�<ϱ`d�A��߳�{�"BDDDDDDDDDDDD4`��I���zZPD}�:Ֆ�:�W4^OQ����n9s�������}�%�%5e�p��J��m��N���?�gG��H=�ou��_�����E�ʫX��߅UX�{�����/�[����)ೳ�����o1�z���XXX������Q*��z_�X�?�>:�w��ɚ	���m��^�>y���1��ڈ�����������h�<
��w�;������#w^�^q�o��~' ��V��Y��q$[!"":9�m`������^ ���I���������/���DE�+
��C�T���2���]��T�pY-b�����*M��ޝg�al�*�ˊ�qhH�"""""""""""""""""""�#�Z}��w�����e�r; $�I ��s�Xn`�tO?�4����9�_8F���n���Lxo�ق�}���c���	�DDDDDDDDDDDDDDDDDDDDG����ڿ�g���%I��%����>��0>��S<�䓐���ڔ�y0M�e��<����:����a��@�$ȲMӠ�*4M��iP���.IN�:���q\�v��=�fU^���"&O?��3
,��b�k4`�W_�;
܉���������������������g4��o�)�o��w���������ŋ�u�z7n���s�N"摰m�F�f�a�4���8Α=�,��u���A�B!D"�~d�sRB��x�	lnnbee�׽��u������G��T��	'��i�!�7H����DDDDDDDDDDDDDDDDDDDD�ؼ�����о��]��|����۵�����x<������@L�D�ZE����m�>���<�V�Vk�m�� � � �!�#
�H��5==�T*���E����w��E�����z˅�W8Iv%Y	@�����DDDDDDDDDDDDDDDDDDDD���+�����f����0���੧���v�]��)l�ɲ,T�UT*T*��k��q]�Z�Z[[[  M����ǑJ�|�Z�K(O>���ud2!��O�o�?��Y��<c���N�U�@҂PBq��Рb����������������������A����/�����]����?�c����ws���ʕ+���?U=يg�^G�P@�T�:-�_ض�b��b�����A�R)��i$�I(��w�=$I©S��N�q��ջ�L�6��5��ԩG����.���[�>�(�@Ļ�;�!	�����7�]��%I·��m��o�6dY>�v����"{챣�zW�F�R	�\�v�؟��i"��"��B�e$�I���add����X�/_���J�R��x��G��?u��f
m�9ᔟ�s�:�鋐֑�h�EDDDDDDDDDDDDDDDDDDDtN�����?E��׻ޮ�:���O>��m�T*!��`nn�abve������`Y֑o��y��R��R�Y�122���	�R)�� 4M�c�=�L&���5�nW&�K���S���3�4͓z��X0�+�'���[<,���[������-w�}bb����055�Pϳ���h4z$�k!��"���P�Tz{���<��y��y躎��	LNN"�sss�F��z�*����xk8����U1N8�g�vveZjڷ4xXp'""""""""""""""""""":�v�#,��7aW�������O��O����<�իW��SO!>��-��������Mk?�0������u���`ff�x��L�T
�/_ƕ+W�j���G�g�)#� S�^�?	Ver0%��-�� DDDDDDDDDDDDDDDDDDDD����6�����Zn��׾�?��??�r; 8��+W���C=�4M,//������:��$�@�P�|���{�\B��B!\�|�t�����9�Nr	g�	&��̯@ئ�hp��NDDDDDDDDDDDDDDDDDDDt�+�b�/��^�w�,��������d��k��F7n�8�}[����occc���x�L�����"�y��r9�r(��K�.azz��wj��%o���rr�� <F~�� ����������������������zU�ݿ���{���Ԛ��O��Op���c͐�f��111���v����U
���p��6��dp��)����xI�p��Y���v�S��ߊ_���ZpN4�.�l�*o �����ip��NDDDDDDDDDDDDDDDDDDD�E���Zn�u����p��r��uD"D���:۶������-N�>V�V�~�)��(�H$N<���E���r��h���U8�Gp������nC�cP�'����q��� "��ٻ��������٥-�Œ���6fq60&��%!����KIK�$p�m�p�tIo�6m��M���m��6Iӛ6[16��7��lɫvk��4�r���3#Y�g�f>�׋W^<���|��X�{�             �\��u��Y��^�W��ԧ
Vn�$�0t��%�I�����~�ܹS�����(
i�޽ڿ�b�X��5MSCCCr8joo�ݞ�l��uW�a]귮"9!3m�.�(��              �&���t�O�%#�8VSS�'�xB������u��%�����illL�`Pmmm��윲p���b���n�$���J������a�/�M�=���ws�z�_47�I%FN�Ӽ��k�4��;              �/��l��?~��X(�Xuu�e��3&&&(�	�0��ӣ]�v)�|�H$���>��F���ϧ���)���h@��Qk�;��|KE�JM�X�6f?
�               �⧎����V::�q���(N�XL����<�T��wLO��P8����<��;���Ȉ�;���3]��h��dܒ�1�Qp              e/51�C_^���PƱ��*=��jkk� f����ڵK�@��^o�����4<<,��%��v��TVVj޼yr8Y�;#�tw�1y=��t1L�P|�d����G�              �5#Uן߫�Pw�1�ۭ��r;f$�Hh߾}���a3~�����p8�t�_���B���S��kC����܎�׆��	�Bc_�w              P�LCG��a��^�8�p8�O|B,� f���A�޽[�Hd��b��z{{�H$�v�/x�3%w�={5�)v\���t�=�s/1�#3��`e�V�             @��������e��l6=���Z�|��P
��^}�U�:u*�X:�����&&&TQQ!����ӗ�M-Lu뺖�E�s��tJ������ً�;              (K�������i�c��w����'B�1C�RWW�LӔ$�ԩSr�\S�~�*++��ޞ�0o��Z�8��5�/��BcJG'
�.f'
�              ����_ױ�yD�e��ͮ��z�[���P��ӟ�T]]]��lr�\y[��󩵵5�13�5GU�u�m��$FOf�~ފ�;              (+�HP���;J/\�P�Ї,H�R566���׫��K�=������fMM��̙���+1������r�=Ǜɸ�C]�S�o�@�pT֨��wY@���#t            ��b:��V|�;�М9s�����^���L&��K/��r���^��D���j��՚;wn^�ollT*�R �8V�խ�U�Y�O��S=���A6G�v����;p9�I6[a�             �J�?�����1�r���c����Y�
�f���
�����8�H$�q�F]{�?~^s477+�H(g[d�����h�615����~��lM�>l�              �B��.�����>��������Pjz{{��3�(�Ng-��a��nݪ��5��fS[[��nw�13��-U���-�f������=pw              P�xXG��C2S��c�W����_oA*��P(���׫��_3z�i�ڵk�^}�ռfs8joo�ݞ�6��^9�fx��hOA���B�              ����I�e�wtt����P
��^|�E�ݻW���r8�7��������x��ښ�XCb@��Cy]����ґ`A���A�              ����j���w�\���>&��iA*�v�����͛UQQ!��s�s��^]]����,GL���������@A���A�              ��ThT'���Y�=��jkk+p"�vZ�~�b��jjjr6������k��l�l���TYY�1n�&u��GnG��F"�T8P��0{Pp              %��w?��ĩ���˗��o� f�h4�M�6��ɓS�~���٣����enI��ljkk����8V��5�cy[;�d�_2͂���G�              �����������#�<"��fA*�6�ah�֭ڹs�����t:���ݻ��ݝ��].��Ν���;*��\U�]ܓ1�-գ���;    �܈ӭ��eu���4ui"bu�Ye��Ԑ�cu�ɼDD.v�        �rF<������>��������0uww�ĉ���r��Y�4Mm۶M^�W���yY���F������8kܖ���>�K�Ui�0׼��9}�7���(�   ([�ݕ�N}�6nUL�ӝC�W�6�p���i��4��%�	��mVG       ���~�s��:�1�|�r�\�҂D�MFGG�k�.������|}�4��/���oW]]]^֘;w�"��R��Y��A]�Ш]Å�i$�J���j(�z(~�8    �%����E_�~V�,������u���w�:x       �BѾ:��_e�WTT�����0[��qmܸQ�VCC�l�*�L&��s�)��S��ZZZ2��������p�h'��[ŏ+�    ����G�}z�ۋ%w        ���'d�S���sO�v���{�nm۶M���r��VǑ$E"=��sJ��y����J555���Vz��f6F2�td�`롸q�   @Y��>{Prώr��A�        kv���_{&c���Uk֬)| ��Ǐk���J����|V���s�μ����,�=����a������P�CQ�
+   ��A�}�y�W��Υ��K��gJ�        �����_~+c�f�顇�Z�E�����ƍ5<<���z��L���K���y���tjΜ9�f2����d�˪���I�p�VC1�   @Y��>{m��Qr��ٌ�;        �3��?S|(��j�*-^�؂D(F�TJ�7o־}�T[[;kn|رc�FGG�2w]]�***2��jD��
w�69q�`k�x͎�H    ���g�r/�Sn��(�       ��HP�?���q�˥{�ׂD(F����/� ��'��cu��N��e�%�ɜ�m����ܜ1n)]���^�}����T� k�x9� �x����#2�aɘ�ؤ�tJ�p �\��V6�]��娬��W'��V��Z���  ��A��tl��I��,�#�����q���H�GnӰ:        %g�'���t뭷���΂D(&}}}ڿ�TSScu�699�]�v��k����^�WUUU
�Bg��$���נ��ޜ��V�i*99,w][��B�
����⧎(v���'5>��䰒�A�&�e$�9Y����Y� wC����N�o}�<s.QE�����A  @����[ɝr{��       @~�&�5���2ƫ���n�:�X�B!m۶M���jhh�:NNtww���E������MMM
��2�7=_�4u}Հ���2��������V�VW��w�ĤBc��ܣh�^EN�U������N,�++1z2�	6�<����m�TѺD��+�w�lw  @�Pn/]�Rr��^�(�       �{��G2b���;�S���$����^~�e��)��ou��۾}����r����xT[[�`0x�xU:�%�q���{3�T::.�����af(����N*r�M~Q��_P��.%F{��un����1Ň�i|�����*�d�|�Wʷ`�����y��A �lE����zɝr{�;���;�zd��;        +�ש�������ի-H�<xP���%Yl?#�kǎy�oll����ٻ�K��?�C�Z%����2F��E�tJ���4��YMzA�#�e$"V��#S�k�B][�sյ���[U�|�j/�U��V �ـr{�(Ւ;���q�M�       �\��Wd$���z׻�rqͥ����h��ݪ��+�r�'O��ɓ'��ٙ�y].W�]�+�ZRӬׂ�*B*2.w*!�ӝ��P|(�E.����_h|�/4�o�ґ�g����͖�2��`��kd�?jd�?��ҶL5������Q��5�Q�  oB����Zɝr{���       ��IG'4���2�kjjt�7X�V��bz��UQQ���:��Ԏ;4w�\�ݹ-�744d���j���_�l�ThT.K�Bѡ�����m��ƶ�@���tn�ݮ��:��׫��^~�_uuu������{㟊��i��g�ǕH$���D411���IMLLhbbBccc������E��P������:�W�Gu�ܯ��o�ݝ���  @��^�J��N��|Qr       �z���nz�w�{{0MS۷oW<Wuu��q,�F�{�n�\�2���n���h|��ﯚt@�T4�hԛ���IM�Pp/S܁"�9q�����>�����;w�:;;��Ң��f577���INgn��=�<ό> D�Q���_����������FGG�{�T8����v�O���T�;V�����  �r;f{ɝr;(�       p��d\C�|=c���{{���։'���sމ�m����hѢ��^f�����^ѫ���9]+#���^Q���P\��;����+��h�������y���hll�5�|uvv����(�@���Tgg�:;;���:v옎?����B��k�����m���U��[�>5���^�"�  Pd(���Zr�܎3(�       p~F^�������n�I�ǂD(���1�ڵKuuu���V�)
�ij�Ν���r:�����U$9k��U���@$���S����w���j��oi��R:��9����l�2��moӂT[[�㔅����|�r-_�\������z���u��!uuue���J*4����+ߥW�񦏩�p  %�r;�j���)��(�       0sC��Ռ1�áիW[���L&�m�69���[�����G9����>��g)]���@�=�ke�
�n��	ŏ�;P f:���?����\�;���n�[�]v�.��2-]�T���yHY<l6������֦�k��0?~\{���޽{���7�y��v*|l�z��Y�Y�q5���̹$�� @APn�TfKɝr;�B�       �su��h�k�+W�T]]���O���q    IDATw�V PMM��Q��+�����6���^UU%�ۭD"q���|!m�����z��N*����:�렸Pp�,����������#'��>�OW\q�V�X�e˖��*���n����5�|�{��޽{�s�N9rD�iN��td\�?�����_u���}J5�o-Pz  �k��q.�^r�܎s��       ��7�M��o���I�OǏWWW����)����䤎9�E��lN��&�߯S�N�} �ۀ��9gkM%Pp/3܁<I�5�?��s�tlrƯs�\Z�t����Z]u�Ur8yL9{544��o��7߬@ �W_}U�v�:w��4|�'
����T�}�����
  \4�혩��:���-��;�v�%w        �KG���Ì�͛7ςDȵ��Im۶M�������:ά��k�i���9����jxx8��wUU@{c͚~{ڋ�
��l�t��D�ȱ�İ����d$�3z��fӢE�t���kŊ����s��RWW�[n�E��r�����e�����
��Ӿ.|d������v^��{�V���� �"G��k�/wr/��;�v�/J�        dy�e$"�k֬)|�T:��֭[e��UWWgu�Y)����KK�,�ٜN�S>�O�P�q�=�wL���v�tJ�x�]��w?Ӝ�����~�eo�挋�>�O�]w�V�^����?���������߯W_}U[�lѡC����=rr��|�^���;��xϬ�� ��Pnǅ*��;�v\(J�        �m���������W_mA�ʾ}�422��jJ�k߾}Z�p����Մ�~F�]2��ݧ�Ă��3�td��{����f$"��:���Ųi	Ĉ�5�_��Ͼ����l���u�m��ꫯ���7�өk��F�\s�����a�m۶M�Tj�ׄ��Rןݣ���T燾"߂UL  �C���;�v\,J�        �9�[��}��\s�**�4򣷷WT}}=����b:z��/^��9����p8�N��_V��1���^�JG'�:?��Z-#Rl�[��V|�*Z�V\�j��ƶ�P=����'�y��fӲe�t�m�i�ҥ�3������|D��{���y=��󚜜�����u��ש~�������si� ���܎\���N��B�        i����u|�*6��mB���mۦ��j���[��8p@�-�-G�K�ͦ��j�����ɐ:c:���d�����TB6�;��8PpGQzs�]���c�r7tX���C/��{O*|l�9ϵ�lZ�b���.��� �RSS����=���۵y�f=��3����.��ض(��O�|ǧ�r�gx�	  �܎\+tɝr;r��;       �����^�׌���z-\�Ђ@��ah�Ν��b���[�.g�PH===����ٜ555wIZh�����e::!guc�ׁ�(���c��v�|˅���)�=^9�,J&�&�u����;�6�M�x�;t�]w���� �0S�G��v�֬Y�F�=�]��]_��5��?��_W���8-  �r;�P%w���J�       �r�~Y����V���.�ȯ����Ouuu��|V�)y�i������t*�J�5��ohSB��s�TV��8�2A�E%W��ьr������+ew{�L������JM�����˗��}/��"�r��v�Z�^�Z6l�/~�E�Ѭ�&}�����_�n�{��n��}  ��r;�-�%w���7J�       �r4��_��_s�5N��544��{����^uuuV�)���S}}}N��l���V 8kܞ��]�:��9Yg*�ؤd�7��<�"(�ؤ⧎LYn�$�4N��<���&�#:�G����8g�}޼yz�'�������g�˥;�C_�җ�n�:�\S�����D��ϥ��/�� �rB����[��W;Wf��܎B9Sr��       PLS�?�njjR[[��0�x\�6mұc�rV��������|UUUY�W���i�e��y_��
(��+>�-�<w��Hƕ>��P���������rM�[?�~�_�>��>��hɒ%�φ���|������/~QW^y����z��w���ߨ�Pn� P�(���r]r�܎B��       (����e��X�48�4�k�.m۶M����n:��:v�R�T����|��3�Mͯ1��g�t<��5`=�~�rF"��P��;��U*2���`�2%�u�O߭��2��)�s8Z�v�~�wW�V����^����F=���z�'���2�y������+4�__-`:  J�vX%W%w��
%w       @9��i�񫮺��Ip.G��ƍ%�.C�Z�dR'N���|6�-�Wg:�&[0g�LňQp/\����d\��.���;(1֧tt"���}��\�{~>�yK�,��?�y=������yXoɒ%z��u�=�Ly�����w?�_�ɑ' �tPn��.��N�V��       (u�Y
����K-H�lFGG�~�z������[or�ȑ��WUU�u�����:٤)���z�2f:uz��t������$���7?�_����UVV����>��Ok�ܹ9Y���t��;����-^�x��;�]�>s��_{���  (��Q,.��N�ł�;       �T�&G>�#c���.��f� �,�Lj˖-:|������oR����
�>����k/�:S������}X�+���i�<|�o2f:���Q�4.j���a��u���iϻ�����/|A7�x#?��̜9s��O����<O�s����;����s�_�  ���(6�[r�܎bC�       P����B���_�l�i�f�w�֖-[TYY)��muL�4M����l>��%�+�i��T�3�%w�]�K��� (C����1�hN�3��GN�3�z}p׏u�o>�td|�s*++��CiժU���f���o�ҥK�����b���/+rr�����䬪/|P  f	��(V;�u��{�5�m���Q�Δ�둛�o      �0Ӕ�x��?���DT���i�$Ð���.ٜ.�+|rx���T���w�����c6�MK�,� $���W�������TSScu����ǵt�Ҝ���z5>��ޥih�1�	��l�lұ��Սy]֢���K��*5M��B�B�rTT����N��Ok�'|����ϟ�G}Ts���ET����F=��SZ�~�~��+�μ;t|�ϵ�s+��S?�o�5� ��QnG�;Wɝr;�%w       ��HD�*U*4*3�:�lrTV�Y�(W�9�e�M������3����U]]mA��611��۷���VuuuV��yS(RUUUN���|�wI����-��p^��(���R�#JN���܉ѓ��+e��Ν#4�W�7My��n��w߭u���n�x����v�[�N.Է��-���f��=����&]�+�R�uY� ��D���钻M���Ur�܎ق�;      ��aJ���Q*<&M����JG'��N(~�lN����r7̓�"7�O�Vb�W�SG3�ٽ����^z�%��v��i�����������:~I�!r�Ĕ�dL2��A��,
&�Tb�d��7MS�SG�yWf��Q��wN[n���z��'��w��r;��`�=��Ӻ�+�7Q����G_��I  ���mvx���-o���r;f�3%w�w      �F��V|��&lT���B[nϲF*���c�<���Gw(�v\�Ƀ�g_�pa����h����z�����:.B��r�\r�2��ֺym�3#���W7QF2����y.�����G�,��_��/^�X��Sαh�"}���բE��%���������ߟ���T��~W���Q��D� P$(�c�:SrRn�,E�      �l������z�޼3O�yx���w�H��(��6g��l6-X���4�e``@�ׯW4UMM��q�CCCJ���D�|�|��A�PC�7gkL��{isZ ��4ҧ��F� 륣�J�k=k<���t�O��f��t����{�e�v�7�ͦu�֩��]��ַ�3���%FNj��M�߂�  X�_�m�+1k���5��PnǬu���K�z�	�X       �e$"��أThԲ���R#�l]*wc�e9pZ�Ж����&UWW[��<D�Qm۶M^�W���V�A��i���-'�y�^��O�hu�ԓ��F����.A�%FO�.�7�P:��o�C��5u��S��9�N=��#S����e�]��~��jii�z|��F�����Q/  ��v�ri��	��S���      ��%Ǉ4������0�IEz�*|l��t��8eˈ��=c�����0mݺU�v�Ruu��Ց�9�'�L���*�V���5�c$)��2&ȫ�İR�1K֎���i�?������d�Yϫ���SO=�k����	Q��[��[Z�dI�����:�{�T|�H��           !�T��u���(�2y28��C[d�#VG)K��%3�(;o�<Ҕ���n=��sr�ݪ���:�hhh�^�N��J���ܬ��f9�ΌsZ���y1vp/mܑ7F"��X�215�H�y�74���5�9�����g>�K/����P�^�>��O�n�z<>|\�FE{�8           @�0M)���C�R��+-g��
umQ:2nu��9�j�񎎎')]���z�g�������J$��:�4��UWW��s��n?]Aζ��S)���Eg�6O:Ut7E!w(�#/L#����2��5=�L-۠{�����g=e���zꩧTWWW�p(�C?������Ǔ���[9����            �g�R��.%FOZ圌dB���J��VG)+��w�ͦ��vҔ�x<��^���jhh�͖��Q4L�����y�&����Bmmmr��g�Vp�����g�)3���w�Eb����8LSo��n_r�n�U�Vi���g��b�
}��Q*(�u��顇��!09qJ��p�"Y>�           �,�T�g�����̘i�:�]�X~w%���؝1���$��cA�ұg�m۶MUUUee�������J�d����֦����L5^o��� #E��TQpGΥ&���Xw����&�q�ܳ�|�A-X�@�t��7����\.��P�֬Y�G}T�#�X*4�C_�]Ѿ$           (��P׬ع���TB�#�d�VG)y��V�w�x[[�iJÑ#G�~�z�R)�|>���B�*���d2�9s模�a�s�^o��9��7S&��%��;r�Lƕ�l���/����d�;}���=�ܣ|�ǩ�+W��'>�	9�Όc�����?uԂd            ��
�*>x���HD���iu���푙ew�s�f9��ƍT__ou�@ 0�x<������d����*++�v2�|�~��2���^�(�#��#�e��%kw?��e�H����
��o�6�vX��+�ԯ�گe}�@2Я׿t�#',H           �f2�ȱWd��nxj��CG��Q��C]YǛ���d�J��ڲe���߯��Z�sxC,S,;k,�H��r���M3��f����2c���=�_rf��Kw�Lr|P�XȒ���7�%S?2�K.ѥ�^*�߯y��.�������c�e��=1zR����&�           �l��'#ˮܳQt�e}�r�^pg��ٳg�6oެ��Jy<���AI�o�H��jmmUmm����fnN�r''.*㹘��^�2ە�0Q%������y�|Fgg�:::������B!���*"��+��c�=�o~�2���z�]���N-�_�����    P����!U]~��1ސMj�
<���t�`�V�c��o�C��9J���3?Qh�+[��l6�ݴV��\#g�_����G��~�(�|�.���7�}�\3Si��z|�y�C�y_��Ш�O��y�n��?��myH4=O[�n�<m�J
������    �咓�J���i(ڻOU��:II�ugojj*p�٥��GPcc�jjj���"622���555Mٿ��l;�K�71��3_�f:)����	Jw\<�T|��L�8��9���{;&�qgFkkk��/^�H$�H$�������J=��#����-�-��
۩����~�����m    �]j��Q�w�ku��=*��ӡ����}=y]��vk���������[���5�����/}��E�l�5�Z��o����o{�7���/��o������|�:���y]#�R������h�g?��:_��x��_W�y�<�s��+6����j��'es��n���4�?�ѧ����1�     �;Ӕ������s��%��r��U<��Yvp���ȺS4�P(��[����V���V�A���z�jii��|S=%���XNV��4M�FJ6���'cV�5������|]gdX�5�P�7{����Y,�z��ph�ҥ}�p�V�Z�|0���S��?[�D    P�|K�k�w~(gͅ=^s�.y�3��g���#�|�sy]��l6-���g��%��p���ϩ���Zl�p���+�T�]�Y%��ko��m�
�^ۯ��:>��g��Ϙs�����`Y     @�J�d��V�ȋ����~�Tb�d�X]]�I��aںu���٣��z:q���Ą|>�֮]�ӛE**��8k�ɜ�13���(<
�(f2�dp��'º��j|YWWW���M�C���բE����5k���;��zl�?��S�~���    �tUt�S�c�������}����G���3oΥn�-����i��|�W�Ҵl6]��?���ou��Z>�XA�q7�U��?5�9�wݧ�kxL7     e�4�:Eޤ#JM[��$�c��v��=��sr��S�I���F�Z�z��,Y"I��b9���k]F�֘�iPp/E�qQc=2�����4��z[G�ǨTTT���U�G�pX}}}�z�9s��ښϴ���}�ݺ���zO~�S�8�\�   @�[{G����^+٧�������[��\�7�v�s�5��y����ݜ5���e��1�j|��r5���:����>Ņ�7��5���     �<�B�JG'���W�SǬ�PR�tR��ьq
�h����F����s�04>>�+��R7�p�Y;����3U�����0�q�R�R����|�?�Y7\֖����RGG�쿼�l����x�L&��ק��Q�oy����U[��G��b�����k�����tRG��A%�z-H    ��ݘ�ү��yF�y��-ù�4��yn������K������V�C��:��쿧�8�uf�    ��T���䈌d�vC.w��!)�ƫ555�)�HD6lЉ'T__ou�`0���f�r�-��|��P"���Z������tN���D��4����g��~����7ZI���������z����4Mhxx�����fӒ%K�v���	�ө_��_USSSƱ��)���e�r�    �Yb$�
��3y��L��[�_0g=o�߱�l���o 1SszdF��_�=9�z    �\�FZ���1
�T2�ou�����5SUUU�$��4Mm߾]�v�����:�X(����ڵk���9���=�ץ�ef93�L��{)������(p��ֻ��pd~��l6���O���7s�ݲ�l��АÐ���ҥKe����1�ϧ�\�B�/�矟�     ����_X��0|a��)��jhT�]�Y     ����Hٔ��CVG(��SY�˱���ݭ�7��p���ZE,�L*�����UW]5�פR�{�Zp�����Kw�7#Uj"���IƵ��!ue��---Y�1��%�á��a���R�^zi.����E�>�h�.����F_�gR   @i��������(C����݇��1�����Ħ     �B�Ш�
&�4�V�(	��X�����f���z�g������"f�����,Y�o��v�O&�9ˑ��^��4r�F6��&
�8o����    IDAT�@�L3���x�ŁMZvIs�cs��Qmm���p8�r�46v�C���เ\���+u�m�e=v�[�)6X��   �E���(X%`��?б/=mu�s�.Z��U�:     (c�Tp�i(����������C�=�Hh�ƍ:|���n�	���ب[o���n��w���p�i�s�Fv��0�V��b�BJE�����n_Z��Xuu�s������Pgg�~�����Immm9����w�N�8�C��5n��:�W��/�$�c�w�   @��>���;�N*T�W�����e�}=
����op���
4��kb��VǙ���>��X     �!�4��NZ��R�q9�s�g*g��R߼tϞ=��_Q�Ѩ�n�n��f����u*���&�#�x*���2g�d0�C<�A��%1�[����I��yD�7���VKKK��t�\�뮻���\����:;;�hѢ�����n��?�q�����&&&�:>�S?�C�����   ��i�������^����O�c�zuknS�����:
     (3f""��U<4�a�#��t��
�ǏWWW�����b�z\�T*�h4�뮻N���K��9HuڔE�TTr����3��;f,(]�`�$���&s�v�ݮ���)���X���Z�b�v�ء��	mذA�������/�n'�|��������/�R�y�����j�X����Z�  L綛���5�Y���>6���.�c �V\q����S������j��������VG����4�C������$     �̤�؅��M��8��T7
�\�'ɯ��I�رC��ժ���:�\ �W\��������N�Ř�ϙ��l�lr�g@�(Ѫr�4��tɆ��Zyyf�]�Z[[sr��T�Ѩ:�ƿ��~�R)mڴI>�OW_}u����[-_�\7�|�6n�xָ�N��7?�˾����� ���m�O��◫���u�ظ�!�c ���A����֍�����=�+��fu (���>�����R���     
�H%��PpF:nu��0Ս���{:��֭[e��U[[ku���	�����xG��6��=ec�N��L�l����I!墴�P#o���2�����tGG,뱺�:UWW�m�x<�6hbb"�Xmm��N�^z�%���KJ$��C8�q������-c<6إ�~ނD  `&lfB�A%����B:rl\�ÃV�@���	(.�_
������B ��^Q���}��     �ܤ�V'(83]B�,d�㥰)��ݻ�y�fUVV�u�W�~�hT�DBk֬ѢE��F.�6[�ͥ�<W����$Qpǹ�����XV�v��_�1��xr�x��J&�ڸq����w��z��x<ڱc�6mڤ��ɼe�ӏW���>��C��/�B��-H  f��J���T	��)�(w-��l��z�3     (nS��KwL���O�<���jj2�q��ah||\o��u�u�MY�� �p{��&��Jw�SjrDf�l
�����2��v������f�N��i�&�����5���־}��a�����% IZ�n]��Љ�DA�O ��)��;��2W%w��  �綨��wY      8�)
��(��Z(҆��ק������Autt�[n���:N�̾�[X��;�g�JNl9[*����כ3gN^ɲm�6]؟��v����رcz��gu����N�뮻��֖19�WC�� ����%w��4�K��࿵|�1�#     �2b�g>���ٝV'(i���n��o߮ݻw�����(���X(����ڵk5w�܂������i>����E���=�C��J��d$�[o���j�We�{�^��e��+�����=z����v����ԩSڸq����r��oN�S��G�~���/*>|̂T  `�fcɽ�r;�l��)�(F<�����έ��jU]��<'     8��(��w9���cv��~��mܸQ�C���V�AK$�����u��|��J鹔J��@K�(�WŴ��۽�3qR7-�e���v���������ڻwoN��l�����Ą6lؠ={��0fO��K.�M7ݔ1n$"���,H  ��l*�w�(�v��-����Qr���\������������;     (��cu���;�VG(	Su�R���622�g�}V�h4��b�3C�@@˖-���_�ӝ��G.ם�#��{U��KwL)�HD����.yܙ𚚚��2��`P/��r^�����J�Rڴi��o߮t��FBY���T[[�1��#M�{ւD  �|̆�;�vLǦ�/�PnPf����2�3{c��-ω      ${E��
��)�?s>��ެ�����b��6mڤ��n��8�`0���f�z�Y;`��ˍ��*��\9[#��6�Х��`J��Y�&芅���
���㹐H$����쮾3?�^z�%�l6]}�ժ���7JWEE���~}����8��/�S���.��  �3%���\E�73�혉3%w�N>_q}�8�	�� �LrlT#?�w5���9ϵ9�j���t�+P�d@��������V�(:��%t+��5��    �n�d�Iy�|���ʰԟ����D��I�g��^y���aUWg��
�TUU��k�Z�Ng�.VO��oڞ�y䰤��Qd5
#��h��n�K��p7w�ܜ�!t�i�ںu�&''s>��x���.|�W�J��b�
>����Z�J�7o֑#G���ح���W̢d  `����N��K��1[��,�l��K-[�5��o������xX}��s�#�$���;.�:F���/��� w    ��f���Z���I
�9E1��Q����b����ѣ:v��~�|>��qPĒɤb�����w��rY�,��3��3�Sp/I�q�E'9q�`k�w��1��^__���ʼ�y��A����e��x<��|ڿ�6nܨ��aK�`���lz��ߟ�&���NF,dA*  p�Δܓ�y�д(�����y|\w}7��Yf�l�h�-���N�-q'v��(&fI(�r�@��<t��-�>�mo������BC
-YL 	du��Ypb�K�}��e$͌f_���a$��(I����|ޯ�^������4��9����t���S��'�*��v�&��m��cN����^ע%_�*#}�(F��R�\��G�oo7�""sI--V�0kI>��%��=A�K�A��i����0Q�=��V��b�HO=�"��.�f1]�122��K�bӦM�.����=��C���е�_U*����XE��6�d��eYF(2e�H$�����r���l���8s��y�˃�T],X�5k��b}x����""""���r?�p;��l�3�N�E����&�"Z�}��bJh�~W�s3gNM>�f����-{n�ݟD�"&"""""""s�s2@���@gɶ�UN��~2i]��B��ݻw�رc�B%�R�����M7݄@ `u922t�(��� �[�$Q2��d	�4�"Jb�^�@���h�(�$
� I�?騪�W^ye­0�$I���000��Ǐc�ܹ��겺,�۶m�����^ �����[���ݚ���������������1<�p;��h�]���*��F38��v��c���_BtN�+]�w���߀^���$��[?X����������"��F��)8�/�t�s�Bn�	�短@eDDDDDDDT�do�(A�*s�J6w3�Dy�D"Q�J.ٿ?��(|�5�&��d`�۱i�&�U�`�Ȁ{�P(K�T@6�fAb��J��:
���,%k9l�S>���mݲw�^�b��N?]� ����D�=�����b�
��G
�����s��q�JrO}��u�*#""������t=_�u��b��� }�1
�=���ۀ
ݨM45��ӿ@��t�����nD���*P�}[Y�{ ?� W�J�п�0��������<�DDDDDDDd*A� ��P�^���	��X]DͰ��J�W����p��1���=)��T*�6��*�\�l�p8;V�nzRY���������c���h̰8s �g�xKK�)a���~�8q������#���^��={fe�y��n�
��x+��_��TԂ��������W��e�m�~���Lo-]U0���&WCf
?���xYs��� w��&WDDDDDDDD���t��%�N�4A�g�hz��%�+��}ddO=����*�&U�x<�ছn��p�$I�e���:��Tɰ�OD��1�N�(��to�,և��R644�������سg�*�<��z!Iv�ލݻw#��Y]�2>�7�xcѸ���Sߴ�""""""���Udϝ.kn�[`on5�"�}�*���,kn����0�"2��JN�F��O~��j�������� ���ᶺS9��[]BM�����`l,3u]UU�{�n���[�BEF,ib�xn��7oFKK���L��i�M9����g4���Ā{-�/�ѕ<�Le�p�ߋ���N�P(d�zD<^^ת���v��ra�޽x���k�s"�lݺ�䋎�'�	-[�홈�����ꚮ#��CeM$Ϳ��䂀֏~��?hb%T)}��tU-kn�w�l6�""""""""�o���.�4��[c��e�A� ��ÑHĴ5�z�-���Kp�\����r9��y�p����i3��<�ϗl@�(�Sf��Ā;�QR���'A�c]0[4�r��v�f4ő#G?���^/>�]�vahh��h�x<ظqcѸ��a���YPQ�
��!�Jq��RZ��j�.o�PYs��}y��j����� �ܓe��v�~�S&WDDDDDDDD���4���!f-p�u0�_��:�Ɔ��_���O=�r��^��ǧڡiFFFp�WbÆ���]����\.Wr<V���;��$�i���L��#�6�C�E�fto�u���:4M3�س��f���Ù3g����V�D���!��?���tU��""""""��T
#��β�:;�÷n�i��n�m�>YsÏ<Xv�o����mw~��ab5DDDDDDDT��9�[]��dw ��v�˨I��eEc�\�Tʐ�'�I�ܹ===�dר��b1̙37�t�.�F6$�(��̽iDbu�h@�1�N  -����Td�k��1��	��c�Z�ΝC86����(����>��Ǐ[]Y���k׮-��El�cTDDDDDDT��({n���L����ck�?~ȴ:��⯿���e͵Cew�'"""""""�.��6��eF��4u��z�l[Rr|hhhF�UU���
�|�M466V}n2W2������-[��^[7���f�Ec��#��F)���-��wP���ɓ��T��ESS��k���7�|����f�   �H`�Ν8p�@�v����r�-J�����?XPQ������޲�6��v����fʵh	�W�]J�����1��V���+{n��~�c��������t�9+ �6��0��u1$���2j�D����i�ȑ#صkG�t�&s��yd2lܸ+V���S��d�,'I�6��(E�1�^�p' ��/��ɲ���zo���a��T���F(��_|o����u���˖-+O�~�S���""""""����*����B���5�~�Se�?\~�y�C�������6t-�o��+"""""""�z'�]h�����%O��.�˨i��N'�>88���~�T
�@`��Q�4�h��ݸ���!���u�\��^P*�>���ݰ5JL>>YG�� ���M@W��#�øb��h<��6=�l�6������ v��Q�v�Z8��]���lڴ��c`p׽p/�ڂ��������5�r;��oН�Bt��0�^Gl�.�iko~xd.����2N��~���ໆ�-��h.34_D乧[�(���êG����k�RG�B��C��)+��R�����/�����=���brUDDDDDDDT�l�V8[!;P��l���W�y����}}�5t �\.��_~�F�F5*�a���X�n�ե���.�r�D���@J�߼vAf�Zŀ;AME+�����m�qc� �rG��o�EQ?n5���o�>
\u�U�tΧ�a�ʕ�7>��1��߀��ZT�o8�/���2S����߃�͠�?����oPSIS֙L��<F~�2�6N:��k<��B���������!�ʚ;��AW�o�0U����U3:�w��h�����_|C?Ԡʪ��C��e��2�2�6����9S����)n��I�ij�\j�~w�$"""""������
9�#=V�2%�(ó�j�66�4�����-;��n9w]ױo�>�R)��~�J��J�����e��K�#�����P(��0�L��6�kUm�@S��GL_C�5�i)�z��ns\��ĉ���8x<>|�=�����.�L �"�����q-�D�ZPQ�N�|�+X��g�Zl�V��Gv�=�去[�e{��
��!�֝�D�������]�
�a=���&���]s"2�8�F��͓��Ϳ�K?����lg�"""""�YC�й
6o��J�&�"܋�Ar��dE\Ż���a���	?�ԩSx�g ߥ�j��(H$��kp�WZ]NEy�G2Y��P��\��:��3Д��%�>����h܌��ؽ�<6�~�gΜ�Ν;q���K"�]�������������8;�c��{�
K�~�q(�HYsC�����T9�΃��e͍��*2�j�Y� ���fu����w ]/kn�C�����g���!w"""""��D�^����+�� ��^|dO��R�J���Ec����:E"<��3�F��u���F��ՅM�6�n�[]NEI�d���T�Ή��#io3l����{�b��Ω�XE�Y,\,�e��;�ؽ}�DQDcc#��0v�܉cǎY]������//O�|��,��������:�ׇ�o�[��s&���Ѳ�Jn��������������z�·f=D���2,�>q#��.k���F�G�4�""k�67Z�nP�s$U�(�a�j8B�dB��	�k!���.���)9~��ٱ�
�޽ǎCSS�2ύR}����z�����.�^����I������N��(E���t���.����GL_C(�����'��o���cǎAUUC�YO�L&�s�N�B!�\��dp��\s*��� �|��-��������:���������劯~�A��se�m����IF�oo/k���ӿ��ZUG!��в�+�D�}�¿acYs�~���^�*wJ��K6O������-{W3�=��'Dqj�5�+��	�+`艃3/��������p�]	�@��!�����Ȟ毆h��ϳ�D���� ��ߏh4
��Wɲ�
e2��v�x�u��������T��7���>o���lhS/p�c��@�oa������Y4n����(��n���F(��_|X�z5d�O��+�@CC�����ȯƜ��]���������jE������WdN���G�<�&<���t���pw_��ѷ��V�[`on-k��������L@�E�.�2��A��)�,�t��c�nފ��@eD�$�ЧR�dcw�.�+A Ʌ��w�!Jv�6A��<�ln�>�MӴKT���DDDDDD�ao������P�1KkD	��.8[2_a!לdt%7n��ɓx�g����p;�'EQ��fq��W��,�1�##;׫��L��:CoJ��-S�ho0w��u�R/�\1 �qcv����uN�>�\.7�D*��{�'̫��
Q�f����26�k֬�K/�4n<>�ԙ7�^�΢ʈ�����,"�m� .��?V|��#;�
�@�G>���~mZ�n�������֨V�O=��w��u�?�=,��ߖ5��ӿǀ;U]׫v�q�f���'�X�� �Z �.������q�MH�    IDAT�P(�&�NDuiGؗ���;DD�&	�' ^Q@�l��U��F��#9��.���Ed.���+^���
ל���َ��+�:�Ƹ�!�hR�X+V�@kkyMa��f�!�H�lB�W0�����st-c����ل�kHJ��)��n�]s����ѣ��~�����}��!��c��ռ󱊬]��(�\��΀;�#��7Xpz�ǘ��	��tn���?��lvJk�����Ʋ�&��ԑ��t�j����{�˰\��`��	d�s�W����H�W�ʈ�OQȲ\�!w�͉�{<�����ݰ���c��~[m"��[i;.�F"�	� ���Ӂ.�p��訾אD�C��il�V�O#7t�Rz�+#���m]�=M��E�s/��(� }}}X�h��
����q���c͚5V�2�ٽ FFF��EA��f��m.�W +�gS3���R���Ga�@ ��Op���p8��zq��a�ܹ���V�De���*�����0�-�����������2K�U�)?����>?�n~���h��.�T���#N���*}�j�V�b9-�F���w�o���L�������UlvTeꝖ%�>��B����~�MN�uds9�G���?�?=Ʀ3Q|f��]�oMDed��K�[���.��`|CFA��h�o���,����Y��]��G___�+��.��!����n@ww����JMM�>Ǖ�m�:wb�|C�y7A� ���A�b�:�r�U�Ozϓ� �B��l�os��	C�G��f����gϞŁ��Յ��N�ˢ	���U�V��_7���ԙ7�ŝ�����w�o"�莊�k�`�?���l��v'���#;��O�5�e�]z���\Ѽ��eM�2i����"ٳ�0����x5�@��!���"tU1�����w����A�&?=����ǿF�����Yv@Q ��}'A�������ʼ���j��DDӗ��ql(��<�9��z�i�f!A��hY G���
#}($�����>��A��6O��6_�5���m���co/�Y�%��!�Lb���p��V�3k��hh�]�u$ō��' x�}^������uJ͚߽�4�[���F� ��r�pႡǤ򈢈@ ���A�8qs��EWW��eQ	W]uUQ� F���w"""""2\��������S��ׂu�o����chX�tҹ����9o!��N�u����pt�)k��/������J�8����7V�Qsr�=�<�$���>�\A�������?�m*#�?6�JajwA� ��g��i��)�ۉ���L��X:���Nlj��k^��EQI���关�5Z&5���MA�g�kʥf�
H6�Qr@t4@rz :=�FV���e�#��ָ�X,�t:��~=�Y,CWW�Νku)�^SS����T�xw�~�o�m.�� k1�^��l��5|ѣ�^V������Ι3gJ>IRe566"�H��C0�ʕ+!���Ycٲep8��r��c�@Ƕ���*"""""��~�����s򉂀�;�,;�ݲ�������eϥ��w߽e����BϷ�-�6�*��#�P�<��O>  J�ax]/�����ܓҰ�wx,�.�ϟ�n�DD��i4M��������r�f�H�����~\&���Y�v7�����Q���h�Q��@r[�k#U�o�梀;p����ŋ-����L&�e��K��P���E�Ѣ1EQ0d�f'E��9T�}p�SZ:�w�" ƿx��jgΜ1�x43~�����^�����ի!�|���,����¡C�ƍ�N��B<��Ţʈ��������O~�ί�9D���z[�}����+���g6#����O�8�ā�eͥڕ��+$�	Ϫ�&�+��h��v<��
TFT_DQ�(J�t�P^�eQ��1�NT��֋��.Dcc�ŕU�|>�x<�D"�X,Vr'�D*��Kg�H0�{�v8ʾ%�����]v#��������p�3�B�B6l�����t�(�hjj2���X�h�ȉ�[>f�:�H��<�W�C����L|7�Q���7�r�\�v�N&�6�xd��I��ꫯb����d2V�T�V�XQ<�k���l�!"""""�cJ,���'˚k6#���&���C�����{;���e�������Gd
��	M/��%J�?�v�%�e��4�8�p;���v�B!,X� �V�������z��麎�C|�Bo����DDd2��7C���̽��TCV�u�x˗/�ƍn��`0I�;��(H$�-�J� ��sɢ�	��sdT�xE��٤�k�2��,�+ohh0t��g�z<2^CC\.�|�M<�����V�T�J��x��tM��A>ڃl�Q��B��>�N����ב>����;�B�"�t��Z]6�Z��e�m���� h��'�:���c�珖�6ն�_������:�/B`�f�+"�O���T�%:���(���r%�U�J븟�ۉ�%I�� ������]�95�N����ty����?�K7������Rm��b�Bؼy3|��\"M������E"���
���uJ�\�7&R푭.�*O˧M_�)u�X|����s��z<2�������#G�J��b�
���X]V]	�BhiiA87{�E�T)�(��(��K���n=-��ݍ�=!������JDDDDD���������9ҹ����蘃\oO������y�Z7���P����J5LW
��}��������w�x��h6���@.���8A�}�犈��ܓҰ�����r���z�����z�����za��!< @�e8�������z�(ʸ�������P�P@>�G:�F:�F*�B*�B:�F2�7FT/�n7-Z�L&����#��MAEU�_=Cw4�/<�;���W�d��ܹs6~��N��p8�e��K�jN���������z���o���ė&:<&�@��uH�g&�4C����qc� ��r�F"�@45�xT�,����ܹs8x� ������iuYucɒ%E�B���Sp�.��*z/��Cn�<�h��@�5(��d��㐜؛���Xb/"""""2��c�c����sE��>���ǒ�n��ɲ�?�`�s�>���O\�{_�������Ѱt9��W�2��a�9���_���l>o�1���8D��[i�����x��ڊ��V�������@`,�>����޻vTJ�P@4E${�F�F4������P(�.��0.�K�.���0zzz�(
�K7��b�������[`͇p����wo�v��y�k�荚6l����������n�C�k~�}vp��סJtp_�-��t:!��ak���v,�<Q088��Ǐc�ܹX�t��eռ%K���_.O�̀�,��3��F~�t͜��l�ޣ���=0ζ%�NS�"""""�b�Gw`Η��4��֏܉���tU7.7�t�e���p#{^�V�T����(Z?Zލ��,N}��L����Ȳ���ؿUUC.W &�N7Qw"�]��^}DQD[[�̙����qa�����n�K���6V�Dt]���0z{{��ׇ��^�������f+X1�q�� �~?Μ9�x<>6�R��Jh�_���@���yh��
��ƍ���"���n�M� �bժU�����'Z[['�8�h껮W ����uJmϏ��댮䡫��k�^�]�\4nd�v �x��#�$�I�ڵn��֭� pK73,Y���x���m����P)��!7p��I��`{MC~�
�p�,��m1 �d�Ut]�^�_�4�B?s�.���|����z�Dd�|F^~�7�4�\{{��ވ�Kύo��v�ev�	?�@Qg#" ��^�n�(�|L�C�q�_����
TFTlv'UA��lD����=)�3�>���n̛7��������ŋ�`�8�3o(��*TU��(Pe�ߚ�A�u�~}��긿�~AƮ�	�0�)�$IE�$�����R7�
��P(�P(�U�V�?���ɓ�p�Ο?��'O���g�{�h6�eK�,A__����[O��Yn��Jo�CDD&i\󡢀��i�p�-bs�j622���N�Y���RjJss��7�"�|��W�%���iv`���h���k4�K��0�$�(UU�;�>ߥ>�w�����ի!�|�2R(B (�"&y���;U��B�����Q��i��G>z��U�<AK� "�g��������.�mA/�ifr��>\�c��l��m͐�ʮKd��#;�
�@��;��-��*�cuU��cO�>���0���_{�sE����|�+PQ}�e;���K6��C@�N��C�DT���� ��Jkk+����p�B̟?���GSSӔ��(
��<
������G죡v}�ܠ*dY��f+���n��n�ݼ����~�z�_�~l,���ܹs8{�,N�8��G�2�N�Z{{;\.Μ93v��.begl�FDT)M>�ޟ��E�N�b��Je�Y���͛7�)�	�̙c��4M���p���Sa��]��e~�x���3�M61 �O"Fvp���ۉ����p���^{��`ݺuU�U�l�p�B�ݻw�X����0d�-��@��8��' X�Z˥�<�*�]p�/&��JDDƺn?j�ڙL��`ȝf$W���`��� PP���dȝ�Rd�(�aM��jӖ���ZP�tӿ��uhX���u���A>�?�Z����woYw h��w�����˙\Q}�ٜP
9 �Ρ��I.%vo'���4��-&�"�̙��˗����������#��#��!�ˍ�����p뺎B��Bίl��l���p8�����%��\.tww���[�np)�~��Y>|�Ƒ#G�H$L�������]]]8y�䥝4�Ǐ;}�1�GDT��eh����ƍ_�p�|��N�dMӐH$p�5׌���X������Kf7O��_�)A!����C��u�ܛ�4�p�$����f�ћ"8�T*��k�"X\U��7o^Q�����7�[q�5E�1]U�:��D��=V�u �J:��5�FDd���r���2�>�!w�V��`𧏠�_�t� �h�����  ��d��yp�5R}�����'�Z�xҹ�`�[?���~T�ʈj�$����as�! Г
�_���$$������JD�;�[��v���˖-òe����U�ժ�"��"�� ��"��!��T]���!�T*U�>����	��������Qԡ��r�}>�@�4������Ɓp��A��rn�K�,���ǡ�*��,�0��DD������8w��,YbQU4�X�_~9��ڬ.��ݽ ��Ν?�l����%�&�9�j�uF+dM^@A������p�L86�x4�98�8q�x˗/GGG��eU�y��O��π{�i�<R�^���[]ʄ�x�����j�2O��a$�����Q��t̆p�(�ܩZ<� :~��@��Z�߅��}�ǋ���u�|b/�i�T�t�~��weMo���p'2��9�+����v�B�����M?��	;�W�(�X�p!���
\u�UX�bE�.����J���f��&�jN�����NEN�N�.�n��(�.�":;;��ى[o� ��ߏ������طo�i�w1'z���,Z�'N����8;�O+����DD��.�<�����]�O�:ŀ�,����ֆ5k�X]J��z��7�-
�F�E�.$ /i2t�R��䓨f0�^g��k�gѲ,X4nd�vUU�D;UI���ۋ#G�`���X�h��eU�y��A�>n<}�E�']�!y�h��.&���A�ī�,� �!w""Cͦp�(��i*riք�G1�N�({��{��k&�뜿��Wõ����-[Ï�>��4{�}s���������W·nC�"�/��"�N�� d��⊈���Ii���vS566⪫��ڵkq�W���M8W�ud2�R)�R)d2��	�� Q��PӴ�kCV�4�tz\@]�������BCCdy|����[�n�֭[Q(p��Q�ݻ��կ���S�O��������q�� ���ql��m�=ֈ�j���
��[0r�q�===H��hh(��)UN>������&����1Qԙ(ڭJUU��b�>3ǀ{}a����j�nn@ůC����DfUx�*O466"�a׮]hkkòeˬ.�j�\.�A�O��oQE�GW$O��*���l�S��r/�<ODDS7��r�r\
�����1�N�(�Ȏ�� �r�]hX�]ށ5�?4�ʨ�h��@�g�T����?�̩�&WET_ҩ�� Y� �N���ꒈ�B���ٹ��(���k֬��5k�hѢ���(EQ��֣��w7̮U�$H�Y���|��EQ�s��xg��ܠ���c���i�4��BUՒ/
Pe�O3�_TUE2�D2�s8p���z�p����6�+W��ʕ+��O���x�װg�9r��_C�OMMMH�R��Hg2�������+x���������+-���M�4$�I�]�^���r���3�{;p)��n{�̿���Mr�!H<WVO�P�#fwo�&1	��D����ʥ�����N��k�.��n�Y��w������豔�=���`3�*��:R�_���[]ʔ�����g�:�"�]ծ�����bȝ��l��bȝ���?ǂ��Hމ;H�
��aRy��b�����3-��H�������A�'�P�t�-��.�D�"���a�fg���^ܓ�n7�(�����ƍq�ע����<]בN��L&�Ǒ�dL�K�$�l6���qo�c���%��z�YWU�q��|>?�����t������v�v�\�x<p���x<�nZ�����m۰m�6��q�ٳ{���޽{�����hԜ9s�L&�N���pI_ ��҈��ִ�\x�Q�=v��D,Ò%K�n�:�K�;���7��###�v_u �p�q�Љ�{{�a���hJ�r�5���N�n�[H����E�֭3���ִ���СC��tUA��(:�������;%9luӦ�������m�եU����C�gw�}C�TJ5��G1�N�D�f0������OO:��p; �����z���C��'����'�"�~�V�"�:�~xܗ.��Ճ{R�g��������p�M7�����B�0hO�RP��A��n���{����x��4?ѵ8M�����<��,�٬!�2�2�!��z��������p��7��oF>�Ǟ={�k�.�۷��=�7A�`�>|�B���~܉��&�v�n�,�~���A__���-����$� �l�bu)u���~��a𾾾�c���0?����7/S�ߢiR����(ߍ?�U�Q�ѨaǢ��v� ���:E��u����7&z�8ɀ���� r��.c�r��!{�|�HD4�nŐ;�S5��G1�N�d��e�˥D#��zڰ�Q����w��euz'��S#P��7$��沺$"2ٷ�:;���h�}���%�}�viO$H$�vi�ey\���r��p��&^�DQ�y�Ѱ{&���rӿ���:R�R����a�������z�v�!�����n���_�믿�d���:v�ލ7�xc�1H4N�mmm���Þh���w���|-[���_�tu��ko��6�(
(
���ka��A��E�?n.����P���G{a��v��{7��`c��zÀ{���\�T45��f���N̔������j��u��ϡC����r�J���=&�\���p%�C�T���[]ʌ麎���-�x����\�nŐ;�nŐ;U����:|��+9^�'A˛|>�jR��ב<��+V[]
Q]����A�]A��!"�ݓ�n��P(����}ؼy��;��$FFF022bH�nQ��� ���������4��v����ݙ�K�3���4R�2�
���j������� dY������������`���'iڸ    IDATؼy3�����/`�Ν8��!�#կ��6D"ds9<�����DD��������ظ�g�"�L���XTY}�u�Xk֬a>�b���hhh0��������\.�Ӷ%��oFl�Y�p�#�bnw%և���'�'ښn:��8)��l��l8q���8�/_����˲\sss��lt��r�ǡ��V�a-�Bv��mK�.���*�$Q���Q�׷j��b��x��W½l�T
�SǑ:���%Մ�;�`��t�r�O}���\�-�� ���G<F��A`w�Q-�'��~�ۧDE�\�[�nņ I�M�R��X�}���Q6�m,��v��t:k�E�DQ����U(�J��N��N���d�5�Q�h�h�(��󡱱^�w���m�6l۶'O��SO=�^x��n�T?DQDGGΜ9�_$r���.�DD���[�_p�4�����-��~�b1,\�k׮����'�2�͛g�qUUE����z���3|�w��7N�#�눮��D�dl�a����q�Á\.gH�}ddd�Ǡ�$I� .^��C�a��Ŧl�R-�^��c��g,���i��5�?7p��\���-F���7.�ۏX]�!ƅܥ�ߕ��s)�~����r7���c�7�A�u�ƍgN���O��#;�D#�W�(�����9�6o�7^C��	���z4���1{�r&�����d	v����Ȯ�D����:`��l�`�6m�m��V�yO:����b�،B���g,d���ֳ�lhll{lh��d29���f�t<M����� ��X���]]/^�ŋ�3��^|�E�ڵ�6�����ۋ�x�f'�ϣ��w���D�¡q�G���ի!ˌH�!�J���`˖-V�B��`�S������v�RU��A�|I.?���zįz�ՙo��^<H(�766���###H&�3
�'�THt��P(�X,��;w"
�+���,K����avp7C��$0Ů"�@�4�§�l�ե�Z�n5r�&�LU�7�vs���w��i�������5E�s-\��?����?���E��eW�iPq?�4��'���*�z�+������?������
"C��^����j��""2�=)���2Ȳ�6��[n�ʕ+!���
D"D"�i��EQ�������-�ċf���>ߥsR�ޓ�$�Ĕ�E��8���444`�֭غu+N�>�'�x�v�*jET� hkkùs��H��}����'h�������9n8����ѣX�b�E��&EQ��dp���u�,������f�qu]GOOO��+{�B����J�<��^1�^/t�fnw:�(p���~��~$	��q���)o�J��(����/E��]��v��f͚�[Z֪`0Xp��t�	>��J+d��\������Ѻ��-������5���~�� ����օH���<y0- ���j�ȝ%���$:h��N��q'⯿�������'���. �~dǌ�j"��'n`ET��>�|�Ct5X]
QM
��(
p9��}�m|�բ{R�g��=��~�v�m���[��_t]G2�D$A<�>��2v��>���(8O������<��8���d��#�B������B0Dcc��������������O������i�Ն`0��/�tw;k�����t�G����D��������cٲeu�2S4ŪU����gQ�x�bS���ׇ|>?nL�4��@\d�9,A� 7�M_�f'����f~�=��P�����G;!d2D�QȲ\�	$����^y���v\u�Uuq�aSSq�NWP��ސզ���K7�(]SQ� G�9/����ّc�w�U��=a�K�Y(x��S��[��u�뻈����_<�\�Ś���H�=� s�$\��:{�g�B�f���2���E�G��R�j�R�#2t��@ �n�;m���=��s�{hoo�>���}�+������D�F�ܭ]��@����f3�l�e�v;B�B�EA<G<G2�{�M&�ɠ��}}}���hjjBCåЎ���w܁m۶�7���~�38p��O��� ��NM��!"��(�����������4�;��˹3�L��qttt`͚�n�C֘;w���V#麎���z�ݷ��������1��^���Z���].\.r����!IҤw�%���I4���{�쁢(X�n�n��U�����/���E�Q��n��Q�H�DDDDu���1��s�_��?�:��kвYhys�痻S��˚����!:��/����Gw\�u���c��~ductEA~�������������G��OS܉���3�{6Y��i���l���D��;)���	�X�����v��qͰt]���"�Ȕ�
� �ۍ��F�|>�2/��#Y���Ԅ��&h��d2�����q�e�.��*"�"��N'�� � DQ�(�X�~=֯_�cǎ�?�)^~��C�T?���prx:<�oSDD���)�>����7~��twws�i�f���lشiS��ߩ�<�Νkʱ����͎���i^� wV&[�[}�o�u��BqׄrB��PCCC 0�ɦt:=�B�&�r�  D&��W\�`0hqU��xJwP��e.�F)��|�wMT�I���^�!"""�uJ,`ь�!:��Nc
�������#��C���B���e2���2��ʳC�_{��ei�~"�>����9s
���G����.���S#@s�\�v�K""�ݓ�p?��㈢��k�b��������B��H$���a(�Ԯmz<��~vj�"�(�u��4�D�h�����l/^D?�� ������ҥK�կ~���~�'�xb�;P��x<%	��d�dGDT	�dC�m�s���q�D�Ɗ+,�����n��kL�N�E��ݦ�|�i.\�P4��k{�,�XE��r�����Id-ޖT'*����(�O�+�,�hkkCKKt]/��P(�uG=�Q�v;�~?N�:�g�}��+�l��?�Q-
#��Y	[]U@��3ǏZ]¤
Ã�>��?.���&TC�4�|+��?[]FE��w��%�]���s�'d��3IvY]�;��#�2�����;���������r9����رc(;��v���сe˖a���D����ߏ���cٲe�;w.�^oY� UU�q��Q�;w�Tj�}������>�{���vۄ;�S��z�x��p;Q%5o�<��MZ��ۇ|>oAE�'�a�ܹ�馛n��-Z4���h/^D.7~7^UU�'�XWu��\�uh�b��^h����N�9�$�"������Aƞ(���IT)�$!����v�3g�.�ܕ8��FQCV�P1���%Q���Oh5p ��i�K(K��S��e���OL��J	��a�������^څ̩V�ATS�@Ur�z]	NO��%���=��>��\��r�M7�[�����/���u�}�dgϞűc��D��m����҂��n,Z��P��v����,@ww7����p8&�8]�122�S�N��ɓ��b��K���f|�_����=|�����6�ӠY����ta��6""2� �qٶ�*�f�8x�U�d2	�ݎ-[������rh�`д�S�P(ٽ}����?dʚ�&�vH._Eً֢�:������.q'�T:��� ����`��0222��fL�|>D"�ܹ�����>%�p%�IWP3	�˨5�^��������Z�S'p�-����i���!��/�.�,���C�����C��)�d��2[�7l����:����UՌl&���94��.OD�;Q%ܓ���š�����͛7����6�򕯠��}�}�x'O���ӧ���:���ży���ݍ��6v�&C�l6477c�ҥX�d	��� ��G)��4Ο?��G�bh�7�{�ߏ;���{/�㎲��T�<R;�UZ��;�^��h�����va�Kr�r����z�\Y��<j���DWW�i�?�<Tu|(��a_��;`ں�$���2vZ��ƀ{�����IW�p:��#�$��N~�����ewp 2Scc#E��]��gϞ���`��iZ>S�Jjӥp{���5hYi�������ӏ��[����ʠ���;h٬�e�EWU��a���?hb54�Sz�4#h��v4�+����c?�23}�Z�i*.�=���]��f�Σ�*����ս�˖-o���YH�&x�8�0ӡ��0m�tZh�0-eZ�k��)���R([�-K��,M e	�AI��Ļ�ݱ-o�����8��%��%�_�pN�ܫ�|�؊|���<�l�ΐ�vYD%���)޹]TUU��{�ŵ�^;lW===8p� 122���,��tb���(**��f���Ř�`@~~>�ϟ���\���)_�����ֆ���	Aw�ło~����~�/���� �N��EDw�����"l8`���*47�B!���a�8��3��h�.��AE,X� j��������=l��-�@���y"A!�q���6�SE�;����4���}�� \.֭[�y����v#D��D�a�Z��h��{���w�����<��u7a�=:B����r�3Q��u�������%������R��i�~�t��Y�˘���� %����{1�kG*�y�bvmw7��CS��i��YcB�t>�T��!Jvm-�!AX,`� =%�ߌ(x2���K�,�=�܃n�EEE ��{{{q��A���������j���Bee%�N'C��
�F�Á��r���"--m��ݻ���d�l6\z���o~���??���i���(|FDD'g]�������CKK�
�-���p:�8��sa���.�f���&�)fׯ���rB3���n�מQk�ټǓ��4�E���Xwp�{#�\��ʮ��8���Q]]���
&T�����d��`��;�u�V��p�d'B����8���z�]Qr	����c��p���o�߁9����W�u7�H�2fl��eZ�ٛ�=�Љn���z̮��8���Ny^��Y���ãP�l8A4[G��1<x�4 s4��������O���l����w�un��6��� 8�\���5558r�Ȕ�vQ������J�\.X�Vvk�9�h4��� �����ʚ�[���GGG�x�}�!++W]u��^,[�,��`�"""��_|GĐ�m�������cY��kע��@�jh�rss�t:cv���n������a:����{<A �b�5Rb�2�� ��P0b�=���C����a����x<�裏�(
����"�D��C��c߾}��ŋa���.+�I;���q�$9����&�f""""�?���w�B��oA?�ί~�_�
���+C�3�#ލ�G�'� b���_���*+D<���c���8WEP��|�N�|�F��Z]n~���o���8�}�m�}�d���2Q2�EwG���E��
�1S�(
~;����gdd��.�9�3!��v����1�U�$!##S����&�2����t:��ߏ��nx��?W���@OO233!���p��7c���x�G����/��N+E�) ͌�`1��]����0�v��{�n|���U�����|X�bŤy!���v;���cv�`0������]�v������Җ,.�c��=Uĸ{�
F��/����8��`�ʕ+�b�
�ADm^�ِef����͛��ڪvIa&�|e���`G;v�#"""" ޖ&4ݱ�Z���/C�����)��rO�a�>� >>��>�@ہc]��_�o�z�P�v����t�h���T�.5�:�Q��O�������ޯ��N��}+~?ڟ�-j��J;N�?�۸�E�,��!i�ii&ȲQ��du�]EA��۵Z-.��B��׿ƪU�Ɵ7��n:tMMMS��u:���QYY	���p;%A`��Q^^���"��擞?t�����sɒ%���p��&��F*���� "��˻h�����;w���W���klg���J�}���'(�ш����t����F�|�	c~��臡pi��=� ����N�❂�ۇ�����=�o��:��H�eTUUAQ�ڵ]]]p8Q��h�4�v;���q��A���T�NJ	�|�P��x��
%�z_3MN��ѻ�U�n~ �1� geCc2�tސ�_W'��ɵ���{u�_���~}a1B��=�<!�H>܆��v3���k;���@������Ձ���&��N�*��}>������0fp�G���/A�a-�{4F�m��4��� �N� �"";y%�T�WUU��+����i�`xxmmm�x<S��l6��p�j�ƲL���X,�X,Fww�I��|>477�����ٰZ�Ek֬�駟����_��P2�D1�q"":	�ނy_�u�e�x(�[o��/~�Qm�:���n̛7˗/W�:Z��-��͌���A��������f�Uߍټ'Ҙ�!Ⱥ��Gs���
5
���|�3 ���466"###����NF�����vc˖-p8X�d��5E�õ�H��DDDDD�F��N�2^���H�~��8e��C��R������S�20��6�K ����v���ͨð��9n7���Z�l/�F2ƪL"��T������+�����~?����v��|��lFvv6�F�Rr2�L0�L�x<���<i�������f�99900�͸��K�n�:<��#رcG��X҈"0��DD)'�����w��{��&�=z;w�L� ���V���ի�6��*$I¢E����.��(

�W��Ԅ}�%�X��\X��{;MĀ{ʈm�;
!���=ZfN���@EEQSS���:������@ ���z&�	˖-S�{rҟ)�n�AФ�?�\ADDDDDDD�J�a3�ϋڃ��&-��c��,i��Ҧ�[)�]�n7�͸��p�率cB�������=�{��d����l�G�D�3p�\�z�������s���jkk�����	I������n�	۶m�C=����8DDDɩ�k�b߾7�{'��ڵ���R���	�z�X�bEL��(b�0�xW���F���L�x�ݰ���1��x�9����(10Ř*b޹\��U�Lo��t�S\Q�r��~�z�\.������E�2�ٱZ��h4x���}���ONvә!�(I��;DY�
��������T7�Fm���u��v�5Fs�ʕѩJ�p{UUx��w�y����n7jjj���y�p��h���BII	�픒�z=


P^^��6�y����ѣ���AWW����3�<���������W����@�]��/o�Bؼy3FGGU�*z����r��j�*�ۓ�(�X�`�VkL�q��hmm��W^V|;��cA�6-7.sQbI��]jbܑY�u���1�r��O����u����vcǎ��t0����3����?���ǲe�`�Xb>更zܣB��j�w��z_3��{�ҴV��t잶ɒ�5_�ʈ�T�R��n��;���:��1�ǃ��6���z�N��^�T���PXX���ttt`hh(�y�`���CNN�V+�F#���
TWW�@mmm��'""J.��������['�a�֭X�~�:��������`ٲej�BQ���	���9� jjj�755����y1��x�5�̅��T��4�������V��^�n�ٰv�Zx�^�ر�@ .�b����z��z�۷###X�x1G�拴����"�R�#����HDDDDDDDDsE(Dk���4��ىޣ��ݦ�   s�F�S�r���J�]�Y�W\q�x��@ ���v������z����1�0H���F#���188���x<��獎����V�yyy�e%%%���;��O>�$�^o��'""J���+ž�-A�;8�PSS�L��    IDAT�ۇ��T�̌}�X�jw{IB���p8HOO�����a;<�el��-f�H5�m�q���"�wA����Q�#V���z�\��@ ;w����`�ݐ��"�2l6�k�.̟?yyyQ�'Ң�؎t�4���kt\$DDDDDDDD���H���F���������ؽxQ�`M/�N�{�D�.U��yyy��꫱hѢ�1�ۍ���I�' �$Ip:�HOO��n�D��b��b���v���}��0<<�Ӊ��h4\p�X�|9��~|��'q����(9�2�0�kw��+����HOOGNN�
�MO(���0N?�t�LlB��jjj�t�R��_������a�Ͼ��Ϻ�hBNˆ�a��"����.�/����.�rԮ�$I���Buu5$IBOOOL�#��(����hooǛo������^�fSl��I��~�S�܉������(e��C�(P��A��Y>v/H��!�y��DI ��$��_�2����p���Gcc#���&�����t���###��v���l���@nn.4�Ȼ+�A������v�KkNNn��6|��߆V��g�DDDI#s�����sa�P�7o���
UM��v#//�W�f�=8p ��K Fmmm��Ν;Q��
�=7�󝌠�![��6%�S��U5�����H�x4;��:�>F,Y��ׯ��bAOOE���D�� �͆��^lٲ�w��uG"����`���S� ��R���dL� rE%��ބ�"@�����CJ ����D;�nw:�ظq#�����?����šC�0000��,��ʐ��I�}a���p8�.�x<���E[[B�DQ���<��X�`A��&""JE�}ZGaظ���믿�@ �BU�A�eTWW#77~�cR���0>���߿?,4��ۋ�?9
�i�Em��Ц�ŵ[<%~w�
1��{�;8$b��x���X�~=�������FZZ� �z�-|����=9يSɔ<7��&Yj�7�%S���������b���"�@	}�p;ݑA��5U%�ٰ���dL��R!�^]]������ ������G���كN����BQQ�z}<�%Jj�$!77����vcU===8t���� ��q�F\z�\lBDD4C�9%�{�&<���Ӄ��~[��&��|�z�8�쳱x�b��!�tuu���=*�:t��^P(�ǟ{��ߏ�ӥћ!�3�:'%���"M���G",\��|Q��$IA�n�.�.�]]]ؽ{7�f3�|#UY�V �{�QQUU5��ɱ�_'�����d[F���.#.d�"��eF1�5�]ѬȊg��V٠v)D������DDD�dh�(FG���5 ��KZ!,�X���!�C���f �%�d��L&|�{��9��Xh���]]]�>��h4p:���Ș��4�:�����������~x�9�χ��z8dggC����/����q��w��>5�KE���,�y#Z���c����Z�X�|y��R��g>����i���l��b��5���p��Ѱ��^����]���_h3
�6%.vpO��{C�]�#��}*���~���,�[�.�����Q�"�����?�[�n����_;22q��������Fԙ�1��.���7�� ���O�xdE���Zp����W��YY?؅Ş�� ""Jx>� z��b�� ��0�� k-`��(�%{�}ɒ%������p�XP���s�p��jEyy9��Dq������
deeM�s7��}l����B�y����?ϟU""������}�#۹s'����z����p8P]]�p;��Bؿ���������9l����G�e���O����Y�l*FSc�=Eb:����Q�>W�;�Z����������xf*&��^�ł}��a�֭����5�up����=d{��EĜ6=��nѴ�CA\��;%��p{��0E�E�S�Y?؅UC�]9���hv ��Z�)�%�đ��vI�p��cÆ��8�|__߄p�dYFaa!\.����R�(����Fii)����χ��:���AQȲ�+���_�)u�$""J)� ���.�8��m۶EG����k���r�|>J<>�5553�b���&l����6�`���*qZDI�=7�sR�b�=Eģ���~sKQ���1W�c�z=V�\��+W������AR�,˰X,�����͛���:鹓�����*/%�2]��D�2�]%��)�n3r��U��h�n'""�EQ0<0��7"J,�n����]w݅K.��("���---�_��v;���`�q�N"����"77�9���ӃÇ��>^UU����-�g�DDD	K2�Q����1���Bؼy3���c2w ���V�X�e˖�dJ���hll������طo_��~x���Q}U�+��6c 0�L���T!�b��0�D�����t��]+�$I+P]]I���ӣvI��DQ��nG{{;�lقÇ�����6&h$H6g<JL�l�6����2
 �sk��}�S"�n#(
.r�3�Ns��DDD����Q����ԑ����+W���Fq�n�CCC8t�Ф��Z-���1o�<HR�g��� �Á���I;�{�^���x�g
������o�_|��x"""��!w>J��S�&��@ ���:����:g__���q��gC��F�ڔ��92�l����޽{ò��@ �}�y���9 F�{Ɗ�`����h2�M&���iH0E�z��M�\��~"A�d��_��===3��(�A@ZZ�e��޽{�&}�����!�^R��Y
!���"t�%jWAD	�!w��NnÐ;�u�E��(�}�r�x~���h�K�p�(����Kq�u��`0@Q������~�?�|A�t:Q^^�٬B�D4Z�EEE��χF�<OQ��n<������(���Kp뭷&��Q<��G�e��x�����W_�t��L����b���sυ�n?��Q�9t�FFF&=�w�ްsB�{���ChL���Dt�¸�I���"HrL����2���!j׊���r�_�������t�G�xIKKC �?��|��G?tk3�PY�����f�]F��J ʉ�LDsC�4M'�>�!w��n'""�.I�"�73�HzH��lD(��(�����d�[�Vlذ^x!A���(><i�I�����28�Nvy&J���']�"�{�9|�� �ŋ�{�AEEE<�$""JH�����uWG<��z��K/���wV��z��X�f���O�LJq�`���G0;�(
8�����c|�YtW^��4eN�͘A�N43�K�BDI��k�r#f����d��%~.+,,ĺu�PXX���ްm?���j�b`` b��=O��R�>��<�w��	Q6�򁗈�C�4��$�>�!w�kn'""�>I�A�3@`I+��^���h����l�B47$k����w�}7�,Y�Xg�ÇO����p���t��LD�dYFqq1���#.N�$	;w��s�=�`0�Á_��8���U����(�|��}�_#�x<x饗&]@I ����g?�YTUUqa)E�����Ç'������������P����x�8N2� �3�>/%>�[��X����Y�9��̀�$I��bԏ���,�[�,������'� ,ǐ���0�4@P��h`t-� �oID4��\0�p���i�`����(6z:a��  ��A�T���NE����?�|�q�p:�Phnn���F�e�\.���B��5Q����Q�(�����#�<���Ȳ����
W_}5$��g���&#h$��ǳ��_����(^y�tuuMy���~�\.TWW�`0D�TJq���hmm�i������D���{��z�y�.�F��Q�y)90��Bb����ޑ����r'b���l6TWWc����x<�!��H�- �!o~�+I-��	]f��e�2}v$�C�2�(�0�Nj:�p���Im��Fo% ��(J0�s�.��NA2��eY��W_����
�,������aҰ��jEYY�Vk�+%�X�j�(..��bA0;.�y��ݻ �~�z���H��>""�X��]��0-�x����W^A[[[��0�LX�v-�Ng,K���� �ۍ�������;w��-����
�ڌY��)�1��Bb�� �G��<E���p���r�J�\��`p��1Q,L��]�ˀ{�r�C2��.c�$���r�� �$Ő;�!��1��Zn'""�����=�Y �d-�(�Q�J�p{ZZ~��_b��� �=������\IE�����r�s3Q� �w��z{{Î˲���{/��2 ���w�y'\.W�+%""J��׽Cނ���~?^{�������~��V�Beee�J��������;�k�.�e� 2νZ�� ɜ��)R�)D�c����`�V*��D����b�ڵ��F���*TWWC�$����]���*�����j��*h��^�1X`*^�XKD�Đ;�S4��cr�xc����(6������ �� A���f��"�YJ�p{nn.6mڄ��cIz{{Q[[�?|�e�ш��28ܙ�(ٵ��ᡇ��~<A��ֆ'�x���p:��կ~�3�8C�J����dq���נuF<��믣�����X�d	V�XQd,�bott>� �}�]<��C��v�څ�?�A���R�(��(PenJ|'M!b:����+nFF"�v��d�2Q,Y��ׯ��lFwwwT;�/R�]�Q Qχt� H2L%�Q_4W�:#̥+�m�C����aȝ��v""��pw���i6=`�@�OW�,"��d�/^�w�urss
���҂#G�D|��������t�o�EDs���(��y�����|�?������`�O�S\t�E*TJDD���0����s�F<����6�&�)��Q��}�݇}�� �����/ ��݋�w�#�_~5�X
� ]V1Q��)�0��J1��D�� ����Hc�%�2��	��FEE�?�|8�N��� �]%�����7���U�&u�Z=,gAc����E��3!H| BD�Ð;�R,��cr�Xc����(6�v7����E��a���3d�]�R2�۫��q�-��l6������}}}a�i4�\.dggCගD)i���x��#� �(
�y�8p �(���&~��@�$*%""���������.�x<��G��o���(�����;�D]]݄�͛7��ß�� ��:�`m�<�Z�*sSra�=ň��õ�����Fu�����U��������r����1�L4S�nt��hY�+!A��\z&$S��/��‥�,��^�R�(����^�K�$�p���)Vn'""�>EQ��Z�Q���V��bh�s���\���A��_�k���$������Oxs �N���Ҥ����������o�;{O�elݺu<�w��⦛n���0Q$��|T��6�N�x|lٳ�>qw%�hhmmŦM������=J�nP-�.�쐬���Mɇ��;D:�»�Eu�T�!����u��a����ː�ޤ����\	� �0����|�P�e�\�O4��AD�ч�����!w��x���0�N��p;Q�~�4�,] �(��VY�Z����I���%I�5�\�K.�� `hhuuu���a�Z�V���B�㎜Dt������?�7�xc�}q�F���Ç��?���`�ҥشi22��Q$�͉ʟm��`ɤ�lٲ=�FGG�X��O>��6mBooo��9���=�����su�(�u�}^J^������{�~�?��h���G�Z��f�a���X�l<O�;�Sj���8΀�zA�>�����@�tQ6�T�O0�-<֮��He�S4�n3r_ʐ;�"�ۉ�����Bs�n�MZh�h$,�rH2;�%�d���f�r�-���p��MCC����A@vv6\.4���hnS۶m�O<��Y=zO<��~?\.6mڄ��|��%""��$k&*��
��Փ����cӦM���_a���|�M<����3���y�܉����:AsA��*V%XOɋ���{7"��f[�e���]/���z�\�g�}6�� ����.�H���6cd{�
���d��k�usWc� A�.����![�]�-�өP3�>FP�C�t
n'""����^�9�4����6X��5Z�K#�YJ�p{ZZ6n܈ŋ :;;���EQ&�'I\.����(��HSS~�a������|x��G188�Ӊ;����*TIDD4�i�i���5��q�紶�b�ƍ8x�`+�d�����O�g�	ۍ ���+C����q�d�lsƫLh�qɦRja�=ň�B���������6�vG7�a�ۣz�D��hPUU���j��z�iJ>�/�Ϣ��J�j(A�@�Sk�*h��ŧ�� B�(�u��B`w"��r�٘��1��l1�NDD}C�G��Y�4�P����`�AP�� EE����v;n��6AQ477���3�<�ш��2X,�$�D400�G}�w�;&�z�)ttt�l6cÆX�t�
U�}��C���F�n�����a�w�}x����M���w�y'�{ｈ�%s:��g3�q�=C�W��s!��c>�ީM5� A��t
mF7���Du�?%.\��k�"--n���(���������U��NFԛ`,\�5�9K!j���-j��g�����y�!j��6�}��L̥p���i�n'""����~t�F�M  ������0D;���.�+a��YYYشi
����ɑ�fCqq1dYV�J"Jd�@ ��_��o�=;�h4x�P__���o�g�y�J��q���/݌�K����`(�K/��x CCCq.�՞={p�m����1�q}N�߼�Փ_D��,�����9-'fק�ƀ{
��V��##R�����@Ԧ�Z��aAII	���������?sJ|ǭVǷ�6Qk�!�օka.]]V4+��<p m�g��Rv��@�S1������!w���nÐ;M��DDD'�fg�EQ�v� �l@	B��0Zn'J`������{\^^~��_!''�@ uuuC0����E>�%��Qo��6���?bttt�1I���k�a�޽�e�]w֬Y�R�DDDs_ֹ�C�϶@�fMz�޽{q�m����6��Q�	x�g���bx8�sNs�J̿�]�˦�����w���ޗ�3B���u�Ƅ��)�:0��9��#���@�n(
� �Á����\/���� ''���صk�f3�Z��e��"��h�i0-W������  (?������"��� ��{�+�@#A�t��Mufh�VQr�?�^�#\�C'����1c!w �e��\�E�Mm@p`����hx���F �`΃ 0J���-�^PP�[o�������hhh��;q�� ���EFF�JUQ�9t��q\r�%�X,��$��߆���駟����0�Lx��U����h��_���lG�_�HӮ�������;�Duu5���/A�ߤOutt��GAKKˤ�d��
_�gF]�E�	rz>|G'��L��zg)��jC|�LA�9�s�K00���:a���?�7333p�Bff&֭[����ܹ `0ĸ�?�I�P���a����'�&��.A�!�3 3bQ�bȝ"I�p���i2�M_���ٚ�}���m��d�F������r"��d����bÆ�X,���������p�(�((({�FDt��������K.Avv���$I�裏��xp�9���+���(x�WT����h��ea����G�ۏG<GQlٲ���_�����Is��(��?��^x!lg�1��׷~�����?    IDAT3.���5��a��Y5�9Kg�'�.�HA�l�y�U�]�}��a㽽��o��ؕ|��F#V�\���*�A�]�Yww7�@ظ��u*TCDDc!�|�w�)�%R�}�X�}�ǭv)4G0�NDD4} ���V�Д�BA�@�=�%����i}D;�z�T������o��b���(jkk���,�����v"����<���hll�0.�"8�͛7C|�;��\�N�DDD	@��(��1|�^�乶��lܸ������6�zzzzp��w����vC�",�����ct�B�:�)]CD蝥�l�K�ǀ{*�S~������a�����r8�b&�Z-���p�9�@��```@�(N���"�[��J�����!w3�>�!w�p;��x�~���\x�Aw7�ZD�X�.-֥Q<�=ҝ4����J�t�M0��z�������p�^�Gii)w�%���z�����={�Luuux�W ���
|�_P�J""���\�̿i��哞�����/���o[dF�MQ���;ذa:4�yg}n�}n�O*��gϺ9� �eC�sGD��S�F�7�vMn��e}}}Q���-�h�DQ�ҥK�f���f����]�Xsssؘ6������C�-���cr'�ۉ��NM��(�~�I���d H�����%�d������o��`����������%%%�en�ND���/b۶m�A��#G���/C|�[���?�y��$""J��eXx�Nd���I�;r�6mڄ�{n�.ޔ<ZZZ�_�
O=�Ԥ��E�}���{�:S��dt�E�z��Q���Z��{���*a�g���6~�ht؛L&X,��^3�TTT`�ڵ�X,����7Ihtt]]]a��e�@DDɃ!�Ԕ��1��.�ۉ��fK�_��j�2�
�������?Ig�uqDe�%Y������rL&�����Ѐ`08��Պ��Bh4��GD4[����7���͛'�����6��o� �������V�J""�� �Lp}����ϐ̓��
��y�f�x�ؾ};e���<�}�Ylܸ�����g]t.��8V~#&uh�6h�rf�m�<H挘�C4�S��3A��O<��������:��GGyy9֯_���|����=�zZZZ"~�M[��T����(vrO-�nÐ{�a����(:(p�=h��F<��CQBЈ��y�2��%��<��(ܞ���6�b�`dd$b��f������ǹD��w�}/��r�sƖ�������w�f��*$""J�ӿ��w#�3�z�������c��;�@sss���XR��>n��Flٲe�波ֈ�o>����mƼ��$�s!M��֞ٚ�z�"��%���n]1�fؘ�(����a�233ٽ"�rrrP]]���2���]��Hx%s,�PQl1��1�>�!���p;Q��D ��`��c�X�l�qD4+�nw8���[����ǃ����pCZZ


bެ��h:v�؁?��������.���KE�\s�>�l�$""J��|���K(��S����q�F<���8z��Ձp�������@x��1��p�.d��
�����"�����iِg��(ZpOaC�`ͫ������<�N�3��$ ==�V�%K��x��x�.�f!F�9L[�I�����b�!�����1�'?�ۉ��b�
���`e�;Y� �FA���D�l����tlܸN�^�7b�����ۉh�ٻw/���?M�\�����W_�(����k�|�r�$""J�g|��8���+Oz�񝿟}�YƩB:U---���p�����e��$�_��ox��8Vx�I�.�d��drZ6�����Dt<��Ma�in1q*$����&����ݰ;Uyyy��#F�+W��駟���K	�ȑ#��ۗQ�j����g,�ǐ{RI�p��ܓ��DDD��0ҍ�B(�C00�``^� �6Ey|<��(�LD%[��j���[oENN|>&E ++yy��t��a<��Sa������o@�$��g?ÂT����(�H&;\�?���^�>���lٲ�_=��׿bhh(NU�L9r���op��c�����(p�sN���� �ԌA��u��k����pOa��A#�|��@�v*�P(�]��z=222�zM�H��ᬳ�ªU� I�nmA}}}ؘ�`�uѹ*TCDD_�P�b�=i�R�}C�ɇ�v""�h:.�~\H�
����Pzk0�[%�F� ����������.����l�v���[o����������pNVV���U���hz���OO�����lݺZ�7�p

�CRDDD�m�z,���.����7�׋���o����g�}���q�����ֆ�{��v>���6T��T��Gѕ�B�8�Xed�9�quh��!��X�1��8���9g���)l���3�s���G��N,Y����0����a�`0��_���@��*TDDD�'�T��a�=y0�NDD?-�>�B���ifH�&�ǟGD�K�p�(��я~����I��999�Q�hjj��������������l6cÆ���T�J""��"hddV_�ݼ�A�|c����xG���z
���q����(
8�����Ɔ�}����%k&
�~/�r/��Ʊҩi3
�љ�͘��T�" ���x�%�5�����nx��Y,�l��^�N�����հ�������LsCccc�6� �8��*TCDD���[*���0��n'""�������+�@,J"�YH�p; \y啨��B @}}}�=���l�@�(�466⩧����;ሢ�={�`Ϟ=�����7��٬b�DDD�G2�����a��;���sS������;���[n�}�݇�{��4`M��m�6�z뭸��{�o߾���kV�]t+��� ��@�Hq�v���r��,�+!7R(�4+A��?l���@ �4�[���+�ۓ�\.�޽;�פ����---8p� l6[��7�_MMMؘ>��3U����H]c!�ߥ��;�$��?5r�].�M$�Ŋp�#�����'��J�p��^��}�s�hhh� �Ӊ�,��(1577�駟�׾�5h�Z �޻�m������2�p������v� ""��3.Eُ^���mh}����+�����c�������ʕ+q�g�j�}��T��ىw�}��>�<_���Z�]�~�zH�X�,�_6�-��Lq�F����|��l�ܳ/l���#��z�Պ����^��o޼y8��P^^�������)>������6�8�R@���Q2c'���p{8vrO<��C�`z��C!��Ԗ����+W���EAss3<τ��N'�}'����܌g�y���EQ����w���a�����k!��$Ѭ���D�Ϸ���[`.;cZ�����/��������o~�={� Ƹ�������஻��M7݄7�xc�p��5�y�`�]�Q���#�N4��2A2���tA�aw�U'�������Q���ra׮]Q�&͌�n��ի122��?� �׳Sj<��Ԅ/ Dd��uu
"""�#��=10�>9vrO��ω��t3xm(Ȁ;���1�^^^�k���(���5,�`�ۑ���RuDD�UWW����o��F �$	/����կb�ʕhii����+%""J\�հ޴C5���M���J�͐�A|������a4�x�b,[��-�(�/�ɄB!444����Ǉ~�wz��D���.Gο������*�	����wR?Q_f:;kúQ���G=�n�X������ި^�f�h4⬳΂��î]���x`6��.+�B!<x0l�v�y�f�S�"""���!������1�>�1�NDD�.����kJEQ��W"�%c�=;;7�pt:���p����l6���U���(6<����/���8��ӟp饗�_�*�����[o�\)Qb3W�DY�Jx��E�+w�����������oߎ�۷#--K�.�ҥKQVVIb� �~?8�ݻwc׮]��ke�Yk�Y��$s��>K4��݉ ��zK̻��r���'[��N��������`0Du���b����<�Oӣ�jQUU�P(��>�HKKS�������s��U����hn҇����O��G�IG�%1��P�c�}*����v( �-j�C�Y3؍��\pMDDo��@ �ӿ/�������(��.�hJ�n�X,��[����ۍ���	ǭV+


�߫����'�|Y�q����	����~�]v������ѣسg�ʕ%>C�"}�q�}�vt��A���Q��S�@?�n݊�[��`0`�8��PYY�rY���>�߿{��������ͬ	���Ld��
�UA�f�n����w H�����V.���(t�����6���Du.�����\���F��tjDQ�駟 �����#GR��Q<|��'ac��r��W�""���
�ߏ6�]Ѭ�P��6�� """�sf��= E	A�=7Q�$c�]�$���rss1<<����	�-
n'���s�N�L&�]�v|,���3.��"��'?���^���N�$""JZ{�|;�.ڀ��o���ߢ������z�����;�c� @NN***PYY���X��X�w���8|�0<����3� �`_�y8��!�egĠJ"À; 4�4��n�r�j����=��	�(((�,�Q���� ]]]����O����@EEPWW��6�e�^ww7����Ɲ�_�!%+Ef�� �P ������!�� p��c�ESS��� F���v"J��L&V�X1>��ۋ7�|��ո������^�W�*����� j`]t.����hW=���G�=_Oӌ���ގ��vlݺ �p8PRR���"�\.���5����~?�����Ѐ��z444D�SM� �Ry62��:ҫ.��h�n�D���?r�����N$J�3���PhB�9
���Q�N�$���6�ץ�***BQQ���q������;����������t���d[޶<�;lf�(�0�$�R2Ҵ��+m�6���&m�jCCf c��^x˶��W�����@H�e[�I~==����{�o��:�s>_�Ov;_��������ټAe��˂4      @r|�L4�xo�l_j���2)p�n���\�R�]w��Ѩ����F{��&N�H� �_|Q�@@�f��;x���ӵp�B}�s��7��7� �B�ʝ�q�|]�n��B{��������i�>�s544���A�6m�t�w����7NEEE���Snn�rrr��z��]�P(�����׫��Z������T]]]��υ�p�2�ܢ��wɕ7y�**H���J~�����+���_iтy}�+++UTT$��6�����Nmmm�z^������Y;w����ɋJg���IǏ���2�O�t�-H      ���vp��"��n0
��jq{qq���~%	?~\===�s6�M�&M��`�K$zꩧ��zURR"I2MS�7oV^^��-[�o�QO>���I �<�fiܭ�P�G�����W��_�eǳ
7�<��%	��թ��N۶m�3������tedd(--M�`P^�W�G^�W^�Wn���>��E�PH�DB�XL===���Tww������ޮ����?[[[U__����s���0�+^����\p��ʆ�� ���e�˰9��E��N���ٵ���hT555***�5�N��m۶��]YH���]z������a���X�jtغuk�N�ݩ�+?kQ"       5�+j?�R�x<���S!�H�#�X-n��|��W�"�ۭ��*uvv�����'��:�=% `l�F���/��k�*77Wҩ~��������w߭�Ǐk�֭' `�3L��f�Vڬ՚(���N��xN-���#�����{���v�����3�f\���7(}��rf�"�s�^xx�a��N�R�%Wh����+**�R���x4~��a?/����jŊZ�h�b����q7577�����x�%k����?      ���?�ϸ]	��>��XxX2Y)�S��i��������*((PKK��̏7N~?;���uww���E��yM��/~���/~���   u��Tp�_i���м��j�_<����B���2̳��2���3.U�M�����YS��9�����Cw�a�g)�R��u�z��͚�w<���J�ƍ�5Ǐ����>�30:8�N-Z�H�DB�v�Rcc���ӭ�5�lڴ��v�C��>hQ"       �L�M2�2�X��<�s$�@�X�����m��Kҭ�ުE����[}���򔑑aQ2 YZZZ�_�B�g&���>;�XL�<�n��=���z���F-N
 �����R��7)��$I��V�ܨ��o��|��ʷ+�Vgq�s��)��d�|%埲T�)�e:�V�0����͓�X�-�k�J�h��4wά>�*((��6�w����ӧk���I���3Ceee�����B�`��T#CUU�N�8�o<�ҏ˕S��@      @�������'�K�{|�#�;����%%%c��{޼y�����T^^��u�`0���<���SUU���zJ��Gzwߩ��ѦM��x�b�s�=����/�S  I�y���F�ykz��͕�*߮���:�[�5��]{X��Ӝ)���L���]0M���,��d����;(p������))p���뵃͝�w<����R&L�5�^�JJJt�ȑa?7Rkڴi�6m�>��G�*##C�iZ��DBo��V�q��     `,��r�6��};�;��������5�կs�X(n���у>(�4U^^�p���~�_�Ǐ�0 �\�������j�*I��7lݺU�Ǐ���_�}����7ߴ8%  �3�HΌ"�_�g<�R}�ؽ��M'i�>��Z�Hs�"muJD����awɑ�'gf�iyrd��#=Wά	r�ʝ?U�@�y�`d���ؽA�m%b��X�v��m_�������P~~���s�sz���jnnVSSӰ��7e�M�2E555ڷo�|>����KۡC�����o<���to     ��5��I��3������QG�G�P���ˈG�4�v�А�Ln�q{3e�����z��=33��(��4M=��������U[�{��&L��ۙ �߆����ٳgK��v�֭[��k������UY96~& �B��,P`��A��u�+�ӥxO�b]��GB��tz����t�esd�es�d8\Ɉ`����@14�!Gz��M���ў����+�����t��q���&eݩS�j۶m}�j`t���W~~�����s�N�\��� 1҄�amٲ�߸���覯Y�      H�D���]�i*`���%���Ӥ�p�$)z���9�����c��(F��T�.I7�|��Ν���v������������ ����~Z���*,,�t�{ů�k�~������/}�K�F��8  0������c ��3��=�#ô�d���?Ն77����UgggR�t8�9sf��z����KUVV�P(�������l�2��I���,�       `���#j����1 H2e���d��O�2E��G�Dt��	%�޹��"y<����D����y����M7nTii����   )��ŀ�&{ ;%k�<iz���_�n"�Б#G��n PIII��ky�^�X�B�/V,S{{�Ց�]CC�����oܙQ��k>gA"       u.��ݍ
w7���\5�/���>E� ���)##�����v�_���v�N�<�X,�;���5f�O H���=�����Nuq߽{��?��n�Ieee'   `5
�1(GZ��H�Z������o�ommU}}}��-,,T^^^���9�N-Z�H�\r�l6�Z[��6ÉDB6l�7�    IDAT�źq���L�ςT      @���Ty�iU~Zu'_U����H ƨ{�WEEE���UGGG���Uaa��� `�:z��^~����6�M/���b��>������[�   ��(pǠ�S6_�:N�6N[����~SG�U4M��S�LQ H��12��y��iժU���jii�:�yٹs���{��+k9��       0�,Y�+��R�PHuuu���C'NLY�( ��|��>;V����zJYYY����-L   �j����nL��|��x8���Ǔ��i��5k��nw����2m�4�^�Z�`P����[ߍ---ںuk�	��Ļ�+|i       �|eff곟����N�8ѻ��a?~���	`�{���4�jnnֶm۴l�2�Z���d    �D$N�tze���l��Y�덷�����Rkkk��u8�3g"/0�'O֕W^���ǫ��5�;�x<����+����]�i�K�Y�
       ���0}��W PUU�zzzz�


���-L cGOO�~��_)�H:��wӦMjiiѽ�ޫ��L�   ��8#GFQ�ֲ�zS������:t(����n�f̘!����B����U�Vi�ԩjooW8�:Ҡv�ء���~�`����u       0�\u�U*++S[[����z���Ҕ��ma2 {jkk��K/�>��lz�'������|��d    �B%/��tzd�e�l=ς?Փ���o<
����I];==]3gΤ������K/�Teee
�B���:R555ڶmۀs���l�`�       0�dff���V$QEEE��nWQQ�C��d˖-ڳgO��X,�W^yE_|�V�^ma2    V��C��(L�b�M5��k��]��*++��֖��3224}�t���u0ry�^�X�B�/VOOπ;
�ZOO�^}��w1H��ae\|��        {>��O������B�h�w|���r8&���g��kơC�TSS�{ｗ�3   ����ݟ���܅3��x�ډDBP,K��YYY*--M���N��-[��+W�n����ղ,����:::��ۼA����        {�-[��K�����O���l�����������i�Z�n��^�������t    R�w�3X�Ү�Ew��^�7��ݭ�&}���<:�Cҩ'eeeZ�j��~�ZZZR���]�T^^>���?�����R�       �����铟��"�����{��n����-L �'N���߫H$z�W�h�"�X���d    R�w��p�H�_v��ݦ�x��TCC����!''G3f̐i�S�M��իW+++K��ͽ�����J�7op.k��Zz{R�       �B�v�Zeee����w7a�04a�^+�z��t����ǇVMM�>��O���Y�   @�p%g�,�a��l=W�$�ޔ3`1��Ç
���!++K3g���%�(..��_���"555)��]]]z��W,�wf�ӄ�=<�k       p!�={����
�������w���@n���d p���z��'���#�Ԏ��>��222���}��t    R��]��f�#X��5�}D��~g�"�X,��{��v�H���͞=[v{��1:�+�дi�����{��|E�Q���K����?i�*���d�e�Z        \����>��qUUU��eg�pwc @���f��⋽�c��6lؠ���Z3f̰0   �T��g�ȑ�Ha�
�P䢏���_�7
�t�����HOOWYY]:0�`0�K.�D���S(�0�,lذa��$��/+m�e�u~        p�m�ݦq�Ʃ��Z�HD�d��5n�8����m۶m:t�P��{����C��w��   �1�w�=Ð3k|J��rt �Jmݶ��\cc�***R����j���JKKK�z}�^�V�X�%K�(������ϱi�&>|x�����T���1       ����|�x����PSSS�xAA����  ��n�:�B!I��fӺu�4q�D�Y���d    ��w��'MvozJ��/ԋ������+//WcccJr��v͙3G999)Y����ТE��r�J��v����y��v��9��3k�&�e���
       �k�ڵ����������Ȱ0 �]mmm���~�����S{���wܡ��L�   H&
�qΜ��e��/��V��ս����3�H$t��uvv�$�i��>}�JKKeFJ���d����ʴz�j�����WTTh�ƍ�v������qc       I�'�N `��;w��.]�����מL�Ըq�,N x��۷��{�ƍ���뮻,L    ��V��e8\rd(�Ty惇mQC�ݧ�?�-}���L�b1�ٳG��͓��JI���|y<���;
��)Y�״i�4m�4�������JOO�i��I���Y/�������ϝx���M�8�q     ����#3-��#N�4mm�:0♦�O|�
��jhh���˓��0 ����֭[���ON�S�i�^К5k��/���VG   0�(p�yq��)�٬xOW��4]>5�}\O?�?�a͕}�����ۧ�s��f��$Ozz��ϟ���;7���b���Z{���n���??�M����\vo�S      #[<ԭx��� F�+��R%%%*//�m>��x���mq2 �@Z[[�~�z]u�U�N���بO�����0h#1    ��iu �r�!Wv��H�ά	ڟw�^۰��\GG���ۧD"u��:�N͙3G�'O����IAA��.]�6���c�c�ˮф����d        �]>�Ow�q�:::���&I2C�ƍK�k^ ��۴i����$I6�M�?���L��K.���d    ���8o��#{Zn���L��7b��g��~s---ڿJ��%���P��͓��M��zzz���}O����{��k���˰��        ���nS0Tuuu�XNN�<���  g����3��vk���־}�t��w��rY�   �p���Q(ӑ�_}�.�Sb:q�D����F>|8��|>-X�@%%%tsǠ��~��A��:2
U���e��)N       ��UPP�5k֨��Q�PHҩ�zssS��	 p�jjj�y����6lPFF����ZS   nT�bx�\�Ŗlۘ�����cjhh�7WSS�#G��<ӻ�XΛ7O�@ ��cd�D"�����C�8o�k�_>/g��'       `l[�v�L�Tmmm�XQQM� `y��W���&I2MS�ׯ�G>�^�   ���`ؘn����_�0�[�����jnn�7]UU5h!q��|>���i��ɲ��d@_�i*==ݲ���y��۷o�y��U�矑w��'       `l�2e�/^���:E�QIRZZ� 0ʄ�a��w��}|��A�l6�z��   0�(pǰrds�R��aʻ���?�ީ�~555������B]|��***���=N����E]�9s�XR���ӣ�~��ڿ���ݩ)<����)N       ��w�w*���
l�


,N 8�w�Vyy�$�f���_Ԛ5k��oAS>    Îw/Ð+�D�iK�ڦ]��_��Z����~���'��g�d��5i�$͟?_�`В�`0�hƌr�\2C3f̐��LY���.=��C:p����͡)�����^��L        \(�O������������l�\.�� ��s�=�x<.����mmm���,N   `8P��ag8\rf��lm��/���8h�����{ɵ���Ӝ9s4g����Y��B���5{�l͙3G>_ߝ�f̘����---������G�8o�6M�?����뒞       �ѝwީP(Ի��nWnn�ũ  磮�N[�n��^��.�L�ƍ�8   ��E�;���ϒݗa�ڦ�+㊿����:::��766jϞ=��b�{O0TYY�fϞ-��oi��&--M�f�����1��ô�4M�4)�Y�����o~S�6�J>�ce.�HRs        p��5k����TSS�;���/�͂� �j���vxokkSee�n��V�S   8_�#i\9�2nK�6�VY?������ͷ��j׮]
����+##C���WYY�233��3��[�~6���B���%%ϡC���o}k����d�]���_)k�]IY        �����٩��vI���>m� ����ե6H������r�J[   �y���c�r�M�aZ���p���o�g������|GG��o�>`�w+�[��`�����4��
�4����y���M�'O����\�7o�w���nd�|���u�X�'ú.        xς4{�l������0S �Ӗ-[z���B!�8qB��r�ũ    �*h�T��-g�D���^�~��UVV����ڵk�-70�ϧ�S�jѢE�4i��^�ՑF$�׫I�&i��Ś6m���9��f�iƌ����+���'�ԏ~�#E"����5��/)m��        �wܡ���ކG������ `��bz��W%�����k�i���8��Z    �w$�ݗ!Gz�uL�|W~I��Y�}������bڿ�***,78�á��"-\�Peee�������4M���h�ܹZ�p������c��x4u���:G(�#�<�_|q�c�Y�5�o^��t�y�        NoѢE�:ujo�v�0���oq* @2�ݻW'O��$uww��ѣ���-N   �\Q���pf��I�.�a(�O�Ɋ��qc��D"�cǎi�޽�F�<���4M�:UK�,ѬY����+��fu��0MS����6m��,Y��ӧ+===)keeei�����ܓ'O��韴gϞA��N(ӌ��!�        ��7߬�������`P.���T �dH$z��%���i�ƍ��KTPP`q2    �w��aȕS"�a�E���k�ѾDO?��MMMڱc����R�lh��S�=k�,��v[mX��v���h�̙Z�tiJ��'N��`0xV�y뭷��o}Kuuu��^v���u9�έ�        ]ii�fΜ٧{{^��; �����:x�$���Gǎ�7�`q*    ��nu \8�]��)�zG�x̲�I���7S��������t:�̇B!�رC�'O�:��l����ɓ'+
���Y���jkkS8�:��l6���+*���Y��0M�>]۷oWOO�i�����c�=���z���]�9M��J�       �
7�t����z�eff�{M 0��_�^���2Co��n��v=���jjj�:   ��@�;R�t��Λ�J$��p痪5�Kz豇t�Ջ���b1<xPMMM*--��>�?U<�<�
%�*�oooW[[�:;;��٩X̺�e���^�|>�|>�������e���z9͘1C�v�R<���r��G?:m�v��ք�VΥ�HVT        �yyyZ�t����%�jn���km( @JTWW�w�ь3
�T[[�믿^?��O��   �,���]�9��/gv�z�Y����v�W��o�LkJ�5޼~�444���]ӦMSzz�)�ݻ��`��ݭ��N�B!uww�����Z�}.Ð�����}{�������b��M�4I��3�������;��̙5AS����M�8�Q       ��\��
�����$eee��pX�
 �*�ׯ����e�6lؠn�A���/
���   `�(p�%��L%�=
7WY�0X~��?�N<��������{zz�k�.���X�iZ����n����"���Ѩ"�H��c�Xow4��o��eF�6��OQ�X�Ⳡ�@�����$UVV�g?�YoǗ��Qɟ�\v_F
R       �w��~]q��;�������S R���N���ӬY���֦��.]~��Z�n���    #X�D4�H{��Q��!l��������U����wLee�UZZ�`0hA��r8r8�x<VGQ�L����v=��Sz�g�F=ְ�Ux�ߪ���H��K=        c�5�\#�ݮ��6Ito����{͜9S�ij�����������    �g���Ƙ�̚ �?���$g�D�G���Uڼyˀ�twwk���:|��i�1vttt���Y/���i��]9%����*��)n       �v�]k֬Q}}�����V__�}��I�������t�EY�
   �PQ�k�\�Ų{ӭNr�i��=zնL���o���=�a���ڲe����R��Fu��Q�ܹS.�K���'d���Zq�f��.���HqJ        �K/�T�`P��͒Nuo���� .T���z�O6l���_ou$    CD�;�gr�N���:I/���j_����[�wuP4Ց#G�s�Nutt�8!�%�H���R[�lQeee���3���ϱ���~�7����t�S        �Ϛ5k��بX,&�0���mu$ ��jjjt��I҉'4{�l[
   ��P����0�Λ"�*6�~yV}AO5N��ϯ���>�qmmmھ}����?h�w�---ھ}��=�h4�o��k���ٳ%I��?���أ��R        |@II�&O����FIR0���8 �j7n�$���͛7�kj   `d��#�aʕ7E��ku�>��V��ү�/і-oz\CC��nݪC�)��0!�W{{�v�ڥݻw���s��N�<�{@�_X���?.GZn
S       ��\s�5jii�}����  I*//׉'$I{��ե�^*��cq*    gB�;Fôɝ?U6���(}���?�W��臿|N�����USS���~['O�T,KqR����v�ݻW;v�Pkk��uvv�g?�o�`�Qٯ��\���D<�I       �`�N�V�\���IR �x ���.�XL���Z�r�ŉ    �	�q�&w�T�<iVG��]0]�K�J��I��������h4���rmڴIǎS4MqR���ۛ��=.�HhÆ��G�Vuٟ+��/�pz���p<��       �`V�\)�ͦP($��� ��:���z��͛7k͚5VG   p�cd2L����Z��?Ӯ��U�E_�w^<�W֯W"���X,���
mٲEǏ���hnn��ݻ�X�.������X�E�(��o˝?��|��IѶ�;�       �Թꪫ���(Ir��
' �$�DB�7o�$���)''GS�L�8   �ӡ�#�aȕ;Iv_��Id�ɻ��ږ����׵gϞA��F�:q�6oެ����3�I/l�x\555ںu���٣����_QQ��������o�J�}��ǆ�N*�ÿ%        V�8q��N��{�?''��D ��hǎ���i�z��7u�5�X	   �iP����0��)�ݟeu�A9�&H+?�g:f��~��ݻw�c��jkk�m�6�޽[����v��	�B:v�6mڤC����������џ��~��Z���QY+����>'�H�����pF        Ct�UW���U�XL�C��� `�H$��۷K��=�+V��rY�
   �`�V ��0��)�iw*�Rmu�A�&-�&-Һ�;����U'���t��[ZZ���"�á��<�������0������ب���3vjWmm��{�w:������(˟yvkF��?*w^�d�        ��á�.�L�������,\� bӦMZ�d�l6�N�8�%K���^�:   �P��QÑQ(��R�����z�8O����룛�����Ь"͝;w��#��***TQQ���4���(''G�#��G�D"���V��թ��A�XlHϫ��Һ~���Re���r}�!jW��JΌ�s>        8;˖-���Pgg��Pf��5� \X���t��͜9S[�nժU�(p   F(
�1���Y2�N��Q">�Bf�x'-Rt�"=[�M/=���si��%����kkkS[[��=���t���*33�b�x�����Q
��C~��ݻ���{T��@���r��a�i������֧        ��e�]���FIRZZ�i_� @��~�m͜9S��횵�#    IDAT:u����z��    9�ʃQ���]8]=5�����J��R�mn�כ/����*�X|����}N"�PKK�ZZZd���233���%�כ��#G4UKK������بh4:��vuu��^ӖõJL�Z�S����/��p�L�{��        ����5w�\:tH��� �cǎ���QYYYںu�.��=��V�   ��cT2�SE�uG��:ΐ�9�/�S��]�����l|E�h���2Ms��%�������r��
�JOOW0���L�{�:�x\���jiiQss�:::�H$�����?�@((����pN�Ҟ����SwT���1��) ��=#S���rd��0mI]���;j߾%�k$�3'O��e2].������ijPw�E��#Ir��7c���:��V����H��'N�gr��:vmS����H��i�=�X��I2N�:����DB�*���|g`O�7k�Y?�c�v�:ړ����œ���S��N���-���9G�����9��R��N=UR<>���"��9�3���+�Ѯ�w�*>ĝΆ��t�7g���
WW�c���5��x��P6�_�Ǐ���;VG  �i�ҥ���T4���P �: `H$ڶm����
>|X�W���   �(pǨe�r�OU��B��:�����*���z��6�v��:k�tA�rss�����n��Ԩ��F���x���.�߯��4y�^���wc؅�autt���Ummm���P�^����[o������[��_U�3u]���z�˕S��5�N�ͮ	_�k��	vGJ֬����w��V���g��x�t��,��c����O��̯���R����I�/ʺ�:�ݟ�q�?�+���R<ԕ�L�*�����җ��KD"���t����6���(�֏)s�UI)�>�#_�K�o�4��~?��9����g��}C���P.}�J�|��2�w,t䐎��Զ�)��*(R�~O�����N��Y���P�S��e�+|~�����Vp��V��#�ަ��?��_:���E΍���K_�=㽎���Gt��?���!Cb*��~���dz޻>бk��~�nT  �o�ʕjii�D�v ��پ}�.��2%	y�^M�0A'N��:   ������aș5^�˧p�q%#�;ؙ�r'I��TkϾ��{�w��i��);;{H��B
�B��MӔ�����������>2>�c�������ե��Nutt���S���.��c�m;P�j�D�f�$���
c��h���ɑv� \�C���=e]s��IF4�f����L��VZ��LS���R�@��|J�7eݯ%�t{4�O��s{�\97�*���ڿ���ws}?gN�f?�Nμ�>�á�{?#W~�}�3))��<S���+���e�$}��?������j}sCR�:��GU?zD�H$%�e]}�J��2l}w��L.��G�;�ݭ��&5�#+[�~�\EI]G���e]y����V�'�u�_�AM�{6��8�@�&~�r�����央���U�7_�7�.����>����Um[�Jj�3)��ߩ��O��ϝ�ٿX�ݷ]������  �GZZ�fΜ��0
� g���K��fϞ�͛7k����   #�ȨxΓݟ)��QO��#=V�9{v��3WK3W�@w���ޤ��͚��Rٜ�������������g��p��v�ys:�r8����7�H(�(����G�pX��ݽ�B!��ϿO(���۵�p��l��L�D���i�\4U����t���`ʺb��C�{˝������fj�/����תu�)Y�����/n�������O���$�@&>��~���}��jz�y5����}
���&~���p�f���T�<��W,Q��3%k�37_��ܠ�g~����Y����ׯ��]�á)�xXۯ\�XG{�r���/�������5�����Wu���Hc}�3 8{y�ߣ��׫���r~g~�&~�k�Λ.ש��W/K��H([8`q����M��ok�]��T  `8,_�\J$JKK�#E�' Ǝ�[�j��٪��Ԛ5k��c�Y	   ��P��1�tz�.��p}��]-V�9g�;�����������o����5�Ѧ��k֬Yr:�g}�H$�H$����nl6�LӔ�f��n�i������޷X,�h4�X,vֹ��ɓ'�k������ ��k�zʈ)j�D"��͐a��:��������B�(�8���5푟h��ש��;I_/�On�1�ZV�n�=ʼ��3�s���45�o���[�J�Ҏ�e��J�}2�k�I�ݟLI�{��e���EGf�2W_������ͦ�ߐ�sU�C�T��+:p��վ}��Y M�-w&��=�d�����h��.^��7_KJ�3ɾ�#g<&��%r����
:� 0��X�B����D�v �9)//Wss�222�5a���   #�S�&W�d���n�P"�:�y1nf��f�R}"������ŭ�W��٥��&j���r��ò^,S,SĢ�jT]]�������K5����s��y�N�ҭ7�XD=uG�Ο*��q � ����0*���������v^w���}o5�N��Ɵ�8��6�I�!m���M8c�$y&�� ��4�s_����]��#���7k��.Z���7%uO���7eZ�2؃��I;�P9�s5��_���Q��������S2y��XV�~6)p `��������u��9��� }��v�ޭ�+Wj�ΝZ�|9�   �B�;�${Z�LO@=����:��0��K��/UD҉XD�T�Q��{��U��S�y�0a�
�>Ruvv�ȑ#*?qR�=N�+S��i�|B���Y�ź;n��3s��Q � �N�#�
�����)���[�R��<��5��nt3l6�%��5���!w��^�'*��3�f�ww[���������C�����$-C��SJ$Fč��ǫ��D�o�V]�Y�iĻCI;�����d~m<���las{��  ��˗���C�DB���2F��I ��i�Ν�Ї>���Z}���c�=fu$    D�;�,�ᖧ`��-U���Xg���N�/�����zI��Zt��o�Pz�E���
������9Kcwuu���F�mlUc̫V[�z|�r�-�{ᝒ�1j�i������˰:
��m�X���#^ۖ��Pbu���w�m������fu�o�lu�Ae��Z�	��>Qnu���w�Աg��s�YEҩ"�i���vݰJ1n�F���ɽ  �
˗/WKK�$)=}4��
 �UYY�q��)����PUUUV�    
�1���E�y��/W<�:QR���O_)M_)Ij���jO�	�S��厴�ot+`�(���k7����������@  ��/��3�.�HD���
�B���Rkk�Z[[��ѥΨ�΄C���(�͖+�T���d��-Ir��m,7����t����P����ʻ���x�t������i�w��N�!W�8�TUX��=-]Ӿ��L��]e�6����߲4�i����X�����I���?ҴG~bu�^��U��t�߾nu �w�T��X  `X��~�������r�\rq�-  �k�.�7N;w���ŋ��SOY	   �(p����]4S��*E�ꬎ�Z�]��Ir�L�J����E;�*�ЮxE�b�f�zN*���n�C�]���Q)a�tyI2l.�l��l�	��2d�͒�|�ː�O��>�$�1����p��Q � ��Z���>�(E�:rH��t��|�Q_��.�L�;Ύij�7�{�3�D������J���9�$�O?����W��۬��TM����������VG�UpϧT�؏���0��{zt�/�S��cVG  V���WGG�������q  c��={t�UW���N˗/��   !(p��0mrf��ݟ���㊇CVG�K��B92
�����=�' g��c AZ7����
�\���Ųy}�|.g^�ٹØn�h|��ܿW�w���<�ΑU��<U�:�9�sR�cɸO?��ˮ�d�D$���U���T��(��mI��a���{�m������t�|[�o���;��;}����:���4�ݘb�J��$�0d��u��Tѽ�ձ���Y?��Ļ��$w�DB���oߢ�G��БC�]  �.Tkk�$Q� ]]]:z��JKK������nu,   ��G�;.8��'O�E�ji�Rb�w���f��rf�ȶ:
�(�P�}��3����O�?�F���T�O���*[�{yK���8��LA����4�3_<���C]����a�ꩮ�ד��c����D,fu��k��Z7�1���׶˙Wp����fu�����t��]����Q����'�O?��|G���!?��T���U��:  ��f����T]]-��-�(�� ��ٻ�8��z���3}f{/�MOi���I'�$�+�^,���赣���P�'�4��( �-Bؔݝ�}v�����Eʞ�̙�����l��|�	aw��9�o�x�W4k�,���K�u�]�����   ��t�e�[V����rKL�A��T+8i��  ��@�������;b=�zq��r��4�usA�K�R�*:�t����D���z��/�o~Y�����ٶ����   P�O�.�׫d2��� ��z��W����֦=���t    b���(P?[���ry�����)�8G��)���  �q������)-�}M2�k_<Cï��`���p�9�+䍎[W���+l�k-��k<    L�n����~Ib� �V�HD6lP<�̙3�Ja    ��U9 �*Sp�<���e�ܦ� GYn��5Sh�#���t  �c���*�3/�k6���x�)�����V�M��-��TѮ[Y�߯Ƴ>�p#    �l��v��ࠂ��|>��: �<��+�Ȳ,����1c��:   @�c�x�e�[Z�`�<y��L�A�\n�*j���  0!�����NJ��?ߢ�eW;�(w՟�9��F"2��W��v��3嫭w�   �BUTT�ɓ'+������g  ���k�)�����N;�d�   P�p��;�p'͕���td1˲�-�V�i����ŧT  ����wה�/I���_ӛ߾СF����c�o0]#o�-�Zc�6[Y�߯�3�u�   �B��.�hxxX�T^^n�  ������E���Z�p��:   @�c�._P���
6Α;Xj���eY�W)�4_��)��^ӕ  @��V�j������z">4��_=G��a��.��U��g���7���z�m��O9Sުj   (D��������L� ������r��������   4܁q��E
��R�q�<!��,d��O�'�TY��  &��x5��W�W[o��dRo��W5�����R�Ȉ�l�I��8ئ��/���.������Í    �y��ixxX%%%��  �غu�$I6l�ܹs�   
�M.��u3h�͠{��,K����ol��>  �~S���*�}�r�o�u�5�n��7����me=��9z�Í
GbtT[��{����g�[Y�`#    ����R�PH�d�w �������٩����Φ�    �w E�@��u3j�/oi�,�����r�[Z�`���&�c;  H��NP���R���G��W�:�(7�^��l�Y��,��6��}�uko��uCj8�\�   (s������\.����L� �u��)�i��馫    ��\`�,�_���m�����ӕ�&���M^(_U�,��t%  �G���ӌ����kk����d<�P�����=��l��N���O�h�B��.���}N��J   (;U\\,���6 �Z�~�,�R$�����   �)|�N��#oE�B�䯞"���Cr�eY������v��� �aSO1Ǉ��SZ�ٿ�Z�@��5�XT�v���]6��x\m˯��o8����������;T���>�p# ����.n^�  �f͚���1�� ( �7o���6mڤٳg��   ,�7�t�\�T+�8G�Is�-���r�n�q�<>�*l^ �����+ ���cY���㌬�u\.��P�yJJ�����h��'*�{«�)>�o+[��O)8c�Í
GbtT[����|����SZ�`# ������z�5G��;f|]  �^~�_������R� p^<��o����^͝;�t   �`1�8���W5Y��寙*w�]E��e��)�|o���Yn�� ��ب����u'�*e�(ow�H�Gk+t��Y�_�X����5��R�M�:S(GŇ��f{a�R����N�7h���.��%��y,>d�붷�V�|��6T�h��ll�ރS   �v�a��������� (6lP"�Ќ3LW   
,�<�U
4�P��*����nU�,˒;X*�T���$ʹm��[��j  l��診��V��4Ye{��F�Wu�r�{د�ε�1�x�.�t�S�fx����ݯ;�(��^���l�1�婨t�Q�H��i˕���o8�\vq�T�o���;�T�|���S�Q'��F;���1� ���3g����ٽ �Qo���,˒�����   ��by|��)�8g۰{U3;�;̲,���U5+ؼ@��Y�WI��  �%�f��l݉�w3M��EKm��·�ܕ;�X^�f����n������������8�,w�nnQ���j+�
T��4������^R�����p# &<�F�Xo+[~���kp��{*=���M�57)�:�  LԎ;��~
  s:::��߯��V566��   $�<,�O���m;�7͗��Y�P�,������S\)�T'�@����r{MW �1}�=�H�F[��C������B������b+����k��p#3���B��ؿ �����"-o9W*�]��l���dyy=�.��1m��W��g��.�@�
���V�r{Ts�I�yO�"��%�
�Y�l  0a.�K���J&�**�t\ @fmذA��ݚ5k��*   @Ab�0����-���n�BSvR�~����ry���˲���Wޠ`����_3M��*Y.��� �ӒIu�bo�s��U�1�.�M�b{��KR��e61��xU��씮�r�����_j�?��xDC��d+뫭W�aG;ܨ���Z�ѭ�me=�e�;�Lg0"|�
%��le�N<Ur9�����*�c[پ���e  d�wv�r�p*  ����okttT3f�0]   (H���r�,���Y��y
5/��f���5r����e�wڽeu
��ܶK{�y+��I�e�"  F�׮P2���[���.�_�G�`+�����cJ�g�����v���h�o~�`���v�U���g��`��F�����7��y����7���e��&�l�O:�H�[|���9�����  �bڴia�v �---r�\*+�dB   �܁,fy|�W�W5Y�Is���u3�+o�;X"��1]�q.�O��
�*�h���נq�|�Mr��إ �koU����ă�g�d�=�Su�Q��ʆ�ܤd,�hS�N\b;;ںE�/8���
�:�\�hg�V�h�B�춗Í
Kx�r�n�d+�)�P��'9��	���mgS��8�ۣ�cN����������  ��ԩS5<<̀; ����.(�ɕ��    �_�O�y�r����*��_KƣJ��(16����(�(�L�*���������C1� @��W/WŁ����-Z��g�t�K���ɤ�kV8��$��Uɮ{��&�1���s��v�U~I���}��j:�"[��3���?�p�U�Hƶ��>�~f+�pƹj[q��H8�@&�>��F�n���i�l�!G�[Y�hw�#]*?}�|5u����Tbtԑ   =��
�LW �M�6���YMMMjii1]9��g��#^Zi�F�y�a�R9�t��I�܊ox���T�*�l ��[�N������IG#�$W2��_��p���7��29
�8��;�;X���I�u¿    IDAT%ccJ�ǔ��n��ؿ�U2��R-�%����������ey����Ǘ�N  䛞��Uc�6�j���V~�6�������#0u�Jw��Sv���P�孴w�Es��ʶ^w����Í�S�Mת�/���������
4OQd��hV�koҤ�lk�50e����G}O<��f 2&�Px�
5�x���zU}�"�^�GG��.��C|*;�  3466&���  flڴI����:u*��-�+���-��k8f�[jj�u �Ow�7_a����sƿ��v%�����.9�w Y�,�_n�_
�|h$�)��I񘒉����{��D|۠|2)%��Lķ����?k�dY��ro�����w�{�@�ۻ��{  pD2Sǭ�4��/��u�:�X���.�=�-�,�V6�zY���%;�n+����z����_ѮNu�u�j�;iܬ�v��Գ����9_�@$�Qm��4��?���8�p܁<^�LM_�@�{�?��-Z��k/��|򜯡Qe��o+;��S~c]Z�  �UTT���"y<��	 0���E�x\��ͦ�    �e�  3,�G.o@�@�ܡ2y���-���bҶ��&�W=E�����N��v��������k��_3U��)�U6�[� oY�<%��U�(��`� �
�����X�"����ey��9v��l��G��ݝ��"�<�Vn�4���p�����?��}_�x��%��a[x�
���ۅ��Ӈ�~ @�kkU�#����T�.{��C݉Kl�KRxU�>` @��:u�"������Hr @�immU,Sqq��*   @�a�   �_m��>q����孬��1�0����V.�:��=�Mo����T���f��-T��z�Ŵ�_yС�VU��vܺR��Ѵ��m�Q���M����Wm��w�����5?�����n���\|ɸYc������|Q<'�->-����t+�Ѯ�W^Pbl,�������*�� [ٺEK4�̓�[��R��'ۊƇ��u��[  8bڴiQmm��* ��H$��֦)S�mf    }p  @�(^��&�[*��9�p��#��W/�5�+I�'.�[��f�֮]��v6�zy���F��
[���N����믴�����sԶ�j%�q�[��[Wiʅߖ\��3�w���U�A�:r���z��Wm��eyc�#k��}�=�v�����c��'�(�ߗ��+�?H��I���w�Q|x(-�  �477+�+�� (p[�n�����"���:   @���g   �4�K�/���|����dN�K�vUϤ�{�=0Vs��r��f��a�����Vv�٧4�ƺ�����6��M1d���E�������ɪ��g�-T`�]|�y[��snw�H�G��n{@S.��,���m��:n_m+�
Tuıi[�vQ
حZ��u �sd����  ����Ujnn6]   ((�   ��\���Ԥs�Ϲ�vI���A���2�f"Q�kme�%��:쨴�[�h��B.�l�d-II%nR 	���'��3�u�Laz�ހ�����&@a��5~�?��ﮕ��3�!�j����u�nђ��魮U����^���q  �9�e������ Y��'O�l�
   PPp  @V���o���Mט�����d�n�+o��Mǀ��v�渓le��C���^�w�57)>�o+[��>*^��Í
K���i��R�� ����C4���y0p�75�̓��E��h��^����ey�����>  攗�˲,�U  PGG����T]]m�
   PPp  @�*��P�������R�uWY{x�+z�[ْ��Rp���Z�|���o�d+�y�Ň��k=��ć^s��|���lSxb��.p3�8���Uk���tk_��v����|�βT{�)����p  ̪��S$a� ��ɤ������MW   

�   �Z���M#���C2�����C��:�4`v��ᰏR�x��lxղ�Z�8�7\�d<n+[����kp�Q�p��r�ш�M HR�W�!������oS���V�������Ô��I&O����m�  f���2� �*���r��
    W1�  ��䩨Tپ��11��6����}��5:�\�Dd�V�������&����V��d+;��������ݲI=��V��xUw�i7*��&[�X_��M H���A��u�����V�]R��Î��Zu�Rx�n5� �+jjj�r��v�MW @���ѡD"a�   PPp  @V*�� Y9�Ff��O�}��-��t���u�����
Ut�֩=�TY��l��&����믴��;�#;��]v����t9��;*>�#�S8E�nђ	��)�P�����F6���>9�u  @�UVV*��)/  �[8V$QII��*   @��.   ��Uy��9�D���(>8��GR�W)>�����I�v���^��ޤ-��Z���u�^�L5�.���]���@��,K�ǟl+��D�y����ۂ�g��#�g��/�X[k�������Kϫx�N�f��U�>��W�����Vתx�.��C���p �L�ad������+/�h�q�%�����yc}Jk�w���g�W.��ɔ�  ̩��P�� Y$kttT���Z�n��:   @A`�   `�=�y�U���������V퉧ꕳORd㛎v�VT��<�O�?���]>J|hP�p�F�zS�/<�d<n�����	�����3f��-�� &OU�e���������v�s�b�}����οHM_���Sڗ_�S��v�4󧿶�m8��m�3�8a�Gc�����/:�Ȝ����M_�[Q��C�7竪�@�^s���p���N�ۗ�OJ��=�[�d4���V�to  `� �l3<<���>���2�   d�   ����/��p�;��M��ez��O)q����K��'Q�e?v�G��IS.�d��e�������پwݢ��{�f�l'4�y��Ͽ�t�����[4�o�[];n64s���}0��e��3mE�]��l��h �Z���ȺE��p�����p��֔��#W 8n������?Qbl�ֽKv�S��;��v���]���  �<�˥��b�㿆   �:;;5u�T�5   ���2]    ��]\�Ƴ���䩪=��5���u�����l�	��ޅ�S^��Of+��������,�󔖩��_7]#+%�Q��t��|��:�&�Up���f��v�w;�">Я�{�l+�)�P�A�ھw���[�v  䒊�
I���3� �������   �A�  �}��"��c����7m�ѮNu?�[Y_]���;�V����������ju@���*2]#k��t���������Y7�OM_���l�_�t�	�l^��v�v�[9wI��;�Vv�u���v  `^}}��ɤ,�2] �������ɳ    ��   xOY��\y��M�NN�՞p��\2U�m+m��<�U�+d�hw�:�\k/lYjX���C�ⅻ�ʎ�nU��:�@6��1E��`+[��
L�:n����
mݳ}ՍJ�㶲   ;���0� �J���r�<�   ��c�   �Ǜ�y���h�[ي����c3%����ٶ����_�괕Ej�a��^뵗�>=�渓�)�p�Q~i��mg[��R�x��6 �N2�������c��=�ރxJ$�q����   k�;.  +uww+�H��   �  �B�H�c��3��w����.�^��v���q�L��jï���'��u��[���F���CU�`g[��Р�W� (D�+��EmekO8E���W4o���.�u�����p  ��PH^��t  >���G�x��F   �a�   (�)����-^*�>���RUv�����nU�c������W�����Z���v�~�ٲ<S�˲�|�E��m˯U|���B �U�3��﷕��5�|��>��Sy)�C5  �P($��o�  ����ӣP(d�
   Pp   
�X�V�=�����i����ć�X��'�ںO*C�����Ҧ_]�d����o�j�7me}u�:��7�}�j{��ȰZ���Í d���嶳�qJ�+R���ٺG�3����g{M  �=�� ;� �Vgg�JKKM�    
��t    �^�\�8�V���%�{��'�jo�DBkW�����Pǭ+UqС��7ھ�a��r`ǡdR�˯��o��V���/��Ϸ8\*�Y�&}�����R����B �]�C�k�u�|���8�`�j�5n{�ǫ�8F��[�׮P2ƃ_  �P($��g�  ���G���jmm5]   �{�   ������j�l�g���ʪ��/�����==���-�Ԍ�nQ۲�S�����
c�]ۆ��t�<�e�f��-T�.{h�٧2�,�T|����d+R뵗;�@�K���m�&}���f-�G5ǝ�-���}����?�XR�5<` @�bw @6���W]]��   @Ap�.     s�Ѩ:o[e+ky��>��}��p����e)u�Tx�r���3�u�M�,5�煶�m�_��� $I�K���lݢ%��o[g�R�λۺ��Gy{Ä:  ����(  S���
Ɔ!   �i�   �}ՍR2i+[w�����+R��ں.�ա���7�~�S�n����l�!G��4��F���#U4g��l|xH��_�p# �bts���x�V��4Ye{}�����G�^�v  ���R�  �H���
�k    �c�    ������{Z%��1n68}�Jv�]�=��#�������5+��E��*�V�[7���{T��ώ���n՟z�����3�,GX�&}�����`�v �^�\e��g+[{��=��\>�j��D����U�}wmOE  
���3�q��k���t�_m���|>���  �>���r��)]�,*��7~�P��]�}Y]��   d
�   @
�^nk�]�j-��sO�n�R{7O&^s�v���v����%�n�i���_8�(wT}&����z��7�k��S�z~$OE�٪����U*�� [yI�m����[ ��PR�De��K$�Sۍ��� �n`` �k�.�)~M���  �l�2]    @�u�u����_}�1*�uOﴫ�|ߓ�*����8���'4��s��������F9²��ůَ�^w�b}����Ѩ:�Xc+ky��>��-�������+&Z  d���"�  �X��æ+    �w   � %F��y׭���`H������^�l����h��O���g�'�ݏTu�Q
�0�V6>Я��t��\^��v��/�t�}le����^{y��  @�z�r��/ @K&��F��k    �w   �@�2`�kh���������&Z	Ȉλn�XG����i������FY��R��j;��� >���W5�³����ɲley� ����xp d���Q�   ���1]    ��/<���^Vќyi�gǭ+��D�v?�	�hT�7]��/�V�[U�p����� �-�z���Ň��u��i�  ��8�����5��E)�].� ��766�R�eY���t��{▥��    ���   @�X�"��8�}�u<�aG���o��
���, t޹V����  ���,�����X���x��7  �E&�=E����_   @��U.   P�:n[�D��Tx��z���+$�q[9���t�����X��&���R�kL��zՇ���me��jc�v�)����Q|xH]�ܑ���W-K۽  �9n��� Yoxx�t   � 0�   �X_���+-�b�����]�r��F��|8W0$OY��l����6f�^w����ޏb��j���l�^{9��#�X��N>C;�����������_��T8�x��^����U�/>��{  ��� ����LW    
�   @�KǀY|xH]wߞ�6�#��a+Wq�!�ܙ����%G�&cQE{{2�(��X���6]#k՞p��3f����������3ӿ�SM�ޥ
N�)Ir��d�=4��?�nV3~�K�]`�e�x�)��n���~�ih  ����3] �q���DT    o��(�F�u�-g��K�	�+��� � ���c��k ǹ������?iyK���&|��;oQ|�ϣ��h�f[9�d5�q��^�{���SQ������X[��H8�Ȝ��Tپ����uS�k��/��o��r��ldV�!G��������W��'��������j��O����J�cl���kn��o|o��'FG�yǚ�  F1� �ccc�+ ���u���7�s�q6*���  ���_*�v����t��]�dB�C�yT���k  �\�L*��fM��7'|���ei,��}�vv���dtL�ˮv|�<�<E�s���M����<�h�z�O#�xw�fHe��Y?����%��^voGީ;�t�����V��{k�u��n�V�nT����v��㖛5����k��l]�C���4�  �x�^�  �@nE���� ���16��6�5�  ��L����K�5G��[&|�����Ur�B3w7筮�p��<N��w6]�]�xL����q�J���:��W/W�.��N����_ͩ�k�>���:�嫩7k�=��������s�=mk����q�B*^��*92�A��Ik���L�m�՚���nb���Q5G�����r��qOY���4��9�u���woy���濫��g�5T|��b�_B�wL�_C�&�������G4ڶU�3'�x+*m�i�Z�n������?zBׇW�  ��w @.�g���  �|��;  �u��j�%?����w��F�3�^��'5�?��t��?�Lm��j��G�������T�Ϥ|m��h�����o�A��_d����l=��)c�[���{M�p\x�Mj����)+7]e\5�.����L�@ -��^��������m��؄�u��*���4���hW��6^�|Bo����h  Lq���� ���FeY��   @�s�.   Ph��=@ӿ����� �Ҥs��Ƴ�h��m���S�&1:��;�8�&?�^�E;���T˯~�D����(�&����V��A���_�e�=]6���ގ�y�-��bt�&����胊�lL����˥�3;�  3���
  �ktt�t   � 0�  �a�_�Hr�2�P4�"��KLװ����i,ܖ�5]�C��^����6��2�5&d赗�q�j�52��ƫ��O|��L���K������ն��5 Gtܺ�t���}��ƗL��U�]����� @�`� ��Ѩ�
   @AȞw�  
����d��L�@��!���$㱔�«�9�&���N���t���������J4\0�u���z����ؤЬ9�k�+������d�7���:�X��{�4]c�ć�}�=�k�^�\�x�v���{4���`#  `B,��  I���
   `�p  � �ϟU��n�$����)�0]���eR2i+i٨��w�QH&��.��ϚnbK2���|N��ofh={o%��۷^��kL����t��$�p�Ez�%�M �$�q�~���G�V���t�	�z����1]Ö��V�=��|x�r�   Sp �W���   d;^y  dP|hPѮ�5�"��m�rFd�&�l�lz[}O>j+۾�����.���/��?�0]�cŇ���+�ﱇ3�f�3l+7���pi��'5��s��3c6��H��oM��6�p\2S�W�w������g�4]ɶ��_��k�`�FJ�W�h+7�u�z���e  �� r���6]   (�  dX睷������p��M|k�d�o>n&�ݥ��g�M��vw��3OTx�M��|���V�|�q��;�֛��2n��o�f�M���>ֺUC��h�C��[���T�+�� 2-16��{��K�����V)16f��G����W�[�D$b�JJ��������p�T  �y	�� r���1]   (� o��s    IDAT d���_�Ȧ���<�v��m��]Ȓ�6|�J�sk���W�]�}t ��Ɵ\���@�J�d4�7�u��_p��Z���#i�����7��c���/(���?���F�׿������u���ed�Tm���|>I$�y�Z=ܧ����_�"�/<�7��%=s�.j���m�b����=��^\t���1�J"��?�D�h�##�<��[n�`)  �I�� �.c6   @&��   �b}�zy��{��UR��E����k�w.2]%덅۴���rv��o���;�H���>�������Äu�}����^z㿾�އPbt4�"-o���?�#�ӆK.R��'�����;����C�^~A��{j�~����ږ]���R���Z��s����z��^�-�V/�^��kk�Ⱥ@.�vwi��ֳ���[���oW|��X��7�i����+�q�b}��zl��'���U���?���?���OS27�  d� �\��;   ���  `�X{�^9��v�������4��@���|LѮ�����{��]�?NbtT�������F���%�����S[������W���n٬������f�d4��[nV�-7��t��嫭���^ުjY>_Z׋��*�V��SC����o���۫m�5��U~��S�)�������{3>�ؾ��'5�|���O9�����[�O=��C�Rp�l����;1:�X_���6����׿�s'P ���������y�~Yn��v����孩����ѵ���i���iy�ѵ2�������ê��a
L��DdD��S�O=f�  pX"�0] �qY�e�   Pp  0hx�+^���Y��ч���C�k<~�fFbd8gw�O���V�^�G�5��ֆK.6]�#��zվ��5 ��d<������Kϛ����C��}��   Ò�v�  �����P   ���         ��h4j�  �����D^    0�         ����Y�e�  �w    3<�          �O (����)޿��ߡ&  ��/ůo��J������J:�
   �9�         �����q�mB�ǝR~ddD�h��^  l�˕�����m��   ��p         ��444d�  +�w    �+o          FE�Q� Yϲ,�   ����;          ��� ���r��H$L�    
��t          �3��;{�g�ش5�kh @z����tMrdP#��C�ޓ��r|    �p         
H�G{�QgאG*�O隁���  ����FFFR�htL�w�u�   ��\�          ����
  |�`0�H$b�   Pp         `\ʻ� �A�@@�d�t   � 0�         ����A�  �H�   �À;          ���,�2] �
�LW    
�          �koog� ��JKKMW    
�          ����R45] �UTTd�   P0p         `\$QOO��  |����ň   �)��         `� �lUTT�)#   @yL  �A�z�jL�      �.U�a��M� ��666���^�5  ����"��   � F==e-��k      l��x����L� ��ǀ;  �B!E"�5   ���2]           $����t  >���H�D�t   �`0�          +������-L @v)))a�   � �;          +lݺU�e�� ��,�Rii��ɤ�*   @�`�         @V�����Ȉ�  ������E   ��8         ��0::���v�5  xWII��Ѩ�   @Aa�         @V�D"���2] �w���hhh�t   ��0�          +D�Q���ɲ,�U  ���   �	�         �7nd� �5JKK��L�    

�          �ƛo�i�  �$�׫��"%	�U   ��;         ����۫��n�5  PYY��    0�          k����t  TVV�h4j�   Ppp         �5������͎�  ����588h�   Pp<�H���*�Î*�q����SR*W0��بb}}kۢ��^��+/*12l�����%�:��*���ܡ�"-�}�5��:��l󔖩��Ϫh��m?��-������Nu'�.�dc��}�|�9#k�f�Q��G+0e�,wV|��-�թhgX}O<�����d<n�        %�H���E�쳏�ɤ�: �VVV�����S d7�d�]���9��]T,��*�ӭ�u��*��m��:˲T��~*���VV+�ۣ�������	���q�T��U��'孨R��W�O=���ߧd<f�R�N����Í�mJ��-�W-3��+P��Ǩl�}孪��ɕ��䶹��.��N��Oc펯j�W�x�]U��4U|�<e�����z�_�7������Z�?���U���x���}Ս���o+16f��=�G��i���<�e��x����U��݋��|����=����&EZ�������h�~���O�\�}@D��hw��n���^�Ǽ�       �l�a��\.%reP �w�~�B��LW oU��N9SՇ���ٶ�|�9u�u��+oT|(�N���k�/.W�n{���g���W_���������'0y�f��
�]�7�y���X��_=G#o��x��y4��3��I}�>dd��d�=5����o���i�L���G�rُ4��3�-cd50y����z-��.՞p���vi������ڕw�d�=n�9��>L;����K�\.՝t�f��jYnw���T{�ɚ���~`�]�dY�9v�v��u9��7l�,ͼ�ת?�̜n���J�_��v�ˣ*�� �u        (---2] P�***$���  ������oh��>���/�=�.I�v��o|O����N?'淪�5��nGю�`ŝ
4O�p3���M��nGh����v���p3dJ�N�i�5��c�]�v��^�Ђ֌�R.�ϑe2�Y��EZx�_U��l�}��y7�U�^�󟌽U5���ߎ;�]q���_rv�Z��Wנi��T���͕�@5�qn�Z!��?Z՟=�tG�j���Twʙ��        P������j� ��UVV*��� (��35��j��r��&|OE����4���Vצ��3~���&l�SQ��?�ݸ�������~�������\���瀉�����o���MWI?�R��'k�5�䩨L��3:�x�4����]T���Yn���t�f��szȽ~�Y�M��bV~�[�T�@�V������/|��,}�"],�Gӿ�S�.Zb�
        yohhH�6m����  �TVVjxx�t @(�q��/�]Es��e����n��.ww�͚����-�yw�캧ÍR�9[e�`+[�`g�Í�ie��_�)�M�pT�n{i�U+�
�zߌ}G�~�ٚ��:r��N��o��#�΄�}�����7d�q%��m;뭮Up�i��R�N��n�ӿ�S��        �H$�6���  ���v����� �N���׭qd�����{�j�KJ�~�L(���)�q8�t7�s���K�C%c��h�BM������p/�i7��N?G՟=��5���Q ު��L�xGh�;_����Y��ay����W0?_        LY�n���� �TQQ!�˥X,f�
  ���!�����9�Fp����e���IޚT�*S�ā��*S�9#����MWȘ�c����xpw�u�ey��v�Oy��i�۝�Yx��J����8SF$"#����1�)�Uw��k        ��zzz���f� � UTT(�L*�L�� �cS.��B3wp|��C?����:�he�\ej�R��D�����Q�/�v�����ѓ>w�����^F��)-S��gd- ����æ+dT퉧��        @^���ז-[dY��* �S]]����5  y,8s��N9#c�M��;r�[��gﾣ�(���gvWZ����;��	!b:�@���fzǔ@$77=��4Bｙjl��C�M3�`l\e��ZI�]i{����}!ZY����H���99'ڙ睯�������4��]�#�U��#���eh���ҁڋ�4�CT�q��zM":�PU�c�M��}�[[ov""""""""""��������yN�#"��e�XPVV�P(dv""�`n�=$�5m��W�qg_����N����yw��1Ҫ��貎���^tE����,V�]vMZ�ID�w��h��/f�H��̎@DDDDDDDDDD��TU�ƍ9����Ҫ���,#�����2T�>������~ݺ���%� ��%�vM����V�c�M���uYǰwkY9�O?ר����'�"��єke����@ӍW!��4;JZ�*fG """"""""""�hN����f� "�,RYY	MӠi��Q��(C5\}`�ֲr8N?'��%�vѾ|5�x���PU���VQ��:��qQ{�¤��Q#�W��p{+r�ǡ���ב�6�]z5�������� Բ=���&NA�A�$|�����եB�*x,�EB5f�}y1�^{	E�9y&�ZRjv��9�{㄄Ϸ�W������������000������P��K`""2_UU��0܉��{�D��&U�]�9|k�@��Pr�ᰏ�$�F�E�|�Q��PR(��;��ye��K+���F�[���K���`ƾB�0C�ݏ��/Ď���ki�ّ�7q2j.�<��e��U��n-+Ǹ��6c�eg#�Ѷ�1[Ef<�
��)����3�~�-�tu
� �}�i���8����jp�y��7`�r��hp -��'�1��j��)���B�������������� x�^l۶p ܉��p���(**���1;
e��+.<�]��t�p�����$��?��^�Ph-[����F�
�@`���G9/_����;�[�&����1��K�����|�(R2{�P��$�C�!ݙ��_&<u]�b�Eg|����/s��B�֓l6�]|�P��h6l`s;����  D"��Q&*��ʏ>N������Vs; h�����Qh��.�_	9'G���(�top���b܂����	gW�cg:�GxMǩg!�1N���������������F������C�rHDD$�������*""2D��넧�{��=K��x��� ��ʩ�Aռ��j���M����.���H�&����'�xN��!68 �����ڋĶ�  M�̎@DDDDDDDDDDDD �n7�n�
Y6dsj""" �,˨��D0d� �.�4T�C���n��w)�u\o�*�n���@�ل�(��%�f�~
d)*Ƹ�/��|�n����Q���~�!ᵫ�89U��u�Y�W�|�����B���DDDDDDDDDDDD����ASS܉��P����Z��BfG!"�T����4�������#��~�M�S�kjQu�iB5�yT�O�|�!��b���d]?�9�RX�K�jb�~8�}<�s����^s�eB5�y[7���y�AI�ܶU��P�6������hjj�����"���2Gu����h��$DD�i�&OE�q'
׵��Fl�6���k���]z$�U��2G`�X�����"v>�*���-�E�9��·�d��� �O="|�qg�[y�pe��eK�Km����08��ޗ�O��`��7o00Q���nl߾�S܉��0���@��KDD4���?�޾a�５����Cx���a<*�"TC�ſyC�M�j8��ז�H���U���;Y��Z����H7�}Ts�����=nt?��PM�#�B�y�j�|Ԝw�Pe���M�N��%�ǎ��?iH$ν�-���|��4EA���:�����������������ۍ��&X,��Q*))A^^���4%�>~*���p]��7��6���{��S���8�=�i���+hJl�S�n�"�]i%F���й�瞀�z��^tip��`�9�u>z�O�&6�A�����5n�����
�Q����ߣ照�=���shڜ�Tb�n�
�wW{\�F����c`��iLEDDDDDDDDDDDd�@ �M�6q�.��� �DLNBDD�fg�؍�����_��ڒ���8'�7�S���Cl�~!�P0�	���{oE�Cw�7���W�b�����{��W��ϿNc*J�.��ξ��
��;g���|�^��xKaj�h§̡Ţ��?�a������K�� ���:t�w���~���{���x��h��5�]��������K�j��������������h�r:�hii�,�I5 �����!�����2��q*O<Y����Fu lݔTc|��|���\�_�'|��܃�����jmF�K�c��?D�5;∺ ����@	�{WU���ϰ������K��f�1%�%�|Ԝw�p]�c�#68��5c7�=��K���9�Rt=�@�ץ�0�����}�c$OU���s�}�9H�|(>�٩��������������ߏ6`�ĉ��NDD�)--E~~>���Q��(��_q$�X�fp�V��|-�k���O�s< I	��M����N�k��I_�ƾHW'Z����$���;a[
��{��N�[ʷ݌;�|�**�j�]�?��u;�G|�{Q1�-�0���&������������������������NDD���� �B!��Q&ɭ�G��S����9����7�On���?�w�(�����1.�g$975�_&\��ă)OQ�y��~�Qẚ�/���0�kQz��
�Ӊ��f�l� ""��jp�D"&'!"�LR�u��6��P�v��������	h�PM��i;'��)}�S}�ȩ��Q�t?�`*�ݭ󡻄��[KJ1n��\��������������ҧ��_�5,��Q��(���!??�p�`# �prk�Pu�i�u�wߢ��i��up�zS��~�� IJ��DDzH��]��E���u=����d/�-1�Χ���p!,��d """"""""""""��p�\شiTU5;
e���z ���79	e���
�&8��u�^Y�[��;�!<Ž`ƾ(;�X�2�"�����E�c�P�
�����d\�% �F�ZZ�����5+����۷o�,��Y5e9Y�QSS �D"&�!"�L�SS�������VhJL����~�-Ẇ�o�w"���G��A�E�뺟~QW_2�V���3ILq�x!d{��Y��������������X}}}X�~=,��Q��hs8���A8�&8ᖈ�h8u_9'G�&�Ձ�e/螥����Oq�g?��9J�,DD��jpw�_����5F�#�Noߥ�;����*�P=�!y��������������.��6m��(�8Y����T__ ����M�����SUǼ3��:�Z4�{��up��B�����랅�H�p��d����+�/�|�qDz���s������u��^�n7 AQ���`۶m���yQ���lp8 �H$br""���#F�:ѳ��m��Mx�{�����JDD��O|�����z�5A�Cw�^JH�wC�jr���8�������v�ZX,���T__Y�
��	6��c�t�z���u�n���]�_�{+������4DD�jp��6�],>����E�8���DD]�p>#>Ž�k �l$""""""""""""""#���a˖-�����NDD� �@��$DD�)�.�R|z{�=K��޾K�m��������%""�U�d�)�#��Q�Z,�·��IVǃw���s!���ɩ��    IDAT������|�I�Q��,X

u_W���)1]֒sr�F"��e�5�vQUu��C9������ƈ��rA�4D�څ�v�eX�t_V	�������u������ħ�w��PȀD����+x>X��9G	��_�3l��4�R�Y��Ն�K��@ϒg�l�KF���g�@�y�
��]~-z�<�ۋ	"""""""""""���	�����UC!��y������ְ�����Eep ���Χ�5g�������RT��O?Ķ_]���(������/����
I��	N$$"��4~�x ;���o�S����~���j8��Va���HOwRk���c�oA�����������=��>�|4\}�%��}����Z�Z�u�F&���*X��j��^8�O�P��;nnp/9�px0��lP*"�DZL�e����<�d��-�Ţ���P��|�.Ớrk�Qy��%""""""""""""'��8�DL�����%���z�ߝ�b����~�W���2V��cL���a--�d��d�L��aH�n� N?����c��r�_{Q���AMM  �������������^w<$�U������� Y����b�/~����[Ʋ#�������
H�<��y�ͦ�52����g�'\����i�޾�w���|�J��.���D�Y�ťB�!}^g'�Ws��	/���b��[��R�u&ugS͹��������������(5%�� ��V�.��M�k��s��k�Z?:@�`���7i�n� ��ip:���/`�MDD����zȲEQ��̎CDY�h��7i�p��q"
����z������f���SQ�����P��������p>��A���~�M�5eG���D�9��:?����	5�pP�?�{�)
:�3�P���ớ
�����lP""""""""""""��I���������W�K5�n�*�0ר��D{�t:�q�F�ANq'"�=�$	&L  �|>h�fn "�:ɽ��=�C��u�^C���K�1����:�J���x����+�$�[ >��2�d�	�T�h���	�լ:�4��^Y�Ўm�uz��:ѳx�p�c���!"""""""""""J���O�l7;Ѩ
���ߏ����S܉�h�������`��"�t�o\����f� ��tr��jb7��zԘ@	h�S|�{�ON���c@"��/���	B5��u�vB�e�#������[�ɣ����Ք~$~�EDDDDDDDDDDD��
���l��R���j���X�fdY�$If�!"�Qj�ĉ �`0UUMNCD�B�D�yo6_u4E1;����J ]����3 Mb�k>����	�X
�P|С%"�QI�Pw�U�_�3�R��:�	�S�#��VhQ���l6gz�.g��� Ǽ3�����p��]�Ɉ���Ge[�J�������������E��hf��1�2���BWWZ[[QWW�X,fv$""e���PQQ ���&�!�������Rv(=\��]�F�|�	��$��Qr�aB5eG� �V��F$Ym��{7"�."�VQ���ĸ�.@��Y�KDz��߸^�8#vs}�{:�_�T�u?��P�; �̞�w"�Y�Pv�q(?�x�:��Jȹ�f�J��wS�N������|�	N=�T(�M�̎EDD�ȤI�  �X�h��4DD�	��%ȟ2M�����u��(q�V!��	y��$\S<{����(9'�.��3�?u��q�z�E@�ݒFlpϛ��Ђj8�{+��'��������	׌�����b�cޙh���*f��]����DDDDDDDDDDD��tbӦMp��(**��(fG""�Q"77uuu 8������7Y�� \o�f@�$h��xu�_�pIބI�l6h�Q�(-�e�q�(��;fGI������C��'�tB��B~�!�P0�@z�J�|6���ZZ��]�I�GF6�@����DDDDDDDDDDD ���࣏>��:�/""�"&L�,��4����g!"��Md�9 @�0��;ƄI��]�!ƒՆ����3%E�X0펇�Ts; �<��6����=��AhA���I�1��:����'��({���c�s�Q|�l��&68 ��5f� """"""""""�����ڵka�X̎CDD���jń	 �J�4sQ��w�!6�1(�����U�ao%QzT��wl�^F]�h��o��9b����Ph����I�1B�y������n7(Q���1���ao�`vCy�}Z�[��������w"" �?6���w"""���U6�$9J��H�S��RXdP"������B4EAӍW#���uݑ���bw�a����R�'b�dM��ߑ?mo�cJSt�{��1������������4MCgg'>����
Y�P""�`�,cҤI �H$�X,fr"""�$�}�Q����z����(-���AH�_��t_w�Ou�\��H$�0FP�a�9/π$D��p��Q5w��1׻�Y�6�����������()���lO���nG��2_ww7<֯_�)�DDY�����;{^�^��i����7i*��%)�#Y�ț2M�D�G��L���h����$JM3;��HO�!��஄�b�$���!W~�e���n $���
lހ���c�(���qKQ1*��������{�pg�kMUUtuu�>�$I��ND��$I��ɓ �� 2ʆ5%*����Q��Q9����/;��q���a�S�Njpl�U��Hl"��g_%Q:�Z��A���w3��'����~�Ђ��ʤ�!��!\��x�.�(KaJ���1qva����&"""""""""[7���˸Ǫ�/Hy}�0kx�|������'JVWWz{{�m�6X�V���	��� 49Q�������ǪO;'���ώ�x`�F�֯My�L6��*!I�U��V���D��믘A���{�� d�]�uGnp��=)�M��t#��5C�|5��;w���z$�����]�u�O�ݩDDDDDDDDD4��,~*��E��){%�n���(>��ǜ�/Jz]"=D"���`��՜�ND��$I)S ��
�LNDD������O������9�jP:�ȸǜ�=����Bt�n��i%INnm=,�b�c���7�-[2�ЊѪ`�>���j]�qdA��y''�`��Y)�[�	�ω"Dɱ<O�%�߇·�F�CwA�͎CDYJ����A	����P�> ��*Д( ː$$����^�^ k~��� ��#�,�)Q�|.(�A���ϗj,M�Jt�I$��j�l/�%���bX+ Y8я�2���P�P�PC>(a�h���(��B��v���� ��b/�l/����M��DD�}�^��_��8[�;杉���!�u��HҐ�� \�Z�ԚDz�����;��܌	& �WDDY���q��v�W����h4�����ֲ�!��$=i�q�Hː��p}�^Hj�ljo:�VQ�ܚ:��:J$F�� ���HBD�ISb�|���~ߓ(����qV{ѕp>�"=ݺ�7�7��m[Pz��	/X8� XK��S
��nGɡ���l4(Qfu��@Sb���Uo�w鳈��̎DDYH�qw :�5���ɪ
*4%
5 ���I�K~9le�SVɒ��mQ�QC~D���@	��\�BC� J` �n{�$r~)l���)����ott"��QcaDݝ�z�x U���ڮ��hJл�� ,�BX��`+��5����DD�%�G�믠��Ӈs�|�n���ζ�͆�Ϗ{��%P�����)��vcժU��� �2�^��'����횦!�!fD��H}�.Ÿ�/r�r�<���P#|���d�SΈ{���2N�N@p�V��Ï����H#���:_�n�aL""�Ӎ�g��qg^����#��Q?�R��Qs��h��uYo����-BJ*N�	�O?�l&ݔ�C��<���f6�%�Z,�Ŷ��G�f%Ө*��>D�]�bё�'"ҙ���kE��5$�İk������!ؾ��j�:&�ZP���DD�i@�Ӂp�����X�i���@�{��KA�Ua+�0t"%�X��َ�`��':(!����fX�Eȭ[E#�Q��*��O�mp�������'��{°CO��/J*#����P^^�m۶aҤI��ND�����O�����&"��瞌��n�/@��sѳ���J�������z��.!�m[w~�gw��T��Q��n)*F�Q?�	lݴs'P"J5B�#���{ Y�����JlU��}�^pr���p�r&Zo��h���#6�~����:T4�W�q�p��U�!�!"=N�����DD�����iF�w��7�h*��.D=]�V�^3�¡���F�D��vn�6p�(>�>,�Bث��VV+��$����^����v�p��������"�1	9U��ND������(�}��|	����lڂ�){9昿@���z����6o�ú�2appn�+W���ɓ9ŝ�(�Y�VL�:u�ρ w�!"}��7
�GScQ�\}»e�I`�F��}���s�_ ��^=�츏�Zw`𳏒ʘm���P��~	��P�O��@�f������`�/�`_%��T���/� ش=���߅��N���������~�픳���jmF���Ɖ	/�?u:ʎ<�Uo�.E�������	wu ��܉��(}�N��C��zݘ���հ�T#�~&�{Z�OD$B	 жJ ��a*!�-_��ی��}a�/M����Dh�����H�u�X�΍�� �~_�Ji�>�h'Ym8�͏���` �o�m����]��,y�o���K=��	��Hh���F��>,��g̟BG��v�؁��2lٲS�N�w"�6i�$����y���ӎfDD�^{_�F��^�&�n�+���t�ѳ����E$�4m��vz��'t�2��}[�� j/�M��ƠD#��6Ԝ�p]��7HCD��c��.����Pr��B�ų������X%��7����z�=5\s�pM�[�HBDDD4�����)��?M{s�7E��n\�h�����ivl�w��ion�&%��o�um�g�D4*E\�ܰ2���ߤF�o���5Д�i9��2�����O�~K�D��9��ٳ����%	U'���:է��ٵC��zui*�����r��r�J ��b19!77�&M h����Dd:�nG��s�ߒ7Qv䱺�ٷ�(�c�S�Jx�)�C�چ<�)1���8�|�ȽJ���r�<�'L6 Mb�N�/��\��	ߺ/JDD���İ��?���;�f�d$���|�I�;�
g��폳��BɡG�i��<fL """�oP�m~Q���(  M����-_@S�� �H��������rM���
�jhѐ�q�� |�u\�W��u\��	�w���fG!"���bL����OJy����a��9�	)��_�bE�ɧ�=����i�&�(�������ƍa����5�AӦM�����D4��y������׌��R~���,�N���],�H��m�w�x�����X�[��M_�H�/��A�F��Ն��į�|�	@UHDD�]����V��'�r�܃M[0��{7\}# I�u�j��F���wܶՀ4DDDD�'��w�PL��>�H|[WC�q�f"2�����=�Fasd�׏���A	�����÷u��܉G��m�Qw��Q��2����?��.k�,~*��9�5(=���K�89�5q�9�{2�lDF��wUU��ND�a
��� `砊`p�}CD�M��a�/~��Zý�������F�/�ޡ��D�|nQJٲU����k*��C���Oqw�r���v-���JDDc��֒R]��P�; t=~����쇲#��KEс��Ä�������D��v�߼fT�٬���>�0��$"sļ}�m�jLl��tҢa��~�����(D���H�ͫ�F��6��@��������(#�u,�)���`�q�9�/��z�s������Ӕ�mǎp�\X�~=,$�t�1f̘��y��ۉh�*=�p��+R^ǻ����=�8u��u��Ύ�x����I)[��[���>��bA����h�kڒ�����RD�zHDDcEl�#t�l���	�'p�z�u_�p�,�4\}#����D��7��7��罕�!"""�)ܷ���f�H��״�S�@α����H��o�'�6zo�ES��7}��)�a-(3;e5��j���?�NӀ@�W��T4����PZ,�P[�.k厫�d�}�1�fCn}#[6�����w�3����!�ʎ<9�q��t�-ͩ�F���;�{"m�%+���+V���3`�Z�F͎EDD)���Buu5 @UU�B!��X�)���˩������e���w��~�Oǝ_2{�jm�[�s���s.^MQRΖ��P�ߍ�7�V����S�q�6o3(ٷ9N9�uB5�����JDDc�I��	��~�-�~�cB�5�ݽ�-��d}�{(�=G������W"""2L�݉`��f��FB�m�ES�d��\@D�"%8����Ds�.�����N�>,�B��Q�b��>��i@��+H��JǙ����0��|�uYk�+�"o�^C���벾s�"�]q$��[�K+�N>}�/����2�k%-E�K�뒍�h---�����իq�G@�e��x�E""�3I���>���y``���D����O��u3�[���������Ϡ���D/Ip�;���%n]�O�C��z��7CS�z�.���2��bA�e?E�/�10ٿ�e�����^]��|"��$���^�:|��H��7i����_
��7�����(;)~7-_{7өA/;�`,f'��E�F���14e�M��bQ�}-6���آi�͟A	�̎"LӀ@�(�A�����|����#IB�ɧǭ�k�.��!����W���� �V�Y`DD4�L�8��;O�b1No'����^�z�c�yg;��q�Yq���
��v��e#5@�#��UΝ����H�m�S�Bn��.������[JDD42�w`�wQ�������Q��C����ۉ���Z,��A|M#�OQo/BNޑMDF�lY-6;HҔH��/�ޒ��ڄ����I�T��CSbfG!"" =����xn}#J����K=��	qk��/�3��v�؁p8���~�$����ؐ�������]oLLCD�~ý��U:�����.�N�[��u��^���>��]S܍���v����d@""��7���)�?��p��z�W�a@"""" ���H��)wmB��6;e�Pw�^��F����cQ��z�vn7;F�Ԉ���f� "" �+^�Kwǩ�>6�c no��G�隍�h�Hmmm�������)�DDc����w?�G"D"���g�;�N]���q��qύ�z�?�5@ף�
�=��1r�ĊT��nL "�	7�Hj�	#�����������ON�#"""CD��t�C�Z��u�N��jv݄�6B�rd"ҙ�"ؾ@f����#��76�uZ4�ޗ��{��~[y�e�(;�������4��ݝ�({utt 
���_��ilr'"c�������z���&�!"2���g�3q�v4rjjw�l)(D��s�۳�Yh��!�Qד��)�-���}�_F`�&%.���������uFMq���z���M�_��Y����4UE��k�c�J��m6;e�`�z@˜fMQ��`v"�0!gԐ���
��c3$�(�����7�K6*�������3 ��9OS���������*�����ݍ���
���;Q�~dY�̙3w���1���S��E�e����I����r�<X��ѻ4~�<%g�Mq�>�l��֋�ɘ;�    IDAT*:�M�,DD��jpF����sP|�!�um���_��!"�ۡD�f��]�k4��>b�>Dz̎����J`��D�!�X�&�c�N��o5;Q�6o���O��>�����1�̸�x�}��NC��C__���o#�f�����0y�d����������\��.�~'�1ǩg������Ύ{��'�ܞy�?�m�Lq�srPw�5�u��_A`�F]�%#���2Ž��$��7mF���u�@DDD���"ԓ���55�p��cQ�uo5;�a2�w#��
�l����Φ��Ń�h��Y�T���&MAѬ����ț<5�9���(-�m��χ��{�$�b��������� S���k��5C�7%j��u�u(�}�퍂�g�=��댡�z�>�:���;柍�q5bE���$!�wh��S�K=���k���ۉ�����Vh���1��M�����ߍ��ev�D��99��R�Ţ��0;�a�Haw��1���^�k/"6"��p�� �h_<�02QZ��~8�N|�������j���.""��̙3!�{q,C(29����~Ѿ�;�V�_�qg��Xlp �o�fd�����C���}��w97u�\-\�z�U6o�%Q��op��S���L�&ش.�q&"""��]-fG0��"��2;�q���~���]�f� �1.�逦d����>>W�M��Z�R�c�?�	*���X�OC�E��F�6---�F�X�lTU��j5;���Ѐ����?@�4�Z,�ޗ�=V~�	��;/�C�����` ]��7Ž��s����q�-)_��H/)5�C��q�m�ezLq/9�W|z{�]7qz;"��{#��fG �1LSD2�F����lD���+�_s)~7����DDYo����|�v������18Q�D"�����t⣏>�,˰X,f�""�o����{�w���f;"�]z�_�;	�f���(~�O+�u=�)S���\�^|�p]�[����딮MD�����������Ku�{���k�۶���+I_����hO���oB���-�m?�(9��H j,�����D4F�?����i��0;Q������>��jm60Q�uvv����wށ���j���n�DD��}��6�m�σ����ND���m��$��}_}!�>����z�~�T��W�~.r�ŧ���+>蘈�H)7�'�����9G%5����rz;&:�-����>�C��=ϕ�����������@D4Y�K0�������iw>���s̎�2��}��40	�94MÖ-[�F�ꫯ �V�ɩ�� 0nܸ�?{<��� �Y�0�7�������{G霣R�:8�ٝ+�|_�6�i��.������u�o�+�!�DDFJ���oO����+��	�l��_˄눈�����P�>�c�M�+�&��h��/{�?b>�DD�ɦ�5����̎AD�8I�^�=����A��i(?����b�Z�jν���&����PC�ϋy�p��<������������X�v-dY�,��U*%�n�c����s$A08�k"��L��]��B�O�����3|���]r�%�f�K�k�K��x�����KiHD�����^}�y���t�{�p���=�ih��fL��!��]S�ݫ�J�����Qt���	�v�M�E�����(��Ȣ�0��A����FP#����B�E!Ym#�LD�����i�i�֒*��%$o��r���'NƄ_�	W߀��O�� �>��v�k���q���!68��7_C��y{<����F"�� 2[kk+*++��o`���(,,D$��e�DD��~�����>[�x<&�!�L�3���?�q��Ih���Qw�u�]�Zo��&M���P����a���R��z�ET�q��s��"�n��x5�]
[yE�5���7��k����^�:|��
�M���vMq/���P]��7����@�5\u�p�P�v���,\GDDD�(%�5;BZ�� 45I�V�D�8%�e�j;�>X��NBDc��@�eW���
6���`+��k;KQ1j.���Ά��ɦ�͎���'�g�S#6��lyO4����[�b����o��SN9V��h��hDDYg	p8��z�P8Ԑ�t`+�s��%� �\���O�d�B����ڱco��Y�Ԉ��ŋ�@C)?� ���R��r�<t�w���:�����'����[�k���A�}�4w�?��➈�ÏF����F�]7�ꭎ��؇b�q�SK��݊j8dP"""s���k�TC�S����������Ƙ�{]	@�¿D4v�l��5���P��v�m-����'�j�>�q��"д��D���� ������_c�ƍ�e���XDDY���3f�����(���ޑ��lnJ��ܒ_�ks�
"�m�n���[���=ز��k�@�u?� bn��;wMqO�����.��^�&|��K5*6ft�U	��F�%!{�kp�z�U�7}-\�p���$�|ޕILoo݁�W_�K'�/��?e�AI�c-)��Blʖʭn��(�dc���s"�f�s�ƦM"��ϕj(�~g"�b�h��Ո;M�?�.y��A>�����p���G�c�����x�W��za�Z!%�]&�N�ep�ߺ���v����2�
a�����S���b�!�����������4������;y'�x޸�.Lnz��7פ�����oʛ:ݠ$�˛����
�*�vӵ����$��Hd�{ّ�&7����=� "�.��N>���W����
IprE��ݠ4D�'1�oNѨ�_L��������F�k,"}��R��ߙ�R��ϕ��;�����k����a�_~��6�6oC[��p�]�,����h���-9-�FEQ��ԄP(��K�B�4�tܕ����7c������"��F"җ�X�����N�NU�6���ï }�^�������i�@�u=�`B�|S"S��|�^�P8����}��p]:E��B�����1�i�[S���}_�&��aP��Ǫ���7^E`��O�[�����~�m@ӆ�e�_u�p�P��-["\�n��m��?H����f���������J��a<���PM�՗��6D��WU3q�w�2;ƷLh6;�>��i���@��Ĩ���cCd��LD)��,|�`�;�A��t=v?� %�����P~�q���6����
��:�wP�u��u���Q{ѷ�o��D������� ��>��r�V+b�@Dd���*L�8q�ϊ����S"2���{�#�^�����3�G����76�n��+�O����� :������;�C��������z�>4��Bu�s��ۆ��~܂`����~�?�k�-ز]�@�0�ǆ��Ž�?�$��w�99Bu��[JD4����MC�]7c��*+�wT�tz�>;�X�9�p����t�{먟� �/?C�`M���j8��'2$S"�&O��{���L�n��JDDDd��lDʾ�~"JQ>Wf��"J��}���,���(�h>|�kiʏ9%�� ���J I�K*~B-��k9\��-��[o�3�` �?<	PU8�2�mԉ2ASS����r�J�?���PU�����(���v̚5�[�������h�ӏ0��Gh..A��ǡ��`�o���H��zj��P���x}˖@��w�C�=�@�FP��� YF�Ϣ�;Ӛ���z�AԜ�%�	�H����t�9��������?��y%�k?�K����PC!�v{�5E��n[�_��50����\L��-(;��:-�S���I�w ��^C`�F��&��&�TV���)�������朋Q���Bm-�}��:3|�Z,*4�E�X0��F�	?F�S���v�4LE�rrao����ND��A��^���
��X#���Z\bv��h���	ID4�I2�,k̑�?�!�,�ć�c^6��D��l|���ߙ�2R��F�O�照͎�MQ�~�Mh��&���.�aӦM�o���d�\z����A$�oWj""J�$I��w���o�r�"J��� z_|�/>gv��h:��M������L�I��`������#�u$�eG� �X��s��u�p��H���F�aGՕ��Z�>����V"��m� ?IBNU5�g�A���!��Qx��OWCG��l�C��5���g�uip�����b��Ħ�KV�k4���PCA�����t�w[��~KV�������c�k�<El@*c��0��x��4
�]~-꒸y�,j(������[y��%Y,Д���C/�d1;�1�Ř����$g��LD����{�%g��""";���I���o�G?�l6"&owOD�I�O������?��a��~g�w����Ǟ��cO��@�X Y��,y`�;�~�iR�f�{�E�w ȩ��������ƀT�+�)y��*�]v*N�1r��͎c�vO0l<��Wؼ!��T���]�}���������fGH�ޥ� ��I�Dz��v�}�}�Ԝs��q�h���wb��بJD���f�l���(E�����M�DDD4�������b͚5زe$I�՚��ۈ��p80y���?k���cb""""c)�At=v��rNN��� �~�ؘ޾�k�K��:͎a�����lv2P��Y��啨9���nn�Ho�.��������[[~O:�ZtlMP���"�B�����1O�X0�WB�N6;
�2��nv���s�ق���.9'��7�,���(5�-��7�|�#푦iؼy3E��e���za�X`I��������<̚5�[���n��jR"""���z�S��|�?�8��M����{͎a���n�
���3���[[E��Q�"Բ]�u�kp�z��7�3�C�Zw�g�i��^����@�Q����w��q����?��ݸA�  �i��N��$S��3eg6�rj7��H��&�qR[NM6;��I%ٙ����đ��-ˉ]N$9�aY�Y'E�A A������s�0���O�W��Ӎ�/�G����{�Z�ӧ��~���鏯�L �mz��3#�G Pc�H��+-�� ��ِ�+�s  �gqqQ����f����'��+۶eFУ@M�,K��s���pi[&�Q�Pp*  *�M%u�K^(��u��{e�s��=�%-z���=��?�(����G�::��b�^����NYwy������|��ws����Iͭ޾,}`�N?��=FY���[��S��K���'�1 T+�X�aZ2�H�c �1����3Tp}�Hs�ER���  P����555���Q=��Ӓ�P(�T P��o߮�������*�Jɯ`_ @��<��Z:Q���y�	��z�b����bQ���w���p^>����]'�QP&�e��Cz����{jUn�����Ծ74��/��n$I/���g���}�˩��3-��b�c���与��^� ۼ%� T;��e�ڤ� \?��E2��gh�0�g� p�CfS��WG�X[�#  �20,K�H�-�p��q��y���ڿ�� r���i�&������}_����� ����:���w��Թ�N~���~?�>������=���}���g�9r0�IPF��5�[�u��G����ت�VEʂ���-��oe���̔���g*�Z|9������iez�U�,��ȯ��
cg����\���Gu�	 g3�ZeX��B���
z ��0e77�Av��c� \�P�qNSi�"�"�� �z�H$�.rwG���z�'466&�4e�vУ@M����-�ܲb��ܜ<�h"  ��z�U������3�����#e��r�x����z�Us�����v�c��_(HW�8�[\,�4i��Й���U��H������|���ܾ�I��g�W�'�r���S:�������zUJajB�?�1e�=J��N_��G��3*jq�x�# �"�!��Ǩw ת����\��F�Wډ.� @����=�NkppP��������(˲d��s�2 ��XLw�}�����d2���N @�ƿ��F��O�v����~�e��J;�W�����h��5���3�MГ���:ʟ-��kAqfJNr!�1��w�:���Vqvf�n�bϲ������/k�{�����$t��Y��^_����\БO�/�x�A�rMR{_Ӂ_�Ye�9�(�>��U�Xg�z��Ӡ�3�Zx�Š� PeBm��"�PTV�qV`��Bmk��B٭��Xmv�S��g
�6�ch  ]=F���������o��}�B��& �l��Ν;�KۊŢR�T�S PN?����~O�j������u��t�n�J�~���o�M���g~N����5���=J��<��_w��^�������٧��kP�|�щ������xUo���x�E|�75���Ǫ���|U��}u�/��y����;����9*�[�j���D�>�1&Ƃ�r<O'�쏮誙�4��w�<������\���u���a����#�Yd�5��	ٱ֠�(;;�)3z ��0n�z��3��B-k�  �I�w�u�z��O�8�T*���!���Ң8�p�� �a�v�ءD"Q����fgg����  �������G�=��uߖ37�w~�S:��ϯ�d�i�_�Eo���5���A�r�f�~Bo���4������|��83}��y��F��T`���^���;�s:��_��w����y�&�����{5����[�^��/ױ��-�ĿW~�t&�.s�=�}٣�?�Oʝ:�8�S����߯�}A�Sz�������_��K��$7|BG�ï�w�
N�U�y��KYv� j�aZ�2q��/� ԸpG�#�]��}%���l�}e�z���I  P����;!��#w��t���E��G?ұc�$I�Pc�� �ԭ�ު����fffV  �̑����׉�}V�ё��x7����K����4�ç�0auɏ�������/j���j|l�y���s:�+?����u�h���(�L��oJ���E��
:���̑���r�c�u�?|J��\У��u4�����^y�,�a����@�������G����+~�]��?��;7�V��a�������Pz�[����a(q�N�?���ح��[e��W|�PPn��R�����/h��g��r��������g��k�˒�t���w������T2�	���������9�1���f�����C_Pj�A�s���ܩ���3A����C�p�c ��]L*u�E�N��-k߼+�1 �8�s�<��N!�Q��Eղ�}D� �[���r�·�����gdF��X5�~��u��sA� U��P��_�Y�Y#�R)��� �Z]mmmھ}���>��O���W��Xl�� ��_�/��/=�y6mڤm۶�ض���l��C�E=�i}Νz @-2M��s�:�R���m�Y���`Z�u�8tB��4���k���-4p���z�����e��j�v�"k{+�z��)?1���J��f���
cg*;C�
�]����}u�쿓��$�NQ�/��S�_�y�P��_x�Z���g����*�v]��\�uU�����q�?��f�y�Ĺ���2�b�[[e�[��sr�夒��_+�,��U�]�� �������x�"V<���u�r9�N�wݠG*+�)&�NW$�=On:���������*.L=FYķ�/��#�1 ԁ���rcA�QM}�*ҽ1�1 �gaJ��W��,B��ռᮠ� V�; \��~�vS]G����ڰa���>��O���E���q8�/�ʨ��}�ڵڱc��(m�f�ZXXp��"p ��-u��m�ݥ��M-�+��R���e%Ze�b�?wqQnr���evH���2�a�O��[l��eF"2#ѠǸbN:U�fخ�]o1��bV5ީ������f��p�)-��(�Jx�Yy�{   �Y�UŅI��2�Dq;�U�ZWx    IDAT�ڨ�Ԑ|��V�3CQ�;oz u�n���.'S?���$��k�=  ���������=�HHR�D�N�R<���7���گ��"��|ߗ[� ��ttt���^�
%��y�s  ��w�*�L�83�(5�+��L�8�$8���z��y���:yN�\8_:  �*�c�
w�=��2LE��=�:b�!5��%�1V]S߭2L+�1 ԑ���V� � �f��h<�1  @�����ό�?k��D"�H$�T���ѣJ&�����c�=&��d۶,��4�D"��;w�<����innN�__�   (w  �2h�E�z�U!BP�~���A��jB�n���=�:c5�(�uc�c�3U��� hX��{��#G�(����ɓz��'%I�m��<��555i���
�B+�OOO�;k�    ��3)   e`X!5�p�T�mZM-���� ꒡؆;e�vЃ\7���ۃ@�j�EV4���PӍ���  ׮�#�B��C��q�۷O/���$)
�ݙy �\�pX�w�V4]�}ffF��4   �ZD�  P&��5�to
z��b��bw�`�) eb���tc����Sf�)�I �)ôԼq��
z��]�E�DW�c  �*P�{6�աC��y���y8p@�R�I��^ٶ�]�v)_y6؅�
���   P�(�   ʨ���5����.Y��GP��m������,ڳU����� P��h\�n��3�Z�(�Y�  �Y�#w�}�)rO&�:v�|���?���aID� �eYڵk����VlO���f�M   ���  ��a�y�NY�֠'�jѾ�� *��w��}A�q�7*��`@e��׫i���ǸjVs�bv��  �뽅��71T�����N�<)�u��o~S###�����4u�=����c����E�R���   P��   �w�e�y�ne��Xn�6��m�Y��A����b7�.�-��0�4W$�ޫ��ۂ@��to���?�(WĊ�(�i��
z 8ϫ��z����WD����igv>�1Pa�-���!=׳Q����!�HH���|������E�Q�������?�q�[�N�PH�bQ��=" \3�0�c�uww�؞��5?�����ަV�����WD�ܽ���2�A� ��   `�o�_���夫�zÐ�}�)�ucУ hD���ƝZ<�_�������H�5��� Ttݻd�eGI�� ʎw�y�NOA�>����/-k�x/ژ�ۺN�ahwf.�QPa��?~\�pX�����7��O~����&rP����w߭���g�-������ ��ͦV}�u�|ΌSUN��*�ޛ�	z @�3�   �QvH͛w+Զ.�Q.Ȱl�6�$n(Ðb��)�v���{R�0E{oQS�vU�| G�{�b�ڕ���}�o�M��*�k�w[�۫�/�_Z������GA �[H�}C�\��-�H(�8���<O����٬����iffF�a(
= \���׭[�z�뺚���� eG�^ݞJ���Π�  �8w  �
2LK�w(v�2��y(f�Z����Z{.e (7�Ptݻ�i��zB3V��݊�lz �$��{��=��Z��SM}�*��N����2���G����[H��u�:tH�TJ�LF�<�d����, 5�4M�رCk׮]��u]MOO��&�(��k�; �z�*  @ �}�o�#+�� ����-Jly��ps�� �9�D�Zn~@����|a�d�}�]�� �"͊oݳt�M�/���J���"�� .���v�7���q�<�t:�d2�GyD�L���;�;�jg�������v��433C����k�; �z�  Ċ�(�w+v�m2�p���nY���߫�w��&��e��jްC�7��W����%n�O��d_ W�0ME{oQ���r ��(v㝊o�OV4Q���+A�^{��[=G���СCZ\\���y��r9"w U�4M�s�=����kjjJ�Y�l (���D� �V�L   �2�Q-�~`)tE�~�v�K���V|�.�VmPB�n%ny��7���/���n�S����� j�M(~ӽ�o}�B�=R�_�3CMj�U-�ޯpG_�+�����."��Vϑ{�P�������499�/��J��2C�p��@ձ,K;w�Ԛ5kλljj����q{m#r \;�    �4�Q�~&T�UqaJ�W�Ia3ܤpG�B}����,C���Z���̩8sJ��1���:�n�n�U��O6�f7��޴S^.���)gO�+�V��S�֞�ǖ-k��T=��ڷ�K���\�à��SHKC�A�F��%i)r��|>�h׭P(�������555��~����'>�D"�p8�B� �g� x�pX�v�R[���NLOO�r;��#n�O%��zoz&�I  ���  ���Bm�j['�-�I��IO������HW���a�d��d'�Jt�jj%>P?Cv�Cv�C����df夦夦���p�(ôd5��Nt-���%���f4���[��{��삜���J7� �-^ٍ��h|i?��%;�)��)E ����~�7�z��s��<��o�]333�򗿬O|�jkk#rP�Ѩv��]��mjjJ��:O ���ח�k��҃"w ���j  @�2��Bmkj[�&I�}y���|Z�[��:��ʗdڶd�d����qv8���2�T(ѥP�ki���+����R� �sK�a�2L[����G� *ɐk�kS��&I������r�y�+�s�$�Z�WZaY�f�^@P�����r��K��Ƚ��s��f��~m߾]���z����\���
��*���@n XM�XL�w�Vs�ʳ�������v eG�^��nYZɝ� p9�   ��0dF�eF�/] hT�!3�$3��$ P�L;"�#�� ʀ��~����J�D�#���n�$}�k_ӯ�ʯ���G�P��@ŵ��j׮]�D"+������i�v eG�^߈� W�s�       ��@�^��#�W�ۃxO!��O�s�ҶD"q^�Y����okqqQ�LF_��W5::*I
�B�,MPk֬�}��G� 0����5z��3�1  U��        �<���A����9r���ڿ�2��r��y�I�lۖmsrn ���߯�;w����<��@E�7"w ���       ��F��x����"�h4�T��P(h���J�R*�z��Gu��aI�eY
�BO�^mݺUw�q��s�R�u555E�����; �b�       @�"no\D��=��>81�"r���u�;��haaA���;���^x�I�i�
���� p�,��]wݥ�[��w��8�����yL���76"w ���       ��D�"�ƶ������u]<xP����}_/����qy�'�0
���\�h4���O�ׯ?�B�@��"��!� �G�        jq;��7�z��=�ӡC�499)Iڷo���o(���0��a�&/��6���ڳg����λ,��kvvV��#- �E܎�� ��3        ����\D�#��G���ɓ����!}�+_Q*��$�B!Y�� jкu�t���_p?��f��Tq;.�� ���        ��v\�{c���]�FFF400 ��511�/}�K�$ٶ�P(�� j�az׻ޥ;v\���d2���� &�h��q)D�  ��        ��v\�{c���}bbB��8J����W��'NH�L�T8�A$�"��v�ڥ-[�\��9e2�
O���J<ݲF�ǻ�  w        P���q���۞BJ�[�������~�m��y
=����~ ��e���L������ڪx@����]���fff����@�!n��x:�M� �g7        @U#n��"rol��`G��lV���S:����z����o}K�|^�
�d�v�S�}}}�������t�e��hrrR�B!�� 4�v\"w h\�        �j��Z-G�?��7�z�����~�m���H���/}I����$˲
�d�˶m�y睺��;eY�y��r9MOO�� ��h��q=���1�       ��D܎��Kz��ȽQ�{��y��9��'O��}�������Ç%I�i*�4yIh4---ڳg����.xy:���ܜ|�GY ʏ���� �f        ��C܎�B���(��������}���Ȉ>,�qT(��o[O>�diU�P($۶�@�lذA{��Q<?�2��577�T*�d q;V�; 4w        PU�۱ڈ��N��#wI����[o��L&#Iڻw�y����e)� .�i���{�}�����u]MOO+��0�FD܎r r��A�        �q;ʅȽ�5B���o�>MLLH�N�<�������А$�0��aY�� ��4Muwwk�ڵ�<��kjjJ��Tx2 ����D� ���        T�v��{ck����<�رc�<O�tZ_������O�>o۶
�X��˿�;x%�JivvV��#, �A܎J r��G�        G܎J!rol��K����8�|>/���ꫯ�����555%ii��p8,���b�V-�/��Ba���jzzZ�t:�� 4(�vT�; �7;�  �-�R����      �.c���z��E܎J[��%��\�à�p2�ؠ�Y�����qIR.�r�U�L&�o�>mٲE����C=�|�ڵk�$)
�u]9�� ��m�+Vl�O<Qz?��i~~�U�Tq;��t�[��`z:�I  ��� (�
ˌ4=     �u�E[��f�#(DQ"�B��C����W6l�$=��S:v�~��^�x\�eɲ,�Ey��� .�4Mٶ-�'��8z����k�)��J���絸�� q;��t�[���!r���9�        @ ������Ǳ��GA p2��ؠ\�-m���F�NUgΜѾ}���d$I�������cǎ��
�
�J�,��b�������Q}�_ԫ��*���y������Tq;��3�n�0�� �U�
� �@ZI�>y �1VX�ެl�C      ���Q-Xɽ�=�d;�ﭻ��Wr��l6���zK�������f��c��;��?�AE�Q���p8,�qV�� �c��B�P�}�u���P���|���ܜT,�@�"nG5y&�-����^�@�<7��{���c��?�yM=      *��ՆȽ���,J������%�ImݺU�HD���������X۶m���R�eY*���@e�!۶e�fi��訞x�	MM-��溮���u�̙������Q����~�       ��!nG�"rol��K�����z�-mٲE���J�����������#��ZZZd���,K��Ӝ�X,��_ԏ���A'��}��G܎jF� ���tW�� и�m���{oz     ���w��6�B�cT=�vԂcѸ�<W�E��F��9jʦ4��^Z19��<9��t���<MMM)�ͪ��M�eivvV���S(Roo�Ði��,K�ﳚ;Pf�i*
����cǎ��G����%-������u�o�7q����<�@}!nG-�4˔���z �5bw        Pv����'�������pm%wI�����6mڤ5k�(��멧�ҡC��s?�s���a
�B�؟�X]�aȶ���5��N���SO���åm�dRǎS6K� ��%�� ���        �q;j�{ck�ȽX,��ѣ���Ԗ-[�D4::��zH{��ѻ��nY�%�4W�jO�\?۶W������|�M=��s���$�u522�ӧO�{ 0��ED� P��       @��mj%nGMZ�ܛ���|���1r����9��曺�����+�u��/h�޽z��߯�n�M�J���8r]7ੁ�dY�l{e�122�������(m�������U(*=" ��&��Q��It+�ڝ��e �%�        �lN�c��Y���PTw=Ѩ�����Ԕ�l٢��f�R)}����믿���Z�~����<�8�<�xr�6��)۶e���R)=��s:p�@i��|>�'Nhff&�Q�d$#nGM�����         �4j�.-�o���������'˲t��i=��ú���|@���2C�PH����p���q�ۿ��^~�e9�#I�}_ccc�	    �;          \D#G��kddD���ڰa�zzz�����߯���ٳG�w�i����E�!۶e���Գ�>�T*Uڶ���'N(��TzL    �*�          p	�:�2ǎ���%�P(h``@���ڴi���r���}�Y�ݻW�Ї�e�I*����q����@0.��8qB�=�����K�r�����4==]�1   �*�         �e���J��KR2�Ծ}���եM�6)�hvvV���7�~�z=�����4M��aBw4����gΜ�s�=�����6�u5::���Q�z     g!p         �+@�dzzZsss�������e��N�>�o~����Ӄ>��7J"tG�X�>33��^G�Y��?99���!
�J�
    U��          ����u5<<���qmܸQ]]]����Q=��#ڸq�|�A���IZ����jը�iʲ������y��G?��o��"l��������t�GE �z   �&�         �U r��\.�#G�(���oTGG�$ihhHCCCڸq��������W�Rl��|ߗ�r]7��kf��l�>/`�����/��}���8�#�JixxX���A"p   �	�;          \%"����:�D"���~uvvJZ
����A[�n՞={J��a�m[�m�u]9�����,K�e��OLL襗^ґ#GV�؞�fu��IMOOWzTT��   �&�          p��ϗJ�t��a���hÆjmm���:z���=���~�ڵK��rK)^��Wt?;��a���s],l��r:u�&&&��n`�i=   P��         ��r��_�n"r?K2�������֦o�Q---��S�N�ԩS���Խ�ޫ;�u[�=ϓ��</�O�i��,K�9����:v�^y��<yr�e�lV�N����a;d_�    �G�          ��bF+�_���������ѡ��>���J�fff��O�?����N�޽��53M���;*�R��
<xP���fffV\��dt��)MOO��&#�	   ��D�          �i��(�_���fgg����۫5k��0e�Y����z��t�wh������,}�rh��~)v��b��KKj���kڷo������2��FFF4==]�QQ#,�R�)=   P��         `�r原п��L�~�tZ�������#˲�8��|�M�ݻW7�p���.m۶��u4C�m˶m��+���y^��jݥVk�}_���ڻw��=�bUv��5;;�ӧOkaa��#���B!52A�   �$w          X%����O�q"�K��r:q℆����ӣ��>E"����'O��ɓ�����m۶�{�QOOO�c����q��(��n�y���i�߿_o������W\溮���t��ie��J���ջ�~   ��          ��v���q]WgΜ��������~�z577KZ�Z�ݻW{��պu�t��wk���
�å�_��}ߗ�yr]w�Jۀt����}k�޽z�w�;`"�˕~N]׭�بq�mk��z   �&�         �*#r�:��ibbBjiiQOO����K_���1=��z�g�}�v�q�Z�~})V6��+\.j����	<xP���W:�^q��������ؘfgg�Y�U	���}_}^1�Q   ��D�          e����3~B�J�~U��LTNq    IDAT��ɤ��٩�����I�
�BiU�D"�m۶i۶m���+}������r]��U�Q����i^4j_XX�ѣG���ok||���������466��)�Y$�]`�v   �Z�         @��W��f%�k⺮&''599���f�]�Vk֬�m/�̝J��ꫯ��W_UKK�n�����+yKK+�/��"w�[��.�]��⢎9����ktt������������������u1C�pX]3A�   �,w          (��ŬD�~]2��N�8���!uuu���G����U���d)vooo׭�ުm۶���g��B���"xGm8;h��*�4;;�w�yGǎөS�.�g2��A�B��c��D�Q��;�G   j�;          ���bV��q}o�MD����R����ե��.����b繹9���Kz饗��֦M�6i�ƍڼy�"�H�ÐeY����������]%�4h�}_���бc�466v��-..jjjJSSS�f���0555�u]�*d����   �w        �U��٢�wo�a�i���zm�	M�$���I�:��X�}�
�9sFgΜQ(Rgg�֬Y�����u���w�^�ݻW�e�n��͛u�M7���{���KZ��;�{��!�0�(h��l6���a�8qB�������5==�d����|"��L�T���B��V��6�ݻ�Ju�w��K{�j|r>�Q  �(w        �U�ݑP[������z[������ZZb��u�Y�JDX,j||\���D"���Rww��D�:��jhhHCCCz��g��Ң�n�I�7o�ƍW��l9�^v���D����}���)���ࠆ��499y��A6����fff�J��^���P,�$�IO<���ўPk�������lUk|���3jk�� ��;        �j�5:�����g3�j�Y��;�ﭻ�Ƚ���N�>�ӧO+���]jkk�m��%�d2YZ��0uww�nP�������v�m_(�>7x_~�O��_ne�e˫��<yR���:}��\׽�u}�W2�,E틋���) ���d���\N�:��5�_��Q�U�����3�tj&�Q  �,w        ��VO�;q;P�:��Xɽ�
��&&&411!�0�H$��ѡ�����[Z
�&''599�7�xC������W��������{������vv�~�[=:wE�巫�N�522���Q�9sFgΜ�h�.-}���577���9����4�kb۶���$I�-L<�USG�;q; ���        �C=D���@Y�,fe���?�W��
��dR���
��jkk+��
�V\?�Nk``@��p8���^�]�Vk֬)�-��u���b����m�s8;Z?w۵���/|066���Qe��K~��ZXX��ܜ���/{}����$�Pп��<�UU�;q; ��        �K-G���@E�(fU;�ﭻ�Ƚ�
�Bi�vI��bJ$jmmU"�P,;�����.m3C���њ5kJ����]���4�X�~����}߿��}������]�|>���)MNN�����I����~��J�RZXX����R�TՄ���D"Q��67!��Q���p�N� �U�         �T��;q;PQ�:�
��{�٬�٬&&&$I�e)�H���E���jii�i�+>��}���hffF�.m�D"���T[[�Z[[��ޮ������V}��rD�-��ivvVsss+����U&����)
J&�ZXXP:�&hG�kjjR8^zg1��-�u�#w��u��ҩ٠G ��        �[-E����ہ
�Q�J������b��5&�u5??������i�������bjnnVss�c�|>�3g��̙3��x<���6������U�x\MMMjjjRss�b�����
���9^��8�f�J&��d2J�R��<�N+�L*�L^����+��)��(�ɔn�q�2}&��D"jnn���3������ 5��"�Rܞ$n �&w        �J��Ƚ��=	Аv�rǎ�u7������R�`y�W
���FK���q��V\O��J����}Z�U���#�Hi%�h4*I
�B���#����쟡|>/��J?[�o�|~ſ��^���)��g�y�wݷ%+�H���m.�i�!�@�N� ��         �R͑;q;Pv9��Xɽ�,��333�m�i*�^��B��_��J�RJ�R�U
�r9-..����],�XU���Z��K�7�ʫ�ȝ� P/�        *�#w�v����{��<O�lV�l���۶]��#��"��lۖm�
�B��C�P�'_�u]
����y�E���UY��MMMjnn.��9�~sjH��8�@Ta�����3�t�� P��   \R19%U��MC��5AO �$7;/��z���2,� ��TS����xR��|�s X�����8J��J�ӗ��a��}9�7MS�e��ILg�K�-o_�o�4%-���O���}_��n�u]��+�q�8�y�Xb�b�����J�<���M���whXU�<2�L��� ��W7   \���^yn��F�0���Ѡ�  IR��ѥ��P��d�Z�  \H5D���@U�Q�J�D���X|�W�XT�X}���²,�����������'��x�4 h U��?<�,q; ���A         а�E����ɯ�}�5aG1��;.�uK����h�S@�[^����mE��y��8��N����:=����w��� ���        ��-���'�+T�n]�$nj�.gQ�9+���qIb%w (�p8�x<.�\�n��z���,f�@��58��q��[�1�� u��         `���u��O�g�g���(f卟��D� P6�HD�XlŊ�˼bQ��b �����-�w  ���          j��bV&+����,K�HD�h���K�I'��ٓ���
O   4&w          ��� ��0�B!ٶ�p8,۾x:㺮�̌�٩
N   ��          j��bV��	�󺕑�i�r'�� �z�!�0d��lۖeY2MS�a\�cCs���3����   ���         ���p�_�=�< �>3����u_1�(   @�"p         �����9~B�|V� �z��)�N�éI�(f�   hx�          P�v��; \5��d�uSjN�ͩ�w�	   �O�         @#r�K�}_���.�Ԛ[ԶBZ��j���G   p�          P�v�J��I;�( P�=W1�U���/*��A�   �
�         @�����=     �u1�                  ��                P%�                U��                P�                U�z    \9'3��}/���%IVS��HLf8�h             p��  �g��8����
��T\�\�79)gaBNv^^.-7����\�����2�1����D�B-k�X��o�:�Z�*�f�"=7�E���������O/�#S�*&'T\����R15-y��̜|ב�K�+��e������gF�b��b���ZK�j�Q��_���
w�+��/+�����E��*Ώ�8?����ޝ�GUl�ϙ}2�d��daI!,����"V\����X���W�o��V�V[����j��.��]+
D;$d#!���d2�9�Z�$d�5��r�<s�����<��Ύ:�{�_~tArX!ٻ���  {<�BQQc�B�.
����LIPE&BmJ��AT���$"""""""""""��Ƃ;�؛*`=][�)��O�V_[C)\�V������������ uT*���I�m�D��M�>}&��(�d#"�G[�Շ�s�(�e�7U��XG[ K�:�,��\��� �:#4��Kʆ.e
��Y�&O�6~�jX����Kv;�=��5��>V6���P��X�C���]<�0��I���kb4q�|�$"""""""""""�!c�����h�9Z�`)/���tW���@�Re��e8Z��h�N�<oH����Чπ>#�B���SP"
U��
t�����>k�!�,m��Շ����"XO�w��PA����9?a��K��OI�(�H�nX���Zu��{=s����h z9�k�h�E��]�	J5��S���GXz>��ЧN��T�',܉���F��Q����0��c��T��H���RGK���wwNmbYa�r1�9K�4��9%Yr���0�Jv�rj7�N}g{��c���v�NO>������2g#<g)�S.BX�l
��&��q[;�U�]��FW�a=} ����X�"���]����m�R�����Y�������לDDDDDDDDDDDDX�;�IN��?BG�?a>��͕�����FO�	�Ԟ@��� A�>m:"�_����0��;QNs:�������|�}�,����u�3��?���G���P�#���܋��ڤlG$� "���*���ކ��G�Vd�߱�Fv9`)�K�^Կ�S
�EASW����wL""""""""""""�#܉�����Ղ�Co����<�${��ϩ�����0h�Zh4�T*h����i4 ��n����n���BOO����}8���(��v-�{�GPc���3�"r��5a�{>"
��#h/�:����E>)j�}|�h4�j�P*���t�:�\.88�Ntww����k���Nt�E� h&�4{L�7 ,c ^;7&WW�'>F��7�Q�&����KE�F��z�t:��z��z��j(�J��j �V����$��1�f������Z����BWW\���U^v�`)�K����'P�`�r"f��i�eP�#F�<DDDDDDDDDDDD<Xp'"""��օ�/����^F׉�!K�Q;�B�@\\������hDEE!::F��J��>U������@{{;:::��ֆ��6466���f�yD�w��Ѻ�%��~	�&�3�!z�5��[A��ς�UO�	���3���[]�;<<����+�~����h4�[�3\�$�b��������hooG{{;Q[[����Q�|l�P��è�a��Sa�u9LW"|�B�݉B���m�A��W�U��-�E��ш��Cll,������DFF�h4BG�*;�f����hiiAss�_����eiC۾�Ѷ�u�Vj`��Qs7�4{��Q�,������������(��NDDD�_d�����?�}���3""iiiHKKCRR�B1
�O�� >>���ǭV+���p�̙s555p8C>�d�F۞WѶ�U(��0�ހ���!<{	˛D!��Q��O_D�g/���؈���j1n�8���"11��GX���qv�c�� �8q⹱�?��/�$I���D{{;�f��B�����z��=�����&.1�G����Ħ�ƧED~��1���h��*��>��ٮ�z�iiiHNNFJJ
RRR���8�#�`0�`0 ))�Ϙ$I���֢�����C^($���<�:����ߎ����`�SWBP�ǚDDDDDDDDDDDD���p�V��_�����l�qA@tt4������� 22r�z�^�Gzz:�����&I���Q^^���2������eH�u[;����h��yh����,��!z�?"�Yr���;h��[tzk�eMQ�����'"##iii����`�`zzz��j�f6�L0�L�͑$	f�����>ZZZ�v����
���!���0�,A��o"j�5�/����./D��ϡuϫ����>Nbb"&L����Lddd !!!�'=E��"�Y�f�����������ĩS�PSSY�uL�aE۞?�mϟ�2�!j޵���6h����i����NDDDc�,�|�#4}�:��	YZ�-�GFF"!!���HNN�F� tvv��	8X�-�&''c��� ����<y�܇�l��l�%8��{P��}�*��݆�EފOD���Q���A�'����v��)))�<y2&N��	&@��y!��ڿ?�z��sDQDdd$"##���.I���Q__���444����a>�1�_���nB��mPǤ���!"/rۺ����д�װ�.�1L&rrr������lDDD�rJ����ALLfϞ �X,())Aqq1N�<����A�inB�{O��'a�� ��i���՝�����������(D�]"""s$GZ��{4���ꊇ|�шq��!99���P���EDD`�޽�?�H#���H̛7��̓,˨���ѣGq��!TWWjN�eG�篠��W�9	��L�7@>��h(��G����h��EHNې���0eʔs�V�t���;=�[z���G||< @�e477���gΜAKKˠ/��4��34��8"��A���`̽xع�h�9Z����h��w�l�!�?))	S�NŴiӐ��;�������|�������ȑ#8r�JJJ I��a9�,�>�:z�.��Ko�����DDDDDDDDDDDD�E,�ј!�,h��w���#p������HKKCZZL&���)I�X,0C�A@jj*RSS�f�����СC(**Bii�ʛ�_��WC����w!v����LD^&��<�.�y�c�z�yyy�����ɓ�T���\p���qqq���ìY���Ӄ3gΠ��555.q�:�����YHX�D\��#���VF�ۏ�mϟ �� Fdff��� ӧOGdd�S���,_�˗/��lFQQ
QQQq�畎�j���>�����x3��� �Q)>JNDDDDDDDDDDDD�)x�DDDD�䲴���_����಴�~&�	����8q"�F�έ��w�^\|���m�d2aٲeX�l:::PTT�������7W����Q�Ə���ۈ_��&���这�}��׾�������J�30g����@���1H�������{��:��&M¤I��p8p���A�ݻ+���W�.y2�}���+`�P��]��Ǐ�� (%%�={6�����.t�F,]�K�.Ekk+
QXX������.;�w>���1�7#q�w����Qj"���2��fw���n��R� \x�:�l��f���:����눈(���NDDD!K�YP�֣h|�	�m]����`8W8n����F#Μ9����Q9^����<�gMM>��S�۷===���Ղ���E�O q����6*��R�]�c�������A�g�ĉ�7o����j�����9�r�W���s�{�V+***P\\����e�Ԟ@�6��#a��,�y��l/j_����>Z�ӧO�ܹs�����t�-::�\r	.��TUU��O?Eaa!�v{��9Wt��yDͻɗ?M�x�&"
5�8]]嗳�ш6��.�p	�o�����/g7L�5i ~9=�W��NDDD!Gv;���oP�����x���("##YYYHNN�0ʯ�
N�<9�
��-%%�^{-6l؀�������7N�>=�}����~�n4���.�1K�@P�|�h1�؉���Cw��A��j��={6�-[���d/�󟶶6DDD���z�������Ecc#�?����wu�;y��r�È��އ��B_O�1���h+� �������˗c֬Y�h�Po4���!--W\q��ۇ�;w�������ۅ��/�mϫ�Y��W� ��x&&"�����ln��;����� K; �܉�(���NDDD!�|�CT��=5�.8W��!++�'O��`�j���h:tӧO��y�F����`�TUUa�Ν(,,���h=���ߊ��C��9�R&&
]��RԾ��h����������/Ɯ9sB��Y\\�r�W���#>>s���ɓ'q��q�l�~��ԝD���8yR����3|��(����:    IDAT8Z�q�O�A۾?��.����|�rL�:u�M��t:�.]�%K����;w��ѣG!��o%��h���������A�%�!��>NMD�U�/��Œ;�p���~K�DDjXp'""��`�>�����g�k2�����	&@�P� ]����\.(�|
�e��[�~�!>��38�~��N��gk9sR���	}��(t����a4��s�.�秥�a���(((�(�>H�5550�L��q�^�G~~>�M����b:tV��������UpR��3����0-Q�V4��Q���H������T*1w�\�Z�
qqq>HH�M��� ''���x��p���~���3j_�M>���~��E���#"�P�h�r�Y,�E����bɝ��B	�UDDD��=f���A4}�K�n׀s���0m�4L�0�/;j������?��ŋ}~�@�k��k׮Ů]����CqGћ�<�Vߍį��6܇i���,���ߠ�������ӧL��K/��Ǐ�A��QUUP����T*����ɓ'���EEE����<Y�ж�utzI_{ 	kv@P�|�(u��ꗾ{���U*��7o.��Ҁ}�kƍ��o�k׮Ż�;�����u�|�4}��nxa�|���ƶ/��U����܉�����C@c����K�DD*Xp'""���Q�&��p�g��Y�f!--�G���R���с��HG	8�k׮Œ%K��`׮]��=�.-����#h��Ҿ�4L�.�qZ��bk(E���|b��N�0�ׯGVV�����Ҁ/������L�4	Ǐ����}���ݨy�^�~�G�����8-Qp�7����n������T*�d�\r�%�B�@����-[�`���x뭷���~wt�܏��C��o!銇�x��| p��g��NDDDDD4��r{i ���bɝ��B����C�ADDcס�+ѐ���d�ͧQ���Q����c�w^XX�Ν�E�L�\�P���������4rrr�h�"��nTUU�[H�l��}��R�g-��	�qڱ��XY����?	� m�$�h�ۉ��~��_\{cـs322p�7b�������Q�������旫|�(����GNNA@sss���.sZ>yΎ:�g/����8m�s��B�[��#uLD���1��v���P����5�8W���c�֭(((�F��G�.<<3g��ԩS��Ԅ��V�e	��=h��Ehb�A�<ٷA)d��ُ����;F@*ֆ�n}/��6"1N�a$���g��=�dt:<=;6[d�wX|��_��6�����KDDDD�U��՞^�&S�)�z#�_n?���%���*=��-V�������$�eG�m�|�DD��;�QPi��"�_�� />�j5�O����\(���t'""�������w��f0p��WcѢE�����Ç�;���W�y��l|��o�aJ��e9�*s#l�%�3�L��׾�9s�M��[�=0��B�Ѡ�� �������Q]]�y�,�y�s�<�6Ҷ<��k}�(���9���܈�/.87''W_}5���|��F[ZZv�؁#G��o����=�s�ע쩫`*��[��2|l.�""o	�r�Y�ɝ������O��,��NDD�,�_DDDD8;�Q�ۛ�y��祥�a��0>J6t�(������c�L:�������QRR�W_}uuu繺�q��[�y����[(�>NJd�u�����d���<�N�K/�˖-��@������;�h4b��ը����ݻa�x�a��V����!z�uH��3���y��v�����?��v8766�_~9���}���)//���صk���f�y��^�XJv#���p1��AVn?�%w"""""" ��g��NDD��-"""
xm�^G��������ш 55ՇɆ�d2����e�!������ߏO>�d�Bҁ7`)ۃ�[_@D�j�$�/[]1*��ݕ���������0�L>J�<���p��ƍ�UW]�����رc�e�M���/�R��[_�a��$�GKʟ�K����j�Y�+V��"�#�"�/_���|��/Aaa��y���>�Qs�B���2��3�h�z��AXn?�%w"""""�Է�P����Xr'"�`�w興�(`IN�_��;��w� ���ìY��P(|�n亻��p8�V��%h(
,_�3f��+���#G�x���lĩG� ~�H��QJ�S�k��"�~;${w�s���p�5�`ʔ)>L�zzzB�X�Ra޼y?~<v�څ�����͕(��R$���W��B��D����+�z�v���������M��d�����p�B����hjj�8�m����㷽���s|����_���bɝ�����Ʀ/����[n?�%w""
6��yb�/���Xn7�X�v-�̙t�v ����A�d2�;��-�����˲�������[ {S��Љ�?�3ʞ�����o�]E�Z�
>� ��8p ���1�"..6l����!��k��B��?E��+��l�qB"�sۺP��ͨx����z=6mڄ���1$++�����j�*����ڛO����'}����[���2�[����"�	�Sn?�biGs��\����(�pw"""
8������X@�2e
�̙�2���h4����D5L����4i^{�5|���tW�ǉ��F�� "o��y���e?߀����IJJ��͛����`A��rA��*�J %%;w��j�8���'8~�LL���0LZ��D�ak(E��/GO���M�6�]w]��(��T�s�����?�������@�Kw�|�cd���H?$%�`!�rȕ��:���$�;	��rȕ��:���$�֕m��(�w#����B��r���;������Q��X�x1233}��{�j5<�+V�;J�
�M7݄3f��_�X�tY�P��K�|����^�{
��������f�8~v���k��b o***�^��w�HJJW^�]�v�����g{���W�����D����[�xf�֎~�h�Zlܸ����a2
T��������׿��v�� ���?p��矡O�D�*PS�B�����	����DDDDDD^SY݄�����.�.� ""Ph~&""��㲴���+a>�q�sbccq����Κ&�	�������w��������<���(--�3.Kn���>X�� 󶗠�G�!%��ɒg^�6��y�sL&n��L�4ɇɂ�$I�Z�!�}e Z��W�Ƒ#GPXX��֛�ۅ���EO�Q���D��X @!D�Q��GP��� ���e'N��-[� ::ڇ�(ЩT*\s�5�<y2^|�Etuu��ck(�ɇ�!���"z�7������-��j�w""""""&Y��������D """�՗��Cs,�O�:�]vYH�A@MM�ǒ!MTTv�؁u��A�g����7q��h��q:���l������ӧO�<�r� 9r$$��F^^֮];�������?Z
gg�����օ��֡�{�-����.�۷og�������|����%���uo���;�DDD�W���8����5��q 
�,Y�y��AC����dBaa��c�Q�v�Zl߾F��㜞��8��\tW�q:��s�ס��K�Q���q�B�k��[�nEXX������VG𫄄\y�HJJ�wNw�8q�,X��0��8;�Q����8�V�s�mۆ���
��(���c۶mذa��œ��ڿ<�򧯅���}@"""""""""""��-1"""
xͻ~��������z��֭CVV�������Dww��c����,�w�}����8��l@ɏ����{>NF4t=g���C��]��{�˖-�q��U\\���H��;�V�5k�`�����q�ע���y�]&#���׬����3~�x<�����M� X�j�n�
�N�qN���P��
8�M>NGDDDDDDDDDDD�Xp'"""���8���!��ǣ���a�����8����z�۷��1B��d�=�܃���{wۺP��K��ѯ|��h�:������ ��j��&L�}�݇����8Yp����w��!�".\����{ޡ_>^>~Zv���tDf>�1N�`a��� �`��ر�[hئM���}�{�^��r�3�|p.��>NFDDDDDDDDDDDzXp'"""ߒeԼ�]Լv/ �����`ݺu���>�aaa����w���T*�y�flܸ�cqS�ܨ��V���'~HG4���7Q��epۺ<�/\�;v�@DD������j�\=���Ŋ+�T*=��.*�M4�󄏓��m�k8��j���EQĆp������M4X�����{����q��\��/EO�I'#"""""""""""
-,���Ȓ�����z��9���X�z5�j���R�cǎ�;FHZ�|9�m��V�q�����.� 
�����'7@r���	��u���뮃B��C��v�ԩ~w*����^d&˨������|�ȃ�=Bų� ���z=��.�Z����(�i4lݺK�.�8�h�A��R�׷�������������B�DDD��ˁ���E�ǿ�w���ӱx�b���~�͒���������6�F����7��׾��TD}5}�+T<{d��ϘJ�7ވ�k��!Y�kii����/�����Ω��C\D~ռ뷨xf���I ���Ď;�����d4���k��7n����eiC��+`>������#"""��%7*~�m�^�wN~~>


|�*�577���\آ�IMM�w��]���y��aT�p; �>NFԫ�GQ����,����ؾ};fϞ�d�����c~!�`���a���HMM�wN��?E�Kw��|��_���n��8	 III���{��%˗/ǭ��
�J�gL�YP��z���dDDDDDDDDDDDD�����Wɒ�^��=��;g�������a��g4�w�^�Y111�����~�oM>����q*����?}���h�=�܃����8U�0��0��4T*�ϟ?�������%�T�;����o���"11�7o��d�q2��O���[�B�V��=(}�2t�|�dDDDDDDDDDDDD��w"""�YF�﷢mϟ���p�B����0T�]]]���.Tn|�)����>NEcY˧@Ջwy;�(#%%�ǩBKQQ�J��c�F�n�˖-�wN�{O��o�.�Y-�~g^�����իW���~�!�V���X5e��s�=�3&ٻq�KXr'"""""""""""܉���;dU�����)s����ɓ}*�h�Z�;FH��t�뮻����q���᭟�8�E�_��{ K}����~qqq~H:zzz<�K������Y� 6n܈�/��߹u�?�������}�߿|��\nOMM�%�\�J�R	�Ʉ��"B��>�����tl߾�ߒ{�c��]��n]G *�� ����!�ܟ!�ZA�e)F��s��m6nW��ݽo�;��̀�������_������7版�]�k����g�/((@^^�'�ш��j�7��QB�F���m����O�������W�ex4bo�C::����_^����->>۷o��h�C��r���t:�*.��@�UE���*(�J����׼v/���.�՗1i�<�.�yd��q|ܸqX�b������v�Brrr�ڈFKjj*�oߎ'�x���獹��8��jd?�)t�\�KDDDDDDDDD�DBd�:��F <�?�7��v	E��w�Y���՞;��vA��z��Cv:{���/;���/����)lk�N|�D�w3��8�)b��8�	@l��x �4�������N'����rs#�|���k�[ψs�C�O���Y�0}�t&
^�(����w/S�ո�����_��N�:P�q��7C���i����e)��[�t��E||<v�؁��H?$-.�2����@~~~��/��rȲ���{��d�;��10;�)i,���EٓWBv9<�gffb�����/R���.|���6m��A^5P��eié�W"�=PG��)!���ALI�z{�1q�zb���*�_�^����;�z��-M��
��@nmR&�`ł;��Bb2��4 &��e@0F�;Y�J$$CHH�8.w�A�,�\S��rE)����W'� �q�-T�|w��yyy�9s����(:t�����N�O>�$�����%7*�����c&��K>�倠T������J���rH���cccYnEEEE�����T�V+���=�mذ�,�����;(K�xf��K�a�</��pz>V�[}	J]���q|���X�lـ���A@TT*++q��I̛7j5�V�;RSS�o}O<�lgw������O\���?�B��q��d����Z!�!��!dL��>��[�<BR
0��|M����=~bN��+䆺�>ae��2��27ӥÂ;=�aR��)'M�����t�C���0� �Q��6�U�JN@>uR�q��⿐DD���r?�����q|�ԩ�;�?��`�����	�J��(!M����;����>������$�eO\��?�u�wԗe8:��27C�2��_��eiéG.�����Xdd$��n��G�$I����h�w���v�1mڴ�lذV��w��3&9m(}|=&?���	ފه����3�&L��5���.KJ[Ww���I�&aɒ%�X�U*�0سg�Z-


�|��HOO��ߎ��z
.����������0�;��|Q���{S%T�	Py5"""""""""
M�V�eB��W(L�!,D�?��{����ˡ��f����Kz;�r��W�� Ƃ;!y�����@̚�X�G��0i2�&��Y� �9���⣐����;������as���4i��S����p�ٳ�/�w������>�(ZZZ�sv6�������n��'e���
�m����g�����yɻd��O][}I�1�N�m۶!&&��Bӑ#GXn����~
��M�6�j�����ϸ�����G���Af�V�^�{K5\�V ������L�d�eOn�����xzz:/^<�b����}���>	���>�c�'++7�|3~��_C�����'>���oE�Ϳ�Ygg��u�eζZ(�����!� a��S!fM���2���� !.�?���vHg�G� �T�;"ѐ��N�O��0)��9��B���R�E�i�@Z&�r- I�;�;�`!�ғ�W�D%"m��eO]����x^^6mڄݻws�P�Thoo���� !22��ַ�ӟ����/ڰVF�/���{ބ *�9��I6lM���s���ۡ�vB����y��N��&�O��s�Z�Ɲwމ��T?�
]mmm�������e��ك�+n��tuu���o���$ʟ��w�b�w~� ;�5�Cr�璋��Ns#T	^9'y_Ջw���'�RRRp�EA�J�L&477�������z���ӧc�ƍ�ӟ��g���K���Kvx5�,��h�:��,��Z��+m�&!yęsg@����~TЊ0A�� ���?���!�t� `���%Q�P�cx��!������lWo��ۡX��,�0'|� �1k2KV@q���%	BK��pM\���<Ǡ���7a>��Ǳ��l۶J��������Z�]�C�P����Ǐ�w�1�`0 33���}vܴ7�Ar� b�
�����{sd��gL�[�2��tgb{c9d9�C� mbp]��_��͇��~�(����T����tD;<�Emmm�9s��+
̘1ǎ��l�3no���"b��ь	 p[;ak,��r��l(�L^+�{�l��d���|C��I����;Ơ���4��S�c			X�z5����wZ����DRR
�-b����j    IDAT'==����}ƺN�!k!4�^9����Pz�@�١����!��ُ����u��p��k��X�ӆ;��JDDDDcW�ƀj���1��-�eG����1h�T*�3
���j(o���+{��q	cn��a�� �ˀ8gk.�09�!r[3��s����8P,\���B��� Nˇ�o>#��BH˄b�(V���2�w���F��) ����yo?�q,>>;v�N����B����>ea<�V�Պ��(G���������>u*t�9�wBY����Ά����:���Xp���(�Z��6`���~H�<x�{N||<����t�J��S��/���n�3n)�]rt)SF'�,��Q{k5 ��Osڡ4�s	�G���.T�z�����H\z�^](�T*�V�Q^^���N$$�* 4zrrrp��466�? K�<�/D͹ʰѽR���{c�yW�*����'C��c����DDDD4ֱ�N��� &�&M��k��u��CH�4�Yӈ�"���y�P��b�L:=���Xv����;��f�b�
(�q���1�h���5*u�*��K �\11��z��D~{p���Fų���Z�۷o�S�NHH��'X8&A��Ѐ���J�#���p��(--�3�y��Q+#INl�p�+��ۧ;��>rNsN��b�����͟?W\q�R����j��n>VA[[


�u_�N�	&`߾}�uy�����(G@v�`o����z�.;�0��Ypgg#J^	wO�+h�Z�]�aa����Z��$I8~�8�j5"""|r^
m�  //G��s��у��O��z
��O&�pt���V���@�s%�Ѕ���Ă� Xp�`ǂ;�u,�S�c�=Ȉ"�)Ӡ��5P�r7+.��1Pyo�1M D�B��e�}ʴ޿�z���J�D�;���1�+���!Κ!&��v�j��!.������H���	�B�.܃���%?^汌+n��6�?��}�J%,K�ä��PWW���$G3���P[[����wV��6t��F̢�#*�����k�����������YpYr���W�Zu���ĉq�-�@�U�F�_|��TCd4?���L&DGG�С�_������z�*Ͱ�/9��7����k��U�oQ��>|�ۅ��ף��X�1�R�5k����5:�]]]())A\\�Ww���A�Tb�ԩ(,,��q��>gg���0�_6�s�n'��pyXT���eX��O�2�����66Q��(DC�va��:W�"""""+b]v�Ԅ����(��]��Y_��+�By��ޢu�x�ټo	��x�3
 ���q��- 7�%?`��|F3@���o@�_ۻ�J�7��N1k2��C������/O4�XpR���_^㱬	 W\q�ϟ���#""PRR�6p�V��j�"..*�(��H$rssq��aX,����쨇����/�����zf��w%��v&f�}d��� Z��B�ۍF#��n��z߇
q��Ͱ�l\H5����3gΈ��RRR�t:Q^^�g�ei�����C�b���
{cd�5��ɒ�(B�5��Cł��վ��h���.��b$''�8�� �V�3gΠ�����\�D#��鐖��}��A���?k�!h&A�:uXǖl�J!9mC����œ����ie	Sl],�SЉt�pS[��� �����(ie	��],�S�	s�pS[5�]vG��|�[��-P޴b^>�8�B�8(]��%�F4�v�"�`���NL˄��-P�ݭ="�ߑ�?� !.�E_�"�j���w2
a,���wG�O{�5k����#&&uuuPr�Ӱ��j���###��Q��R���l�ݻ.������%O�.eʠ�'���7��eiv&�a����,����g8���,`P(ضm�_K��l߾}ܽ}��j��}=fgg���---}�z�ZyS�`o�������Jv+���������y�mT���c�f�BNN��y�R��R�p��)�l6����;���(
�3�Qs��2lh??sv6��r�0w���6(t��û��b�}`,�S�a�������|,�S�a�=���P�Z��@�r��q 7�	\#��W������0w�;�8��k��)Pn��o�!-��On�����7���HPS�fY�����z��O�P����öm�UZ�h4���f�}DQ�Z�FXX��������8x�`�1��`:��3��5��,� *�5�����l�<r	\��>c7nD~~�R�>�ٌ��(��cк��1gΜQەZL�2������>Ι���y�B���)��7����9�@������Xp:WWN=����g,==.�C��i48�N;vaaa0�u 
M&L@mm-λ]v�a)ۃ�����Yr��|Nsӈ3IΞ�œ4l,�_�V�0�օ�,�S�c�������3��)X�����((�\�߅�?��}�`"(�2���R�Sg ]f�u��E!�K^ht)�P,Y�O�����@�Q��E�˴:(V����B��i��NDD~$ٻQ��7 {xsO�R�[n�V;���ܹs���5���J�C��;ƘSPP�������m��S�W��Z`k8�=:WHq��X>'��;`o,�s�̙3�l�2?$<�J��AE�P������p�z���v�����e�m�DO�	��ݣ������b��n������&�)�'���QUU��?�===��CAH\��0�L}ƺ�Q��_���[]1\��I�[G�XD1�����
�QzMD4�Xn'""""�3S�c�=0	����~�W|B7�	v¤�P��}(�ą�npI��;���P(!.\�]�A\|1��.�LA@!�ˀ�5��@��:����B wp.������8��o|S�N��DQ��j����xc�^���lFLL����)999(**Bw���K{S9�Q���3�,��\��7"�AT@��� ���е�7Լ��}n���ĝw�	�Z�T��f�����W�͆��|����L&������>c��j��0�OZ�g��� {K���vBַH:Z���д~�
���a��
֬Y;���x�D���HNN��E�4*�
iiiػw/�<�YJv�8u%�Q)�벴��X6j�&ϒ��]���<,��}�t�ɝ�:DDDDD�Ý�)P��x��t(����n���ܓ9��&�����F�v�U���>�M|���E�sB��3P޶B\����ӡ��ϡ����ѝh���EӇ�x�>}:.\8��N�<���%p$jkk�v��.�>�F��n��c!����}v햜6���_��h���B�@�47���n�s� زe��x�=o9p� 4��c��9�����ի����q��/���Ĺ?�nl�p��z%����(�O#�l�C��wz[�p!���|�hdt:�j5v�܉S�N�;��'b�ʕ}n�%7*���i�ʀG{-�͕^Y�(9�pu���q�<�N�hXn'"""">��@�r{`��A���A��_B����j�Bt,7n����@��@d=�F�_A4<���[߃����D�k� qFT?z��k �_D�Lv�Q���C�"<<�6m��sssY����H�;Ƙ3n�8�_���풽����܊d����bH��e�%7��F�������Ჴ��}�ʕ����C��A�$~/"�Á�|W�E-�]T>w K�V��N��c�jgG�W�O�S�����"�����]L&�f3>��#���g4x�ׯGZZZ��muŨ��O��Yv;ak8g�(_�+�_�yK�(X�!"""">��@�r{��R��zT?�b�%����~⢋Xt�a�W����R3�ǹ��Bq�6��NDD^P��a�+�8�y�f������			�Z�#:�X�r����]i}m�ʕ?~|�ۻN�B��?��V[c9d���[�������#���W�ܞ���u���!��q���?DV�u����d2����|�~���ޝ�Gq���}ffW��cWZ] 		a0 @H�+@>�}'v�:�'N�8����m�iR7��9mڤW�����i��I�Il�q�������}#�su�1���fH�������x�h�f^4;�}}�s�U�.| ��w�z��	��ִ^ZZ�K/�TB"{	!�D�ꫯ⩧�B*����TU�>��|>���߯cd�6�cC=�
�cC��1�id���zDNaɝdc!�����hzxOM��ܞ#�K�����=�wP.���f��k���O��跡,X$;�!^E��E+O���_A46�NC�FQ�^q=�o�ԛo4Mv""��ȁ�8������K.��/��<˖-��ؘ-��P(��{Nv�B�}�{���T\\��Kv�l�kY=��`�k�#3=5��?��i]Q�u�]��5����r��WH��,Z[[];_{{�iZ��(���P���H:;�����|Lˎ��~δ.��e�]VP�I�ߏ��2lذ�?���8�jkkq��כ֍l3w|Ռ�p���8�������;��"�=xoM��ܞT�����B��@Qe'�#��@��c�>�U��Fv�#,�ӹ��v'���Ǔ����:Q\�����uȎCD�e8��,��H��v�m�
�и9fZJKKq��a�1<���7�x�����_���2���vC�x��reZ<Y;�1~|�i�ꫯFSS���<dǎ(++�#������s�y�oN��D"��g?�k����m�}⻮�Ȍ�CO��12�闐�3o�jii�̙3%$r^II	4M��ի�o�>�q(�]���5k֛�����}�{n�"�D��"�=�DϤ�I�p�|D K��>p�������{lr���EK������sP����씶�����q7ʎCy�w:+eť�=�C��x7P@����u�>�Uh��*De��4D4E=����X�ܟ�ٟ!
�z�D"���[��%����_�Ó���Z444`���x���,�6��Фv���S��=����q�zMMn��f	�����Gv��b�ϟ��yKJJp��c޼y������O�D"蘩`����eI�u�\t�ȁ��Z�}�z8FGG�o�.//Gww7V�^�d2);�(EQ��������=�.��" �ؾ��qa�;�)�$Cy6��@8���
�7DDDDD��6���vɪj�}��>��u����N����|;|��{(�NC9N����a�!(E+�}�P��.i3꠬�b|�����(��0���Dv���c��oGv�\���b�M����t���P(������NnRU7�|3,X U=��k3|�x9=���k������֧����m;�]�̘'; `�߿c�^7��s�=������;^�uW��P������&��˖-{���Vs���ڟ�3��n ��{�����
վ�Ǥ{C������F(��� ��]߹�L?u��W#K�>!�� �=�={�����t�@�DP]]�w���F�o�z�A'|3pbНk��g��P�|o�|�܌�{��#,�Ꮑ2�+��C�cᆈ����YC���$^)*Ũ����~,�K�(P�;|���v�AY~	D�������H.�;L����������5r������=�m��9���y:�#�wش
�p�w8v�y�桯�ϱ�{AOO�٬��QTT�%K�`��ŖE�2-����Z#�Af�׵�0������ߙ���8ZZZ$$����ˎ�wf�r�GUU�`�477c޼yP�(��|>�z�
�m��k�����x��z}�i��.�̙3%$��������ׯ����eǡS__����H��s�G^�u�����`8=p̵s�U4��{��,���
��DDDDD��79��vyDC|_�h�� �/��
�[�c���vAg�z���	�_�z�}@0$; �4��x�wC�|���Y�w����<n�s7�t���=�ҥK�N�C�*--����e���H$���6��� fϞ��k\g�"�&L���v.�3�,�烦u�ߏ�n�MB"o9t�e�&��ۋ/���s�B!,]���� �@ ���zӯkmmE���#;:�J�L�F6�ʹ�LO���Ŵ����|�r	�rGII	��4�|�I<xPv�L�4,Z��gφ��hjj2�"Àvx3�_���a�Ԩ�S���p��~�%w�6DDDDD��=8ٍ�vIT�ͷ����@\��gL��b���/?Q� ;��	��C�;(��NC���oC44�NCD8�� ==fZ�1c.��r��_YY�T�otL��i������c��ŧ�5MCcc��תz
���e��cȎ���ݿ��zɴ~�M7!�JH�-;w��m)555�����
K�.E(t�&ꆆӯ׭7���u%�a��$�]9�����1�����߅WUTT�ȑ#X�fFF�N/*))A[[����\�����X��?���aDJ����p�$ITɒ;ل�"""""9x/Nva�]���o|�w�&;81o!|_�.�kn�0�w*�@������!���E��	�G�����x�3z�%�>�-��|'TUu%ǲe�X��ߏM�6ɎQ�4MCKKfϞm�󵵵���y�>�,1����� �HNˎ���6�G�Q\y�����n��a�1���� -Z�ʹ�hnn����-�EAss�i����H�q#&҃݀�޵�k2�}8���6���a,\�PB�ܥi"��n݊u��A�uّ�%���X�t����$ �l�-3�����Ȁ�h"���N��B�\�'��b�]!�^�6��<Q7Kv����?�C�B�s��ױU�aJ|��}(K㲣�W�|P����D�K��ˀa.�,Y�---��(**Bqq�k�+D�p��������YQQ1�B���ɴnd�X��\�3dG�,"9��ﾃ̠y���
��c�(�(9)%%%����|>,^�uuug�u�h�HĴ~��c��;�4F6��H�+��#?{��>���e���;�`0�`0��k�b�Ν�㐃E�ܹs1w��	�FRZZ���J�zf�'Pq���L�k�"�;M�4DDDDD����4U,�K���\���Bp`.I"�A��� ڗɎB��D/*
@�����Pj~�1��Ģ�|A"��{7�o�/L늢��[ou=O{{;��Y:�*EQ�k�.�1
Fuu5Z[[-�k�i��f�֏E���"�s���8��������s��-��@B[[���	��hoo?���V�"��z��;ls:k��y�
M�x�>t��{�zuu���;�.cxxO<���SY
MQQ�,Y����s�ڦ�&��Ⱦ-���j'�Y�$OXn�&rK�4Y,��ޣ�d���>%�	�7��s)'��0|��2�����e�!	Xp�Q3�G����dG!:�(���@��>@��S"YNNo7L�˗/�̙3%$�̙�"����rl۶Mv���(
�̙�/�pR�f-�{����C��;��s�w�Ef�״~��O8���u�V�81bR4Ms�����X�x1��x�i���7�p�����x�/�q��߀a�����%��_�h{���ڵk1>�q
AEE���QZZz^�>Z᳣�X�?��wC�Z>���m,���
�8CDDDD��Xr���r���wC�����{��B@��F�y�f��4�2�=DiK@{��@44ɎB4!���}�/�p��(D�3��9l��i]�4�x����Ԅ��i�/�d��$��S�5�����������)����}l�rz����`�	��elllRj:�g��;����?>�Ν;�VӉ#�z�:�߮�g��w;���������kb5���󡴴7n�ƍ��3���ף��e��,7Z��߆K/��+�9�ZI��%w:�p6���0CDDDD��Xr�sa��e�e���7�p��(1k6|�](�����Xp�!��|;�O}��Dv��i{    IDAT�sR,��k߆r�|�Q�<��/�\���,'��)���=���ذa��y'����kZill4�z+ܞ�N�:���,�\o��&	i�g˖-(**�#���iG��t�RTUM�`QSScZ���0��ߦ�e�{-�bCSs��c9����]B��
���*V�^��_]v�UU�p�B̞={J������զu}l�N�6�=;>=5�ʹ�΅%w�ȩr{4��������rK�4���%f_ �׾e�R�Q��-�v���q7`1�
��]0�/�򎨨�����z��dG!�c��o����5M�5�\#!��"�2���y������Gv��QWW�ŋ���M�8%%%�S���>Ի��0;6==���<@O���o7�ϙ3s�Ε��[��,�٬�y%�J���͑cG�Q���!
M�X�S�C�$��}�s1�dF�?�d�zн�M�3f���v�TTT``` �W�F_�Ԓ�JJJ��ގh4:��̚5�r���q�|���2C���rK�t&�ۉ�����˩�{9K����ݥ^q=|��<\�(g����rس��\�Dm|�(�岣M������^h��7h9�د�0t�zgg'"���Df]t�ɤ�y���c�֭�c�<MӰp�B477���Se9�=����#��|d�z];W�;�YNo��[$��-[���؝)��bxx�p��c
!0{�l,\����r�@ `9�����ট�r�s�������ǆL�Nm��*!��˱s�N<��3���jjj���j�S4&����AD˦���|d����-,��),��H6�{{��N,��IQ�}�cP��4�i��DY����53dG!�1Z����}��53eG!�6嚛�}�a ��� ����쿛�UUŵ�^+!�5EQPUU%;F^+//Ǯ]�d��i���Ӟ�y���ˍ"��>T��m=�D8i�&���'�gZnnn����%��004d.��Ĳ�,�,Yb�q��(���m?�DS�g��#5b��Δ��eIx:��!t��;�zEE�#�f��&�P(�u��a˖-���[̝;�r��TM�u4z`;�]�Δ%#�Fv��)���N,��p6͒�Ǳ��B�ԗ�\y��(D�&f�������Q�!,� ��"h_�:D��S��dR�����7�
{K�Dt=�=�Q�z"�@ee��DkiiA__��yK����C�����Ç#���~\�2��C�v��sY�3)�i�49���#��֯��j	i�gǎ�O"/t��~��ĉ�l6���W\���~e���d2Ü�>'���#���ŋKH�-��� �5k�`����� ��������c�ATTT����G�M!P��|�����Xr�.�ۉ����
K���r�{Dyڗ���!;
�}JJ�>��PV\&;	9���^�6h�3��Mb�l�y��Yv��ad��^�O�?���ͅ:R@��H$�͛7ˎ����48`�q���
�L�Kʆt�������wMk�hK�.���{���eG�+�a8�d��{�:r\�A�g�F��Z�p~�V���i�Z�}�Z ��9s$��H$���.<��������g��.Mq׏���Y����rM&�,�ܽ��v""""�������Q��oA4��z*<�����B��N�Q�f,�
E�v�}P�{/`㣏�r������o@�_$;
QA���?H�5�ϟ?��l3g�tdj�����ct�<��N:r����l?n]]�iM��a^���Yf�0W�U�Ǝ����3�_y�Px��]�v!�Ȏ�W������������y�JII	���L�K�ah���L��a��dJ��������@�4	��KQTTTॗ^³�>˧�H�J�p��a[��QRRbZ�ڃ�M%B�z>+��#;:��y���%w�`�������0���,��GY��G�����9B@}ǻ�������ME�v��P��^v"W����(�q�Q��^�S?�\���+]N29˗/gA{B��{�9�1r���ؿ��ǭ���,�����SDʦ��;~�B���ߚ6tvvJJ�-���!�466:~�={��p`��&��˗#��	��e%3���y
��'��r��/t9	��v�Zl߾]v�:x� �����n�̙�5CϢl� fU�m=�D2��or"�K�v""""��ƒ{�c��=��8�OeG!r�z�M�>�i@QeG!����4�'�rIn�l�/���/CI\$;	Q�?��/�1�WWWc�����P(ĉ��
�p��1�1rVWW�ɤ��T555��p��aw��bij�L
=�ô�b�
�|3�i����I���ży�?����?n�q��(��ik>��c���~�3ey���t��o��i����r"?�+#�Nc͚58z���&r���8p���Ǭ����89v�,������ `�� ��Xr/\,�yK�v���eP����ˎB�*��r��"��';
M�ayL�|�}�,��wq�Ѵt���i1 \r�%�L���+V`ppPv���i'y���E$ �1c�i�гXpg��Sӿ��I�0�_t��ݰs�μx]�%��ծ�����Lq���5�]q��H����u�����&��3?��3�����Dp���^�###��x����m}��(����p�#\��]�2�,���n%�K�v"""""oaɽ���|��D�2h|�<����( �3C�/���H.E����\}��$Dy�г8�̏M뚦aŊM�uuu�c�h4�W^yEv����ۋ��a[��M��JF�)"e�����o���ȴ��Ԅ��	i��ĉ�_34���AW��2>>���.ۏ[[[k��PYY������p���g�OLk~�MMM��4���غu+6l؀l6+;�'��Ç�zL��@ �:�*�fW�z��dG�]9�t��^8Xn'""""�&�����Q���G?(�<E�(W����=
�T�|ł{>�A��#���NB������@��:�I��F�H�5�/Y����Mͼy����+;F^;z�(t]�#g<x��cZ��2�]�[��s�Q>�`2��0�����K.�DB�y���(��u2B���f�}����C45��ͫ�街l=����Ⱦ�=��i�����IHD�#����駟ƫ��*;�'?~��}�{���())1��w�E�1���O2�VR�`�=���NDDDD�m,��?��ݣ\y�|��kD  e�"h�y�ɎBS�O��ߧ�1��$^1��� ��a���() #��G���>!D	 �(��7�o ��9I�w��8�g����(��n�O���/���$���ֆݻw�@5E�p�=�:;;eG�I��ݘ5kB��mǬ��Į]�LS[�'���g"ّ�"3?O��Y�o0���֊����%%�d2���b�1����.��"��;::���TV�;1���'N�8m-�቟?�`��S�cɓ��](�滞g���`Μ9.'����O>���VTWWˎT�t]��Ç1{�lێY]]�����֌l��#�����	g76�4��(?��P�;Ur���,�|4w>a��������?��P1}�_v���ݣ\r%��>��6ܑ��>�	��[�0lF
 E��u��E+,�P D T�O�B��dIY��_D��Ga�9#��	�OT�'>��Mv�B��:�� ��O��0�}�Tjgg�]'z������EiB4�1[1�0�% �	��G@&5}�z�i�r��M�o��M�H,��hz*++�c����Ɏ���@2�̫��n:t��͛g��EA4EWW�i�Q�Ue3�=8f۹�����o�Gφ�0�-Y��@@Boٶm���_����D���O�x����h���¹�#��Ev|j���ge��}��3-̘��T����{��Ŏ;p�E�u�!G�E}}=|>{ʵUUUػw��)��w�����; dGXp����{�a�������ފ%���r�{�eC��~Nn��q!��0^;�'Te/������v�d���A�����>a�a� �յ��$�� 2���g��('�Ւ/ڟJ�2�I�YF��0��B��؞L&��r�Jg[dohmm��`ә?��s�ը��D�D7�b �n�*8�
����_@߾Ev��4��w������8�<�fgŊشi��S��$`�ƍ���+eG�I]]]hllDQ�}�����6ܳ���D���o����� ������}���i���CBo���$Y��Ƥ>Y`xx}}}(//��BTVV�ȑ#���Z.���@pV�m粒`��_^�T�a�zss3���i�D"x����H$ 8��V�lG�Acc�-���������?m=�s ���7��n˹&��/\��9��t�����,$Yr�i,��������Q�:�}�,�O�A � l6c�����F��qo���Ə�<��S���� K�XjF�b)���%��G?����8��9ك����>�I(�/��$ߌ���S �Bl��b#�CYY�|�q O�� �q��!�� .B\�Y��A{��H?�;_���(�XM��D"�r�N�����2<x����0p��1ۊH�ɩ�>��35�d�W����م��ӷ鿁3&��B!,\�PR"�زe�AN���t:-���ȑ#�܁���,�����?}p��>����|׷�g�����.'!;���  V�^��s碩�In�s��1̚5˶���զ���g�DcU���w�C��g!��Q�M�C��Ê��s��DDDDDt6,��>��ݣ,Z
�_ ����zM�����lGG�Aف��1�w�?  /��bq:�� p�� .���yR:/�6>��?}�����+[PW�ʥWɎ�/���a�	�B�oii�h��x���7~`˖-�q��z�0.���������W�~�30���(gz/�ƴ^UUekyW�X,���z
�HDv���(
v��ɂ��."	!�Fq�ر��#� ����pvO�>�t����o��Mkmmm�4~�l6�L&c�S
]:�F[[����������w����}sMQ��G0h�pn�����@�Mak���m�2-��~��r�s!���@ww7^{�5$	�7�xU*�Boo/�Ѩ-ǋF�B�8���XPs��n��a��2G�Cd���8K�9��v""""":,��.��ݣ46C{�K���m�� O	!~���o��ف����u'�>�k�֭+W
!�3�z ��&�}��k���"�_�.;
�?��q���@�坲c亃 ~ৱX�Y!DAn���b� |��֯_,**�
�;ø@��t9*T�G��꧀��i�r����2=��qۊ��(����F������,ؾ};�,Y";Jα�� �����{f��e�5`�i,��L
�o�M(=pC�o0����KH�-۶mCq1oo'cxx�pXv �������C�N[[2�	���D`��OT�Ǉ���y�����H�2�744@�cP��(�F�x�W066�K/���lp��Q��+5MCYYN��L�¢�e�����[eٱ$*3�!م�C���KV���>	}�O�D����(ZG~c�����'K*1��!rFy&�ˆ{�w�Ϗ���(z�a.g�W'��7t�Q���`v�C�c��K�{Q��=��gӸq��B|jq.�`���<
��_��zc V������_|��9����y�6n��"�x��= �H���[�Fo�ߛ��R��'R9LY�v�}�c��0�]U՟���=W����tvv��%�_n޼��a�Mq7�� ���V���_F�k�c��I7����\ommu9�3.���^���%�����L��%v�  �@UUd�������ο��KB+�￧��m�9pƇ EEE���%%�d2��2���W6�ŢE�d�x��O� Nn2ܗ,�����{v4ɂ�����r=ߟ
D֊��PTT�u�֡���XLv����ׇ��1[��FMw#�A`�3�Kq�gЖ�LDM����>?�@��'����PܛAs��'��Շ�ʜ�9T�1E���>�Qr^Z(�Qy=�q�{����x��Q��� ��b=7�圃� ��=�"���iK0���g��ਜ�jQ)�jt�����L�����r�DI6�ƇeG)\� ��>D+e'�ENNj�����_j��l:::^�a�l޼���� ����>�L�Q�/� ;
M���9J�͂z�� E�%�lB|����%�����7x��~�x<>�H$~��W��z!�� ��+�(�s�}�!�@���¯Mkeeehjjr?�C��ۑJ���*--ņ����"�]���1�� �B����Fr��l�E�N���G�9jǎ,�O��� jjjd�xө'^ة��EEE���|>T��z+�q^+'ҷ�MkB���KHCn)-- <�䓦�'49g>�g:*+�?�J�8��3�]�S#���D�n�?����r{J	?�h�N=�Շ�ܞ� �[V��Yx=��s��P����M����v�¿T4`��zg�r{�P5�c�=*����/��6�ܞ��B�G�x5P";JaR�>�Y��f�Ir�q �	!����+c�ؿ{���VB#�H<��?�L&k �B�� �7����1k��$4��� Q���G!��B��q!�?��8��c��Z[[���B[[���x��`08�0�;l��)W(m	�����DR�zb���zkk��SVe���`�}�4M3M�����wYE������ch�p�M�옧��?+#�Ar�Ӧ�%K�HH�-]]]�#��00o�<�1L�,m�bu�l.W�u���H��г����:��򾲢�¶�Ԕ�***p��Q<��tv:x�:~�8Þ�����E��9�g:_p7YN�<�r{�c���Xn�},������%���ܞXr?;��sK�g�r{��
��Գ�� �B�/�#g���0�?�����b�dg�E+W����?��bWh5�_ ��Ε�!h��
��}.�+}�Q5h�x��9i �w5M����I$/��/ZZZR�D�?��x�% ~
����[���Vv"iv��r}���.'qފ+04ĉ�S����i�&�1rRww��ǳ��C�,����V��8�l�����=��9�4+�(��e.ٵk"���y�������c����!����bu�lm]��]��z�3�qr21�f��OY�Ϝ9��$$��(������۱n�:d���aRR����J�����A�(G(����:�'Xn�,�[c�=��n���������%wk,���ܭ�ܞ?Xr��z�MP��Av�\`!V!nI����x<-;T����;��|>�,�0�#;�l��ڧ�h��(t������@�[(;�l'�x�������O.]������x<�.��2c����ǌh��(D�\�1��H��ִ�(
.��B��8�������I��,cϞ=�c���Q�W��������)MAQ�s��Mk�/�1�͜9����߿_v����� ;�%�0��c�{a�H��ę����_��<VX�4KNPp�1c��I(�A�A<���ر�<ٟ&v��	ێe�q@��(�������x����r{�a��t,����O�r{~b��OXn�O,������Ò��Xn�?,��G�� �?$;�l:��*��(�]��~);P>kmm�J$��& �����\0�_c9���9D��
�W\/;�LI �� �H�ukk+?�Q"�x)��n�����͢����_�(�NB���gLk����8�������c�-EQ�{�n�7_.���" ˉ��h�����Ҧ���W���ϟ/!�w>|�0��&���/��]�}�TU�r�I�j������t���O�ք������rE8F*�5kp��1�q�BOO�m���p�b~�7=p���� �')ױܞ�Xr?����Œ�I,��7��Yn�w,���r{�b��$���K�6(�@��C��.-�X ��W����Qv�B���2����    IDAT���*6x�g�6�57A��j�1�-���#���>�	�1dI��MUUg������K$/���UB�N ���#E���>X|�KT�ƻ�"�s���`�	i�3o�<躗�v����
l۶Mv�����m��
��	ԗ����
K�fzjC�o0���.r�Ν;Mӹ�쪪�dG8���>d2[�i5���&�L��2����t�]{�:a~�BEEE�n��ɉD"ؿ?V�^���k�M*����-�RU%%�	S}G1��Ԗs���I���)���Xn�^/��ܞ��^rg��0x���r{a�zɝ������;����%�iP5h��<DE��$���u�#�]�Ƿ�S��(�?�J�� x�'��U��s��f�1�|���%�>�y�瓝�uB��B���D�smmm���#C,{.�uX��N(pʢ���u��D�I�b��	�Dↆ$�I�1����R���9ett�ֲ���jCG��c�9&�ei�dx�&����+���s�JJT�N�8a9��&688�ŋˎqV�a����'Zm�?>F�h�y�t��ioY?���)���3g���r��i(//�֭[�a�n:=;�xa�z��#�GI����y�r��ë%w���WK�,�/��Yn/,^-���^8�Zrg��p��>5�`��26���X�Ҏ��M��xIgggo<����- ~*;���~h��2P�ϯs_�e�}��jd'q�+��\�Ů��b���UB#����� x���LnRn�J�2�1�\�|�Ӛ��CSS��a\��0>�˛�����a�y����YD�4�����%i�'Z�4K�g���i�������c�(|�Τ�ş���J ())1�wWWWC��e�y��)�6Ozm����3\NB� ���c�ڵx��d��IN� �u�.Lq絒r���k%w����J�,�&/��Yn/L^+���^x�Vrg����>9J�"���";��Ƅ�R���D��BCv �jkk{=��B\�So���jh���J:�H�^{�%1�1ܔ�X8nkoo_#;����:�ǿ"�X�z_!ڽ�CD*d'!r���Lk����4MBw��aN�����"twwˎ�S���l=^i��p��$.	�z+Fz��s�a����ٳ%$���a�A�1�������e�8/���0��wBX^/�����V�ix�fӚ����P����o�[�W�!�J��t�	���u�X�k%����WJ�,��S%��
���r{a�Bɝ����f�]QeGq���+%w��K��GTTB���e�p۳B��X,�Hgg��0tR,�]2�l5� �s����/�r��cx�$u����.�1ܴ��x<��ܹs9J7�b�]�X�J!ć����2�y�;�����}մ���,!������e�	>�/����9%�L"���v<�2R&ٍ�.�R|o୆���pǂ�s6o���';F^QU5o6�e�Y�z�p8lZ�	fad�}?�����ʝ����z̘1RQ�B���
�w�����R�y�����m9����8�I�@}��EP�WR�`���zɝ���g �e��Yn��͡~^�%w�۽�?�)�/ؒ;�텯�K�,�>���AQ�~�����2�A ��b�Kc��+�Ð�ʕ+���� � 6J���=�hh���x' �����¼�<C����ٓ���[e���B�X� !������v/>҇<d��v���륂��(����#������<�ԩ�2��MV���j���	��,"���?�T�A�zSS��a<`||�Z� 9ell�x\v�I���l�!hvS#ƻ��z�3��y���`d3����F477�+���i������Cqq1֯_��=�>�Y�y�,)1(��ECE ��l��H�6>��h*Xn���P�,�����Zrg��[�`ɝ�vo)Ԓ;���Q�%w�۽�%�����
e�R�1������w��tkY�����={�t
!��������A��!8�M�H���.����)�X���jժU��9%�������+�<^D��n�Y��J�id�6�u�6[ZZ���';F�B�����u~Oy��E�P(E1ߚת�O�ei�O�w�Kv�@ �����-[�XN�����i�1&Ů�ħX7�̙����z�3��1G��/��n�\oll|��ommŲe�022�t���ۤ�+--���X�z5���';�Tv^+��-�dz�� �K�}�5z�m$yXn��t���Yn��B+����M�Trg�ݛ
���r��Zɝ�v�a��L�7B}�{e�pC�0�G���suGG�y�U�Vec���E�P�SEc3��=�5��xG �X����Ɏ�8!�? ��b1�O�)�	!�x<�]�/�lcD2��A���p���/��JKKQ^�7i[ZZ��r��TE"lڴIv��agIaY��� ~#ZO��t������3gZn>���f��d�S�ib�tK��ߴ���6N���|��$�`0���#��Ê�gadY�9��; �K.�\��tN�������O<a���|��dl{��F  �$O�:���2��H�۽�PJ�,�{W���Yn��B(����m�Rrg�ݻ
���r�w���>��?~w��0�%��907���o�1!�?���4��[���ʎ�I�+p���=���MŘ��X,��x<>";M_GGǦ��������I��	�-�d� ������z	I�1c�m��J����; ٺa�jڦ?3����oH�4`���O�;�i���NB�·u�V�	�4���aD"�1&M�u$�I[�iU��Ηbn����5EQ&�VVVV⪫�Bqq��O>�£(
��(^y��[�Γ���*����^�B���'I��)�K�,�S���Yn' �K�,���%w��)�K�,�K�'���	Q?Kv����D"a.�P�iii��b�!��p�$����!|:��xg�2��� �ke�p�.!ĲX,������.���d,[�~ �I���wA46ˎAd�����ּ\�\�lFGGe��[�`�?���9�0�v<��ovd��,"�e��N�ڌ3$$)|v~�x���X�x��Sfw���z՜��g<~�4�3?ث�������Ο?�_~9��,����~?�� �}�Y��⋲�ʮk�����̎��Rp72)��A�V,��)�Zrg��N�ג;���V�Xrg���*_K�,��)��T6�+��-Yn�SN��wy��.f͆z�m�c8)�X,vk<�D���~���E ����QY�wʎ�9�;p�r�|�W�$;�c������X�<ҍ
����1� =��8BQ�~�c���#���qdGM�^�� �P�%,:�P(�cǎɎ��,�B��3��*+��a	��sC�K�oߎ��2�1�J__���eǘ2���bUp��(Cf��������T��c�׽���(
:::�ŐL&m}

���d2<��8x��8���Ziu_�@m$`�9&bx}3���v:S���Yn�3�[ɝ�v��O%w�����Rѐ7%w���LIE�?E���r;�)+~R�����B��~@-��	 W���Ǆ��0䌎��R�T���8E����se���!�EӠ~��\������-K�,����H$����V 
}3
y˸ŔM���-[��As�Ώ�iؾ��� {�H��E�HϢ\u�I^��J`�������ڂ~����ݲ#��00o�<�1���{0h�@\WW�t�a[�s&�?�b��k�듽������Q__��>��@gWQQ�cǎ������ג\3::
]��du�̎!R�:�ޤׯ����i"�Rrg��&�/%w���l���r;��_0/J�,��D���r;Mċ%w���C̾@v��6��x<��� �����={��`�����E���O�f��û��o{D}��N0�x$�߻r�ʌ�0�x<�;�JuxFv'��z?PU#;Ѵ��.�WUU��$�!0s�L�1�Z4�K/�$;�t���aߔ��,"a��NӚ��C8���p�ڵ�HDv����ۋ��&�1�edd�a�@��fMMR��l;�#��	��Ǭ�S�4s�L\u�UH&�ӉFNQ��al۶�֭���kð����:	0ƒ(-v��@^��c�?�r;�U���Yn�s���;��t>r���r;��\/���N��%w���\�TrU5P�q���0c��(+�DAP%k�V��&�� ����"f͆z�m�cx��P[��w�N�Q!��D�a�AH�����d2y�����vEh����D�6vl�i-
���>\xᅜ:M]]][0:_v�6EAQ��pќ/	:�)�w�3�E�Q~@`�}��Ɏ�wf͚%;´麎���F��*���?�)))�2�e�9������uc<���zZ�mii���^�T*��qn����A�A�]�;w�7�g�@vt ᐳl�C�:z������r���r;��\-���N���%w��i2r���r;��\-���N��+%w�����3!�F"�����|��G���� ����,vSo���O�w�\���C>��v6�X,�3�AH��+W��ٳ� �$;�ݔ�(�q�1��e�k�im�%�B��ڊL��ީ
��ذa��R麎��Qێg5Ž��d��IF�ۥM H[L~������p>|���'�����ϗ�v>��.o���N���r�{��z4���E��+�x�bx~�]8���0�x�	;vLv[�u���4	 ّ�;<������r;MV���Yn��ʵ�;��4�Trg���"�J�,��d�Zɝ�v��B/���eP��dǰ�a?hoo�ܹs9������Ou]�@a=���z�=�Sx��,Z
�-!;���u]�&�H���rêU���X�C�a|[v���� �j�cMY��i���JB��TUUek9٫����^d��,mZ��ң(:<i��S� �wشƂ��v��ɉ��dGq8W�9���^�����=��V��>���������W\qf̘�'��9E�Q�߿k֬��#�]�V�& ;>�H��h��NN`���*WJ�,��T�*�o�\�e���#J�,��t�Jɝ�v��\)���NSU�%wM��݅W�5�o���G���@�N�����W蕝�NJ�bQ���wNRT��Wv
���qmGG�z�A(�!�D"�a���b'Q� ��d� ���y�ay9��}���΂)���q�F�1��o��o~sQFq�٧���N0�qڸ}���l-�z��� Z[[eǰ���J���Y�fm=�/oJY�+**ٸR__����
���>��
��i�D"زe6n��0dG����>���	@zje�W޾V�3Xn��]rg���� 𫰼�;��d�%w����K�,��t�.���N�U�%w�ڷ�u�c��D"q�"�ߨ%�uttlp5����I{߽@�<�P���A�U7@�7ʎa� W%	o������ �!;���w�(-��hJR�GMk,l����#ʎ�����p�����TʶcY�GP�t���S� �{ȴVV���l۶��o�'#
Y���w��eȍ��W7��M������˗/G2�����
O(���X�f���#;Δ9�qr�A
�z��s�w��Nv�Urg���"���r;�IFɝ�v����;��dY%w���.�Tr�Է�Kv�}-�?$;�x<�UQP��E�,(+�������!���;�-;��ø&�o��r_<��o��aQ\����z&��Ǉ����9�ݬ���c�-EQ�s�N�1�q���M9_p�(�{X��<��w{��� �3)1_#�Ɏa+���EEE��Ҡ�8[���2�<#c~�s�:���q��c޼y�����	����r���b������g�t]G&cO9��3�?���PpG�w���d7�K�,����.���NNp���r;9��;��d7�K�,���
����^ TP��ߍ��_��r_,�� I�Y좽��@q~_�r� �����Tv��(�r3'��d�b��
!�Yv��W]_�����?f��	�f��`���,LMC4�/� ;�v�6��HF&�����M��6���V�Xp�ǦM�,�m�Ą�4Mv[�1�=#3�l�ի����}ei�{�{D�Q\u�U(//G�k��#�@yy9v�܉�k�������2�^�V��Xn'��Urg����Vɝ�vr�%w���In��Yn'��Urg�����%wQ?���Ȏa!�?�b��e���ǟ�6 ���آ��-�d�(X��p�(�B��F�1�B������A(�!�ݻw�+��o�Yl����q��D��Nv[�����7zN�={6��OS?����������o��Y."eG���y���T*5�k�666�x<.;��t]��5�j@II	2�?�У���P�庌��9s�r�J '�A4�ߏ��Rlذ�?���8�ͮ{K�뤑I!��#Xp��b����tɝ�vr��%w���N��Yn'78]rg����tɝ�vrZ>�����(�����.��$A��x<��w(�ǁ*W��qب
�j�K�[V����'c���d����jժ����{��eg����R�Y�e� :o���}B!wÜ�b��'�v)--�s�=';��R��m��'��\$���<<������Gw� N� )�0A^�,���+v�I�L2Nfr<�<޹2��d'��ٝ�Lf'�����<;�d'���8�lk=�Eْ�Ô@]$ER$^ @�F7�W�4eUM���z���~����k�nt���|I��E�r޺��F]NRΜ9��c�
�B�~Ϝ>�"�����do��署��~])k#��i���02�J��x����؈@ �S�N�ڵk��<���@T��u��6���I���vr�S%w���-N��Yn'79Qrg����Tɝ�vr�S%w���-*����-І�ʎa����_B��@Z�T*������G���S�%����hm�v��c��0��J��O�9Hm'N�X2�'\��e�4�O���D�V��T��9;$	[�w~0;���\�1�=��j����\p/���p��$��\.�Z�R����A�1c�&2]�M�c���çV��>m٣'#��?�-[�`f�z�<�}�dw���/��L��g��ڰQ�u�Q."p�t?����a���fwɝ�vr��%w��I;K�,��v��Yn'��]rg���v��~A��{���X/�ۯj���;v��s�T*�� ~_v;�#�ZZeǨ;uq����?QeB�J��J�~[v��Tj�0��P���ؼMv�U)/gMk�p��l�Au�F6k����B!�9sFv�Ul*<V��tc���'m�s�	�@���uz��MwVU&�A<��1v�+�[Y�lhh@��d�5V�ki���@^���сg�y�Xss�N�'�i��D"��g�⥗^���Mv�+�*���A�_���^I��r;�bWɝ�v�Ů�;��$әX_Ot����r;�dWɝ�v�Ů�;��$KY��%wm��eǰ�] ��+;Շ�����U�9�-D�'Vv���W6��?���vx�0�_B��P���i���)��̗d� Z�ʒ�����
��\�d2�>�@vW�5��Z)��P>7����j2�WJ�*[XX�A)�J{���Qv�+�[�	%��(8[p�����T;�k��ݻw��ɓ(��XZr�g�T���؈���x��we�y�ӯ+�Mpw�-aç�JZ;��I����Yn'��[rg����L4��;���7�Q�a˦5{Yn'��[rg��dS���̗ ���e�0�N*��*;�!D�P(�"�7egY/��'���1�
_Y�H���*��*dF��ϧR��� T_B�+�9�K8�e��D�TY^4�U;����~N�\!>��>*L�9�XX����]�.��^+%��7X�2�t��y477ˎ����9tuuɎ�(�'���_j�����ҧ�J��� �܁{?��� ���l�XA�%�H�X,����͛7e����"4�?H�齒ֆ�v򊵖�Yn'�Xkɝ�v򒵔�Yn'/Yk���v򊵖�Yn'��r�]l�m %;�~s�n�u    IDATxx�y�!��=z4�� �.��>�3�S������'�?���U1�8pMv�_����+��+�9�E��)�)��R4O�d�}�v��a{�O��$Μ9#;�k�.�k��ol�yҦQ)�֪��hu&&&dGPΎ;dGp��ϫ+'� J˶^c%?m��(��@���o����O=�zzz033#;y\KKn߾��~������|p��^���kK��+�v,����Zrg����֒;���E���Yn'/����r;yM�%w���k�Zr�?�Ӳ#���CCC ;կT*uU���v���O�	�1�_a�D{�' ��<������";�7!�aƯ �,;�zh�� Z�d� z8�Ri�&d2�1�����|>/;�+���]x���"��?���:W�^E"�?�k1;;�-[�Ȏ�8��M�+��������&�����3�<�p8����q��� ��8�|�M����Ҧ��u�|�k�'���^I�`���j�%w��ɫV[rg���l5%w����V[�e���j�%w��ɫ�Vr���c�.D��_B��?r����s ~Gv�u	�?��)�_e�!�>����|����A��J��?� ;˚�����Dg���򲳓`�Ycc#N�>-;�+�,@YOpw�e�ߏ�w{}���#(���WvW�]p��_�.\�y3�������O�P(��=T4E4�K/���/�~}7����N���N^�aɽJ��v��%�j�_��I+���N*xT��v�K�����Yn'��R�]��O����<�r�R���{�fe!��/�α��g ����Ұ�����,;�z�k���/~�rFS�/�B���s���ԧ�� &�gMMM0X�X�H$���)�1g�o��9��	�������e0'����۷�L���Z��i�޽[v%Y�/�[���P���j��@ �#G�������|�G�Ǳ����|�;���u�����b�r��j`��I�
�,��J�J�,��J��Yn'Ud� ��e����r;��%�h��O˻�=~����o�A�!���J�_�챼�9��S�c���X/M����S�������u�9�����αf�(�㟐���!�o��=9�>�L&#;���� �~����u��^ta����HV�s7��֣.(Wx����Uv׸q2�a8��ǟ�z��܌�'ObÆ�����<���cccx������]ϣ��Qv��B�+����E`��I5+��,���>Zrg��T���r;�&����r;�Fv�]�4�I���/����?�3��α�g~
������:i��!��>N�φ���Lv�'!D�߃�;��O~�OF�]o���^;]����.;��ZZZp��E�1eWi�0�2R����Y��"���֊Ţ�$j���ESS��JYXX�������{�����apzk��k��>}ӦMxꩧ �����8�a�@ �D���8s挣?�nlr��%�d�Z��vRSQh��d/�Ś��nf���s��J���e#��3�8���s,���ƃ�߭��z,�r;))��q>Ҍ?j��r;)�,�,ً�n��5��Cs���~��"r����W ���k��m`Hv
��U�:i'?%;�z���_���-�J�0�_�αV��ھA�1�,i�q"���ݻ�tZve	!p�֭��`����
t[��|\D����	�BAB����;�u~V�H4u���N�-�� '�;BE-��e3��� >�|>_7����ؽ��N���˗��]��j�	!Pvxs��7NRuoE�,���
Bë�$�zPv�51 �nH�����#���x=���h�n��aC��vRւīI,i���To��^S�O-��+���Çߒ��|� ��b����Ay|Gy=ZZ��e!��'S�s�R���˲s��v��#Y�,v ��v{����o��$^�u�1cW��&�����οo�k��X�\.�hԺ K��J�d�p���W>/�E����O?�ԪLy��{e(±c���ׇt:��tzrVKK���q��)�7��u����R�A�7���^IDDDDDDDDt�~R�b������(;Q*��B���k��H����Xp_��'��ti�_���s��bƯX��e-��C|2"OңM����e	I�CWW�٬�J+�X\\����=��jE��p����"��d�r��M-5E0�i��B�v�P����
�Z��#F�O'��U���Tp����###H&������<L�d2�.��_�����+���o��齒������������*;�h����C�044�� ���cM4��Gd�P?mX+M���ӲS�U>|Yv�����d�XM���I�)�L�ྴ��>�8|�0����ʊ�b8}�������T�P�l8�_K� ������v+���b����R�4���{��{��Ғ��[�t3���@ l+�z����q��q�J%�r9�q����0����ꫯ�̙3�~<���^W�@E�7��}b�J�'�Qvh.��� ;�
_ƽ��ю+}?��߹5; ��.;�Z�ށ��A�R�P�] 7d�X��'}[v!��,&�
珣�c�X��ש���oߖ�V��A��)��J%��\х��QU�˂�����F�S���e�b�+��ϡ+_�d2�'��u*q�	����O�4:t�T
�L�'{�C55�{=��/��͛k~�6NV{]	=����?�>�WAӠFv���	���h�T*u��";�Z��{�Ɏ�,~ڰF��OȎ�V��`���Ad��ѣy!�o�αbC'�����z�ٴf������1??/;��� Ο?/;���,lV+"-U�):=�М��W��7�rb�e�E�1�R*�088(;�v�6�{�������'�ݟ�J��u%���@�hǏǶmېN�e�!�K$������?������}�^[V{~^�h�oz�뽒��������H�? ѶAv���g�T���'---�[ wd�X���]c�Xp_�h����S���7��	4)ipp�O�,;�Zh�������V�u6�G���^�1���҂�g�ʎa;�B����X!ۮQ���B��@CB7�w�Kqs=�~�m46:<1��d2��q�1����nU��f���}�(�l�f|6�u9�\mmmA4]Sq��C�4����ܹsx��k���h�]hȕ�?ȯ�J"""""""""���#��+CCC_����cǎe��Rv���RG���N���k��� 6��!�?*y��B�s�9�B>
pJyH(�sy����o�Ν�޹N���U���&��|nUp�BQ䊫/E���'m
�@�y�;��Qm*�
���+;��p��u�ZY�/3���	6v��2��\��F�={�����(��<�*#�⥗^Z��p8l˵�
�Z(�̒�+������c-!�?B��=������5�Ps��l,���v��#���'"R����<';G�!�d� ���hH��YF�����릠-Css3~��ʎa�H$b�cY6�P�%gք� ��?�����JH��s���v�Z��͡��Kv)�W���\�-���>=�"��0o�����B����طo��4*���H�a�x�B���w111Q���4Ͷ͓��p������d """"""""�/1�b�c��0�������Q�!Ŀ��c-��OȎ�$�X�@44B��/;F̈́����D5�- �5�#Oʎ@�`�\�[XX�������!��ˎ�4!D]l�������lZ�B���:����
�<���&''eGPN__����5��>����;Q����~)���2�@SSFFF�����=R<����q��)�r9���WV*�*�c�:�q�񽒈�������|M�kE��#;�j=@�i�bߐ�`dc��Fb�(P�C�0~[v�Z�R���a<+;G��� ���C�D�i�
�^q��Q,..ʎ��H$�7�xCv�usz���a>g.�ۊw�A,*V766�D"!;�Rfff�u�V�1��{��Ն�����2!��7㝦5�'���###���d2�㐇$�I���x����o׽��	 z��ï+�͓DDDDDDDD�C� ��òS��_�#;Q���� �� ��òc(��i��Ɏ�/�R���A���!;DM�1���NA��P�\p������>�B!44p��z��qܸqCv�u������dZ+ja��8��)�@x�6���쬄$j�z����ٸq��R�]p��_f*�^�Dӝ}|�Z��L��0��dsZ?�;�|>o9A��h4�P(�_|�.]`߽��	 Z(�tμ��n|mIDDDDDDDD~��?Dc�cԪ���I9�T�; ^���V�!%Oy�����Fh{dǨ�a�^v��>�۲s�J?���D
�o1�MOO���annNvei��a�GEBD�Q[kii�	�������!���}V���i�J%	i�mbb���k�N��{�n�1��{C���a�	g�8>�WF6l7��E�fc!�رcx��0;;�M �P�x�l�?��m�;�Mp��_ta�{�'���h�ʎ��L�Re� Z!�r�X�c��=��`���?����R��_�A�V�a������BȎA �t�4�ݽ{WB���m�6�֡��o����k�F�i����6is���8~/m@آ�Y�T�)�¹s� �Z�&����#H%�@,fo�|�=3�NCkl��+i����>�u�'�K$x��������H---(��s���ZT{]���s��.�  ��3���A����f*v���|�{�s�$�ֿ_v
��ӆh)�j&��!w���������&�$�f�X""]����B����֭[1??/;�����P,eǨ��������<�zlE_��&�����I�mvvMMM�c(eaa�f�H$b�f �޴�B���������v+"��{e�s��:�u�V<��S��r�㐇���"brrr]�����f,.9��[�������������G۶�9.;FM�o�";�Z	!!��*;G���!���j	�oPv�ZM477���D�e�rOFB�1T�"]�,�9��~CCCJ�����	�����5��ྸ�hZ�B1�-;?)[�w��#����Ą�4���;� P�T+��.w���{%p�������I�ڶ�z���~�E��;700�C�!���u#��b1�B��3�`B���#����XVw-�\Aw��)��+�����������0�ߓ��h��`Jv�Z�SX�^m�V��Z��!�hǎΞ;L�l6�U wd稅��V�z�	�x�i}||\B���H$L�d�6�`����cԤ��Ѷǲ*��fL-XOv��ߧ�g�)�����r�F��c(%��!��v�+����lz���묤����P�Fh��i��k
���O����tZv򐖖�Z8���nݺ���ս�g��]z,�;sο��������������G�?,;B�& <+;�z�8qb	�������w���`�}��zeU�0�?���'N�(	!�";G-Ď�@��E���t�4����Ç#��ʎ��P(�3g�ȎQ��&��ﵲ*�Zp�ႻB:zU�6��nܸ!!�7���"��J��=���-�[ܧ��}?�Xh[Lq�sG��Ȟ��ֆ��466bnnNv���v�u!"����011��	��|���cq�v����{%�KS3��>�)j"���T*�cF�.��8{t�ʹ}��Z,������ ϧR���C٥T*�Tz2�4h; ;  ��\�d���P�x\v�%�I\���K�X,�@ `�c---�\.��s��%g�[������}����I�� �X,B�u�1������A��������@����9�{+O�@�f��8(�>�Z�ڵ'N�@�\F>�|���kÆ����������L��چ[��S�<����������N��M�
f�R�(5��a���? �=�9j��mi����"�A`�.�1j�)Du�СC�!�/;G-�c�� �j~at��-	I�a���H�Ӳc(K����GN��;73T+"M#�]�6�jCP�R�=���G"��<֓��%444Ȏ!]cc#4���]Yp_XX@����k�$�  �Jl���^�T�yr�4M���144�L&c��ꛦihiiY�?a���-7�T{]lnw��q�$����<@��N��LT7��C�j����4L������غ�^�]3�X웲C�M��b�n��  ���y���IH��=�*����J&��㑚��m{�����pװ��h����PEl�  �i�ƍ�x�a�b_�R�����ˎ�	v�+�{�	,--=�v��uD{�m��Jz��J �YLp��7o���>E�Q?~����0�3���5������0>>��)
�
��p��u�|� !G�ADDDDDDDD�%�u���c���H$�@�T(mK��J�6�U�v��V_ۻw/(Tw���@`	��C��[�X�3OT#rS�{7�p*��,�������Ooo/��}['|�M>�G>�G4��*;��Z�	L.-�i{��O���c	�Z7�0}����W�����rBy�[o����F�1���dV=���%	[/�ɘ�n��Ad�v[���y���M�-�mZq�
�����Fww7Ν;���i455ɎD���Xӿ'�@8���̇�cUpף͸�5?%I㽒�C��Ql۲��mU|06���ң�AR��kؽkl>��S&&Ә�;/;9hg_"���da>�k7�d� m�mG2Q��E\x�'�ճ��ftw��{��a�¥[(�x_��E�����ɡ�ݼy�y�Y�C44Bt�ʎQ�\,{Nv"��رcytt� ���,�%v��\���Xp_m�Zw�0�Rv"'>|xatt�o ���,��i��C��3����	MGl� ��_}`�wg��ٳ�ò�(����O��l�8�����0,.��<
4���U��T�8���}�1���~��Ii�ann�vjP�T�g�ZC:E�4�v�
��М}{C��	�+Ɇ7l�����?����:����J�O� �B��]�zzz���~t��7P.�?X4�a��dw;�^I�c�]-8�ߍ����P|el�l��:	��ow;z{��|ҙ�&��8�Xp�s{:��7�`��~�s%�{~��:�oO7�nJ����ӞTP*U��{�,�׹��;�gW�Z�o��ax��n�� =����$GgG��t���>?G�v#���"��$v�b;��ۻw/o\T���!�B����e��>��R�=&;E-�f��e� r�R8T;���Wö�i�E$gq���E"LNNʎa���̙L�JŴ��1�pY@-�Mո�q����,�鴄4�?�����itwwˎ�	����u{?��:�bʰwJ�N%��ƾæ���q,-���M�p�����#�N[�f ��B!�����X�������6ܜv���{%����3YϏW�0}�����(�P��֭,*p��ML�q��-�O6!�4Q��;s(���b���n�R)ɎB00;�F&[_�J�s�����(�\vӳΟT�&�0p��23���*�,nݩ��յLL܆����2��	��\�gB�S �y��ݖ��G����:�_;q��Ѡ�����- y�9V�OF�M��0�]�~��2�t��!�"�N0�;�#;��d2i�c��[O�����"����>Դ��_��߹sGv��رCvϰs3p�ã��'&&PNn��:+	!��s��ZX���T*���?���022���n�n��W]]]��Ds9�\�͝��v�d ܉L��~��N>Rg%���v�U���uUr_�q��T���U����������e����J����ٌ2�9�A�������Z��E!���*�M�    IDAT�)�T��Y�9VK���(,�?�ء�N�o��@�cǎe |Ov����v�vթ�Ǟ4�X��H�u�c(���.\�����:�ڪ���"/8_҂,!�ݴz�ٴ~��%	i�v횭�9�`vv[�:[�V��??�L�r���K�.�a�>[���F��#�{�rݯ����Ӄ����ad�,�;O��*�-�Y4#��|��w"k�Rrg������r��K�}![ą�7Q)�GI�jQ%w����>J�,��[���Yn���ClSg��T*��2�C�֝U�غ|�e���X�B�_�u�k�V-���n+�/�܎h�^��ŋ%��={�p��:MLL�R�Λ�����M٬T*�i� Lt��S6�1ǯ���h�qĴ~��9	i�bY�v����#xF,C,f�=��ċ�Ӌ$�l��JZ��ʏ�t�B0n��w��e	i����G�E6�E��鍪�4Ͷ���e����N��8�� �o5U�zɝ�vR��>1�ǵk7Yn�1�K����FE�r(���%�R��wYn�9�K�,��~ɝ�v���^ �c�*�ʷeg rZ(:`Yv���6o������#h�����wZ�躮N��ظEv" @��5�MƮW�������z���8}���jkk��,���h+��Y�����w3���iLNNJH#��Ą�'����v��.�����m̹�9�ڤ��\�it�J���0-_�z��ʼgX�� �|�I�ٳ���05�:~��ىp؞����@0х�)�J��^I�h��ܯ�ͳ�N�(Zr��ܮXn���%w�����,��/�Xn'EK�,��G�Zr�v#��I�]g7պ@�u���b```�+�s��b�XpѻYv�UB���|����(3RT��T��v7�]�vKK�}�����N,.:?�����eO|u]G2����fgg-ׯd#�T���M�S��������{��ryΝ;M㟋�H$�#x�����{'^,,,<�655��]�^Ǌ�ҦI��'Mk�R�'?H��q��I���X�t@޵e���z��צ,�f'�+�VG���ձyܽ;!;y�b%w��i%�J�,���Z%�b��;g�Yn��P��n�_�f���Z���r;�c�Nl�";B-��.;�T��
��oK���C�d+��,;ƪ	!�#;����y�yE��'!4���r��)�.9|�07�C4�����6[K�Vw-܀ky��Z���먨a���L�gϞ���}�tMMM�c(%��bppPv�hhh@,f�},�N�N�x�wۚ��:+	= -q�*����废6yѶm�p��IOl���4����=�U�]�A�)ư��|q@��N�Z���Yn��)���NըRrg���S��^,x��-��@�-j��?,�/X*"S���r��Tvi�2+"��� �%��@ܾ�����Qk��́�P$�0�e�VKc��<"�؊�GM�����4��Fe�PZcc#��ǥfhoo�����M����`*c�u�a	�!���=cZ�x�b����w�A �C)�P�F>�a�y��zYm�2[�uvS�np��U��C��<=�wo�����fQ*�dǡ*zzz
�ly���e��֡�\�t~�������!�'^/���N���;���(^/���N���;���h�.���N�����؍���m�&;B-��X�����9 �<��W�p,�?�J?<�a�*���`0�}�V�mu~/�j$?gZ{�wLQ��T
���c(K�u�ŹH$�dҾݳVeM �kđ�-�v�j����i�\.����Ҹ'��!��Z�r9Ɏ�BW
��bw�=�_g%�+�K���i���ۘ�����V�D"x��'�}�v��i�q�B__�m���f-�Cm[p��p�$��x���r;��GK�,��jy���r;��7K�,���y���r;�«%�����`��A��hi�cՄ���@�!DEqZv��R�4XpѳIv�U�������ܐ�cU�������[2�y����"�^�*!��h����^�1���҂�g�J�vgg���7==mZZ W	[�cE�S�*��g 4ݴ��[oIH�3g���a��z���j��#�ɠP(<�v��Dv|���Xai���s���y�����###����h�!�X��ݶ=�u�]��ԅ;i�'�s3��y��~��v���J�,�S��Vr_ȖXn�y��^(�Yn�y���r;���J�,���g��ɾc�T��Dn�T*��ΰZb�f�<����-19�G��)�d��'T��}�v�6��������Ν;9Es�fffP.�]���=��Ғe)��ƕ��mשF����m��@Sw5��;w�T���b��?kQ(8�}�7��΍�A�þ��V�Р�yS5M��������қ���p��	��e,-y�H�W}}}6} V.��ϛ_?�0UD�����:�D�╒��y̰�Nkᑒ;��V^)�/dK�x����(��e�=w��vZo������,���x���r�{DG���&�`���H�N�beױ���]��
�7e� r�ao�ΰZ�ݾR$�z%�>gZE��	~044T�Y7455��^s���d�։�SSS��H�g�&p�K�6;~�z�<�����r�N'>s�"���JYZZBCOC�/� �L���+�a�zy���YI�6�o�T#� ���i��իXXX���E��b���H�Ӯo�{�ؾ}�m���faX|hj݌s7��X+� O"���;��n�K�wXn�u�]r�_n��Yn���[rg���O~��܅��fXn���]r�v#�r��D��Q��0�Q�����Fq�S�}�>T@v �
����;�r*��_��;����L!W��T�����;���X���Õ+W�s�NI��%�L�P(�Z��]�1??�x�<9�	����>�ݻw͋���$c��kY	D�������p����0* _�uKJ��0����`0(;�2J�d����n�saa�4m���ރ�|��k��q3�#��ۘ=�����7�|Ǐ�����###ǥK�\{=E�l޼���Q�L�r��܃�ɛ�]�n�$�Oqyc7�0w��,�H�L�zM�S�<��0\.�pw�Xn��(���y��S�N���v�A��iLφ]���eXn'�+�_[l@�pwS~>W�b��/��U�Y\�Qq}�g�T���$��nR��Z�T�sr�C�ݻ7;:::��i3�V@ ��(�Ă{��Д����� D�(�m�g�W4l?�H�.,ݹ���믿΂���=��^{���(
�7���Ȉ��jll�������\��f�e.N,�v�j��s��*�h��2^|`�ܹsXXX@ss���|�M466ʎ��L&����1<C�utv�
�Ն��s�#z�K�_k%nz�������(��X���YpW@OOzzzp��yܽ{MMM�#��c�=f�cU*,..��Mm8?#Pva(��{%�����P.9��GU��D�)(�7_9'�"��(!����	���6e,�� ���~J�1���¨�]�j�v�zTߖ
���&��&v�P��n�9��$y
ܡi�m0�x��eܮSk��Y��d�@��B�J�S�Z���i�̙3(��#�-�`�e�u���v��ױ{z�Ą�&��Nܙu�ȠG�!�N�h9�E�Z�R��3g$�q����ު�R�`Ϟ=�cxJWWt��)w�a`zz���J��[Z/ �};C�!��`�QD0����M�W�^��Ԕ�D�{����?�q
,/;����:::���f��e2X�l�܁�7ݙ<�	�DDDDDDDD�7
�o:t���É�I�N��`��z��{�e�� �~���wѺA�S!�Z�����������oKJ�O���H�y��Zi��+W�8z�H$bk	�R�X���{�	W,d	�6Ƀ?���z��%�q�{�g�)~�N����-;�gh�����wvv�Bၵ�g�"���wp"���9����Q���zh��#G�������iZ�ݻw��x�E���،�w-�f3=�`�:����������ni:D�}�;I����[�a�өUk��ض�B(�CS�T.��@$�?�� D�Ev
��۷�q�Q��~�	i�m�Ν,�C2�ěo�������B�8�|zz��P�����1�z���Z�7 >�i���[�066&!���ܹ#;�r���dG𔎎�B!���ċ3W&�p����@�׼�)��M믽������f�<ymmm������$	[7��e,..��C-=x��*��x�$""""""""��@��D[����D�h���ϿJ]e���^�ѤN�'_���H!�5�V�������;��K�.YN�&�lڴ�z�"�Z6�5M��C$Ag��GAMNNZ��c��^ˊ�A�AǯSoڏ�������}����ڵkH$�c(evv۶m��34M�ƍm���e�)'�L���_k%!4��&ǯS/�@��`Z���¥K�$$";lݺO=���e��j��~[7N���[n"�t���cӶ]�a�q����������F���\M�N�����2��;�U��^�hR��쩁�~�H�U�T�dD�F�GZ��5�0��+�HJ�_��Î���������폻i�&[KH�\�r�mƻ����IW�So��B(i��:::�\.'!�}�\�";�r���eG���N��a�wrr�T���+��aψ��ZIoH �o�Ԣ���,�3y:��p��a��y�^]���V[���
�+�@�Fq26�=IDDDDDDDDT�����ԩ"�۱c�2 fe�X��q����V!�������i����N���h}�<���W^A�X��ȿ���Q.�e�PZ8��̌m��F�a���@���[������w'b,����h���3�
�7MLL W��O����޽{e���������	���t z���(�T�H�.4=��i���޲,�ZB��;��;w"�N[N���{z{>���Ғi=ҵ������y�$""""""""?R�����5��$S�Wب�0nױ�^�:?4�e ��T*]��a��:��g��i-���������ѣG��dd�PV0ę3gl{�-[��ZB*�J���2A�p.߂B�b۵���A��,�E��_�����/(�A�����4�IX�DB�c'���ӃP(d��޽{����]�t	�m�Oo�=�Λ�^�~�����2^}�U	i�	���A"��ƅtvv�����Ǵ: D�.\����Z�p3�RC���&�`���N���Ph���f�B��X;"9t�� 5�IW�d�h�^4�z´���|��]�i���d�PZKK�\���ǉ�����s�*s�=ܾo���o:�S6�'ܾ�}�0���i[7W�enn�����L����3B��#�����ۦ�Wώ!�uБ�}��[nf�Gk�i�ͧ����(�J�S���p��q @.����H�R�>f�\��i=�ҋ�&�(���x���B1ǯCDDDDDDDD�5
u
�8��1�DeƤ��¡�U�S�j�������feX>�Gmx���&''q��y	i�����;�ׯ_�,��b۶m6%��R�X�5`�܁�y[�W�l�_�~�r���w9�����[�c(%s��Glݺ��������Mfff0wgsA��ŕ��#���_6����attTB"r��i���02�71T�c��O�����|��ك���{��W�o�3ܒ�B"`Zv�UQ��:~:oAD��"e!���TyQ��1E�/�῅`�۴�ba��޽��S�U"��o����������(̇��xc:l뵪�#���+תg��#�m6�loܸ�.HH�6�\�HDv���yɎ����ذ�<����㦵S��{�v�z%4zT��+����_�4�_x:P��D"8~�8�m�ƍ�+�B!����aX~��H#.,6cnq���UÓ���������ȯ�:'$�ѥ"r�*�Z!w�#�a��JH���L�$�P��@���<J�At~��/^��+W�HH�o===�ɵT�B��\.W��e�[��aY����&\�Z��z�pʦ}:>�k����ַ\N�v�����7�t�r�߳B���ϑ�^\\��̃�3��y�olte�N�!	��u�Y0ށ��?oZ�ŋ%$"����cdd�X񺁁������fQ,M뱍����wm�V5Z(
-u�ZDDDDDDDDD�T��"�0�yÐ�۔(� �A�	<�w+u~X*�ʬ�D�����"'C�?m�2Mm��o���Б#G���e�PV,��ӧk���mۆ��4LNNbiiɴ��x=�7f�
�Aod��.�G~��ԋ�W�*Q�,�J,�֤P(pz�Gtww���ɑǾq�i�/~���9r����\��u��o ��v�J�h�v�ލ�Ǐ�\.[�򋶶6�ܹ��ǝ�6��ׂ��{0>���zV�M�W���jt�<r�|O�	� �VÂ��J���'%�?j��uo!����x���ϟ?�)��b1�.;��b�&&&V��'	tttؚ�0ܼy��k��6\���z��I�?Ov�:��ǖ_��7��r�ڍ��"�Ɏ��|>�Fu��tT$��͛y�\.g*n�J%��MXn³��A�w���]H���i��իx���%$"�	!p��A�۷���(�˲#�J�49r��e�l�r�@t�>�|ٝ}��8IDDDDDDDD~'ԙ��F���ABu&K�Wh�w+
���Q���H6U~�"��mx�A�6��9�]�C�aaaAve�={vU���iرc���ܹcYB��xu6�rō��@��m���?D�y�i��իx��$$Z�J���i�kQ*���~�1<c���m��~��i�� �?���V
6:_���Ο����{��$$SSSN�<����͹��������mܙ�a6�W�p�$�E&�X��H�J����B�W��n%��N+%��DNB��d����@CF�lZ?�<.^�(!��i�����1���҂s��=�ۺu+"����.��U���;p�ּ�׫FF��\���h�t|��-��W�W0w6/����FSS��JYXX@K'�@GG�cߋl6k��^,qz:���f�q"���v=������K�p��e	�H���<��S��f���8*�Lb�޽�?���"r9���ho?�on���p����2�]�a�DNR��@�{��Xp��P	U�_B"��{�����O�3�s���_��g��l�ΝH�Ӳc(mjj
�J��ד�$���m����8
�ӓi«s��Mopz�c�Mq�u�N�>-!ѣ�iz�*�
���e���H$��۷;��ccc��������5?��������r��_�*_W�Ծ}����#��cyY�}��u�?��#']LMM�ք���|0����H�+�"""""""""�,Ez����ѥ"r����|�Ƚ�m,�[Qk�Qv "��P�ɈOD��@s;:⟛֯]����Q	�h���(�J�c(+��?���ׂ� v��e�5��"nݺe��lbΏ�SBBC���������� �}�Y��z�~����q�1��N����%;�tB<��c�6�{�畛/
�Τc�Lo8��)�!1�Y���k���[oIHD^p��1���c~~��6;�R)$	�w~~KKK�������vmz{��J"""""""""��?����H��Gsp�%�-�>\+�J�oH��i��2A��K:?�_#��kZ��׿΢�mmm���c(�0d2��Ν;t�����1��eӺ���$*nMool�Pk�r6<�_!�4���i�:uJB�����eGP���U�y�f45�Ow�������"����5?J�8��A�_�@�߶x��g-�+�?���q��Ilذ�.N���Ŏ;l\�00==mZ�BQ�nƵ�ۯiEh:�DDDDDDDDD�2��0xt-�^�RQ�����ͬ�m�(���I����D�U*�����I�D�h�(�?�ۦ��������Ç���d�PV$�*�    IDAT�믿��Zoo/ZZ�n��f199i���>\w���w�v-��B1�|���ڷ��m��̸������ɤ�J���e�@"�@o�yӛ]�ܹ����ֲ�,��w!����u?�j�
�'��ch9�3����I��?����fӦMxꩧ �t?PECC�9��c��i
�3�-Cx�=s��)��6M������������b�3P�.��4MS�[+Թ���w+
�P�|2"�B(�dd(to!j;�����1�?��s�)l�I$A$�Ci��͸y�&�{��-[�8r�+W�X����D\ގ@,-ȟ7�?��h�:dZ/
��׾&!�Y��K����Kv�"�{�1!y�R���ׯ�֟���"6�EG���!K�r-?���ߵ|N��7��l6+!y���>�|>��B;뺎�����[�T*��ݻ�k��8�Ԏ�w~�6op�ZDDDDDDDDD^'��N!�Z�*�v�V:&[�_B"��Rpe�"uMG�Ǵ^(�կ~UB"�ܜ{ӿ덦i�x�"��c�͉�	d2���%mn͸7�4����6���[~itt�ϟw9Ѓ&&&�H��[���9�ݻWv�4M��ݻ���ؘ��z��M\��F��G��C~����m��ԯ�����JHD^
�p��1���!�N�0\�����hmmu�'''Q�8�8�i�=?��5��I� �~$""""""""ԙ�n�]*"'��eu~��&ܭ�G�z�R��D�T*J|Ҫʋ\���C�G|��M�o��&Ν;'!��i���[�*Q����v$	G
��bccc�_�����M�����h�F׮G@���H������/�B�$����C��g_-��cS�U��ׇ�F��#�l�r��{M�>��u?Jh:�Mm�\������ݦ��_~���'�W[[FFF�H$0??/;NU;w�D__�#��������z0эLE�ɻ��%7N}�:S��)$��4M��Np�Ʀ��&�s#��");ê(�y��Ϳ�AFL��~�m�6Nq_#!>���&G6	\�r%��L"��,��{��$�Ɵ�=�馓��x��$$�7��ɒr=�d28p���Rmܸ��G���˗M�g� �������v׮E�i�Ɵ�w�u�0����S�����p��	�J%��y�q��с��!G�R�Xn����=��/O9r]+z�	Z(������������<O��q��d�T*jt
u�-�⧹�J��a8s2�Z��=�)(�ч����i}jj
���7$$���A
�V����c�֭�������ggg1==m��\b^��h��FF�q�������c���|�;�~��ˉ���z�@���,
�z�}[[�l���5n޼�l6��Z�P���9Ķ:z����l��ʵ��Z�w1�_�v/����D�!:���!d2�=0�"�H��'����<�ݻw-_��6�÷/�Q,��!$�t�ZDDDDDDDDDJP���cl��4Mk��a�u�-���'���L�t��OFD��(˻Wp$�S�g�"]�L�N�+W$$򷖖�k�}�v�ݻ���-���{X*������7S�(�YBJtB�v=zP��~��ݦ�J���|�+�����<�aeN\�|>�T*%;�4���ص��|o�|>��7o�ֿ���A���u��hn�Ѓ�]�~Dl���`����7���)��R�z��(�?�m۶!�NK�q��	�B�S[���0;;kZ�"���M�|ǽӜ�H#�h�k�#""""""""RBN���B���.;��T*���N��
ܭT�0y2�w" ��3�������wӺa��?��E	���ȑ#��d����~`M�uܽ{זǿr�
����_�3�������CQ�ـ\�D0�Ϳ�,7ܼy�=��kYΜ9Â���ޝ��q������`%����(Q%J�d;�dK�-;���.I�������4�mӤ���s�$M�:n��v�$�#;��M���ĩ-Y�B-�DJ�/ �}�s�P@�&@$0C����c?��+j0��=i��bY,�:�łm۶e�{}OOe᤟�W��r�M�婳B cu$�R�����#�~���k�� ������l���Qul����"///+ϯ(
���n�j���s�N�U�:!�B!�B!��U���*h#KEHi&[��^��E(���W3ATz3"��ѣGM ���r�)ڹ�%d���;Qr�=>11���zJ@E��`@~~��2r�����}������Vw�799�4(��n�Këz���+��$�߼e�ޟpۯ~�+���d��h4J!�4��a����.C�ٌ��Ȳ��q����wc�~�����q8�c_O_`�e��J�V��Se��{zz��_�Z@ED��n݊���#&�l�a�,��nCQQ�&�LLL$\e�Xր��՛X�3۠3��B!�B!�Bވ{ܢKH�������%�F�)L���M��좋X�$I5�k D$��R+���Qw�qu�ux.�ᙡ����ؼy3ZZZU�>�޽/��"
E���JKKq�m�A��%������f[��B!\�r%�6�������!D2Z ����,�����ӿD�=��q�9������<,K��?y�dV�-
�Z���P��hDKKK�;�{<,z��g��&��L�A.���5Nқ����������O~�455���JPuDK$I��7��ǃ'N ???++Q�t:�v�m(//��s������r-z\қ0��g/�fm�DԽ�aB�(��ğc�%�`�pBV&���=�c�8g`�&z�ՋqI�c��C��$8�20�{���G$kY(��U�&��隘dL8CX��u���	${�v�?,�U�]!i"W����(����i��s^/�BD��t��kH�vV� $!�� ���;z�|7p]g`�9�����������de6mڄ���y����\���h���4JK�[�s��/"�.��z�&\�Ww����BH�D�+B�G]t� �Ӊ#G���@V�V�@ 6�����(�b�Ν��P��`@KK�FcVǉ�b�t�Ң�qppguې_�^�Y_`����\`�x#�}��}��H?�0>���A���2$5���8x� FFF��ݝ�.�$a���p8{�7
��K�Mn�O�����貥 �Q���=]���]VZ�|}~ ���8{��XL��m��()6���d5b�绯����>��d����ђ�d�8��suS3�W�&�N�JG9�:����22@�@���2��(���H�0Y����R7E�Ӓ;
�t[���,�r(�Nַ����IQ*�Q�x�	����[�sm��f[���`�a��Ȣ�=}�Ѭ�)��ʰg���Q� jjj��h�����q��܍8����k?���Ӄ�����7�t�<�,��I�W��0�o�X�mǏ��/���q;;;Q__���55��S*���PR����2�d2aǎ0��Y�����D"��ѳ�o}k�Ǐc:�-{ݗI�j��%�*�=>::�_��Y�h4������h�ARPUU�C��h4�����dYƁ�����(��,2���̀n(k�'������p�n���1x�� +��8uVL� �<�����aLV(����uUH� A/&��p�Ɡ�z����� �`t|���ʉ
���O�"��*dm���u�	�����>��-eE�]!�=zTP-��T(:���>%'���V���z�扬[��z�5���]!Q���hZ�������geL����<������XZ��ގPH��K����8x�`��v ������Ly�Ӊ����t����i�u��5k�3ٺT���\�=�#G�``` �c��v�y睰�l��[PWW��1��9��l�2�٬Z�}||<�9��'����O �^��PXI��s�d�C��&/~�~���q�����]PP�]�v!??uuuhh�̼i���۷㦛n���C8����z=n��vTTTd������^�K�<�ț�54����H��@2XT�">�G!w�R��Nh�=�B�d�D���(�NVj>�>��}�l��;Y9��鰰p{���j���Q�]%�i����&�Vaaa5 Yt)�i&��:�����]B:6�.�Q4��ݩ��
!II�<4|�{`:��m?�����Օ��v�؁���C��,���6�-�ci��fK��q�������!��>��t���q�b���8m�Ќ�_���bH&��c��Iz6|�{	Û�h����3�a $I��f������x�N�[n����c-r:���}^^v��	�ј��|>�\����ӧO��qd�z]�%�r~�j��Y�w���n��s<��#������555hii�^���luu5�+��^����c۶mp��i�4e4q��!���e�B`ffn�;��p�^�Ꜻ��$��׭��X����(�N�u-��-<�G!w�.%G��qr'�c9n���;I��tW�.��(���J�J�=�B��ǝ�6�X%�d��4EQ4���XVYU��8	>5!����t��m!	Yc-�kHw�����IB���t����W?�p��Hؽ{w� �N�CKKJK)���7�	���ѹi�&�z���tI���1����Յh4�p����EV4�J1&�PD!�\g�ߍ����fff���~wՓT�f3Z[[�c����};}dH���^t	�),,�Ν;�z�%����kѱ�r��L�����^��%5�v�'�q��Ӱm�c��~����7�d��U�elݺ���`	����J477C��V�Zb��p��A�����r-�~~>��.��dw���K����v'��UT_H_T�p3!${���
��Qȝ�*���qr'��n�˙p{��I�.�M�L�=�B�$u�n���;IG����(�e?��"U�!Y�8�� 4�UV}2N�Ok��΋�����5�$����Y�wEmo[����÷���U��Ǣ�o$I�lق���U��u�$e��d.b�aǎػwo Z:�Fc������&�����V�T�y�/t$�NrO�}����'�v��9���?_�s�����]�chmm�M7�D�����΢��It����ؾ}��'��s����E+c�b1|��a��cY��z��:S��c�41	>�=ȶ��2���x���W=��b�Ν;�-���aǎ�L!�jhh���9O`*--��Ç����sF(���H�m��*u902��d����\�1	Y��^�s]�n���;YN����(�N�����YY/�(�N�����8
���1LLs.�G!w�
O 7��qr�.>9.��Tm�p�}�L�+�dj�Ԍ[m��8	�AQ��k D�˵�,��T�Y�C�G���qѦ��!<���<��:����hjjJ9�\[[��7�:�e۶m���]�jt:��ۇ;2s����Mx�bjj*q�b��Y�?��:R%��쪎IV�14|�;	ϗ ��s���_N�)���m�6Ȳ������F<x�����
�%�����6mR�=��ի	�$��g��O��'bdc��j��#+�/�@�'��{��/���G����������
�Œ�����عs'�f��$�I�$����n���_0!���w�qL&SVk�F�J�f\1�����ם�d(��&&D-�n���;I&���qr'��z�=�B�$����Qȝ$w-��{���B�4r�y�,�	0������8
�g�����f�E"�f���k{��J,���q�����Yc���Aw�V�,���ɟA2, utt��g�I��,Z[[Wԍ���۷o_�7�mۖ�_.fB^^>���ڌ>��h\d������@��%��nD����v �SIs^?_&X9r�/_N��z=�mۆ�� @ H9��p8p��a�V��r��m�6�ed�N��֭[�5���`ttt��;�+���U�V �vU�du��oA�;��p�O<�s�Υ�|�1466b���i�^`6���ڊ��������}��a�ƍp�\hmm�-�ܒ�U.E���P╮����<?��rԙ��<*!�V��qr'o��p{ܜg3����<����(�Nވ���&���qr'�i#��9������Z	��Q�=;��8WK�*B2�wYZM|�}^p����j	]�-A�N �z�̙�� 	Y�c;Eא*
����R�u��z�m���/q�ر�����$�b׮]��l+~-����׻�/|�v;����EA4 ��n���$ޑI�3oÉQ��Е-��T����v�����ۢ�(��o`lll��Z�hmmEQ��ǀ��L�;wAA��n��ե�g֚���5��G<�[RR�ژN�}}}�������&�j��ta(\]���ݟF�M��qEQ���'�@���`��;PY��I�,c۶mhhhX�s���p8��O~�w���9���n�U���{��JV�x#�%��4JI�텦��qr'qZ�����Pȝ �^�=�B�$��������ΑB��u�
��Qȝ\Ok��8
�g���-s�[E�@��N�<�	@��:RB��%��R4�f���M�8��9�5t>!d%J������9���~�<$�k����lݺ5#]�F#v�؁���j���D��q�1l߾���d��8�,crr~�]]]P��!#W�F�׀�z�M&�(��q%7����p����׾�58�΄�Z[[�"�dYN�Y�q�-����mM��x<ؽ{��2�����v�ZՄ�ty<tww��gE�׋�p��ޫZ-q��zZ�B�>�,��_��`_���177��/((��ݻ36ᱺ�۷o_ѹ��.�Պݻw���6��c�D�L�ctt>_� ����)Č'q�=��E���ٻ�&���Z��[t+F!wr-�~Qs��8
�����(�N�n���;�f�n���;�n���{fi���v�U�d��2�|J;���k	|tXt	�Yt���W^1�%��T�A�%�u�����m���h_���100�h�^�����Q]]��Zcظq#�lٲ��H�z�^te2�p�������e�����IN��j<5V�`D�/u�E�`�A�qIfվ�Q��քۜN'z�!�����$IBSS�������!I+�X�Ö-[p�]w!??EϡE�aſ�\&I��ܜ�	c�
�p�¢�K4�#?}�C�<�B�_
�i��k�d0c�'��|Ѷ��i<���Α�s8hii���PQQv�ލ����>/���
���0��1�P^^���2D"�EvVc||<��}a�zpyܝ��R%���쪏K�z��p{��ׯ����]�$�(�~i=�G!��������f��qr_Ϯ�ۯ\�f�=�B��'��y�K���8
�g]B�8�mG��.d��Et)�VFYut�>�/��tP���+z�� �H��}�Ӣ� $����xy�,���Calll�1�Պ]�v���0k%���b���Y#�ݻw��ZQSS���������F144�P(�xk9�����V����y�痩>.�&���!�qo�ͣ����7��P(4�*���X�_,�HP�����s���W�\�������]t�D�ֹ2.
����D"�����[>	�7�Z���U�:&�<cY���H�ūG���������N�ӡ��9�D������qcc㚜$�l߾6lHz��t:TTT //����&&&�r��e��Yi+:�fW=�JK�T��D�z�V��qr_BN����p{��ן�n�������O����r_��F�=�B��S<ܾVP�=3��8H܈%�Vk��"QcL3YZE[e��U��`��ұ�W^)]!*���`���o��2�`��?��E�v^�>� fffPYY��kb��F������a݄�c��3M����oĭ�ު�q\&�Ky����F����߳�1����`Aӧ����&����^<��shmmM ��,    IDAT�]}jj*c��eYF{{;��߯�kNEQ`0hc�d*c���Ekk+�fu��H�ϟG0\��gO=�������w�Jj�t�k���*��������===x�G�(
,Z[[QV��$���J�ܹ�E��Hf������EEE)�o�XPYY	�N�����fg�יl��m7^�Q�s; ��	'�B2kn����(�~����hd��5$r��Z�`M����!���;Ȓ����p{\,���$"��X�8����qr__�~iM����C�t9�r�C]E:4��"d�:::J4��#Uk­:��w	|t�FY�&f4o�sх���A�5����.�U����3����ކ�wf�6�ߏ��ITWWg��f2���())Aoo/�n1A5m޼/��B�!�\RSS�={��[6�n��Q#�L�n }��A��*�>}a���i\������c��s��^\�t	۶m[4A�gi�\mm-�v;:::�ק�	��
��hk[;*�����Ԅ�<���HgϞ�߿�;�ї~����aq��H�B����I���Ծ�kx����>}���o��|���m�&bxx���:>I��h�ƍQ\���EEE(,,���$ �<�l||N�3�6&�0[֎����,k-�0$��Lɬ���y� l�KɊ�I���2H��?=E1X{�#f]�3��H4���!p���?���cx�;�9YfX��p4�yD�A����,��1 �c>�|����c|p$EY����T ss��n5�`�Q3�# ���� D����kc�6�����.#�i"�-L,
>:V� ���p����:��ٙ�D43��fZ���\����\��CP�^ @yy9>򑏠��gϞEKKL&��u��رc&''q��D�kcy�dv�܉�W���Z)�ɄݻwcÆ���'�B �ބW#�pfBLxM2Z�/�26�>K�N4�����ǻ���0�Lx��އ]�v \.����u���������6���曱q�F?~sss��!����Z���X5I�PWW���*�'�K��O���+J�{U���dJkU�d_���#<3����4��$Ix��ކ}������ؼy������P^^�˗/��r�:>Y�����V��	cv��HSSS���I�7�9��ǓL�ϱ?�!S�ڒ1ci=���!�����S؅hW4���g����%^M�����ϙD�\n\�Y_���#b_m�R�K��m�����_����.C�#��]EN�o3��j�k��Z�}B�j���C ���H��z��x�>�$�	;v��g?�YTWW �� Ξ=�4P�m���hoo��n2�Z������{I��e���-oQ=ܮ(
�����L6�$oƱq1�͌I0�5 B�D=������'Q�Ј��������������Ů}����6��v���o����W-����Ut�VVV���v!+� K���tv⿦�n�C�� �XZ���d_���} `���O}
�cSSS�t�R�V�X��lFKK���`0��@��lhmmESSSF߿�z=*++a�X���9���ؒ��;񣋀?$f�����I���!�B!�Bn�_t�0q�o]!����읢�He
�G�eh� �����&�B��1v��R�9����*ƶ� �������b�,�
�p��9al�^�M�6a׮]�����r p�7&"���j�{�hkkS=�(
�����~�N�9�/���Jk!��]逈a�ߍ�w�'��r��C����	�ʲ���V�w�}������ۍ���e���j�Ν;����Q�<�P(���΄�̮�.�b�[�[T�m��Y
��MT����_Qz��a2�PVV�`���zzz��܁k���P$�n��`4�y�f�ܹ���Y'//o~�H$�Z�}ttn�;��mǑ+&x���ն��
}�C�؄B!�B!��5|�xO:]�1�t�&d�N�8�@��:RŇ(S���m��%�%��͢ $�~7�J3]|t�n���l�(��a�فKE��ȑ��q��x<^s}h�l6�#[L&SN��JJJp����n2� �appp�p{�q���!궄l)�l�n ���s�����X�V���!I��unnN�� �Պ}���;�X,�u�slٲEt+b2�rb2���Gggg�c���?�e(��*$�	��*!cuE�3(���U��_�*fggl���DWWET!�����Ѐ��6͝+�L�e��ա����媍[RR�ݎH$���a���%�7V��`�V���1&�XZO�B!�B!��!��&FE���d�Y)�N���,�rQt	9����W{���e�WB���]!���ѱ@��:R�\� �B�P�~G�\y���w���Y�o4Źs��t:�.s���2���c˖-9_���v�\.�e  
�o�>�u�]���RC4���`Ґ0�d\2l�JP��%� C�f���
�h��K�x���,iǑ��H���###�Bj��@yy9>��o�]3�gggQ]]-����������nZ���Aggg�c���O\�v�{T0�`,� 0����q�ɫM ����@�b7��`zzz������]�d2���܌��6���
�e-��t���ƞ={P[[�N�UwE����^o�}"e[qd�NoP��2�ց�Ŭ B!�B!�B�Z��%��tl|��ZEAH6q��@t���+=���y�-�r�a��>�U��s�����Qt�dc��kH����,!��Bp�"����w����x��/�3�X]]]���R�̤JKK��ֆ��&�L&��dL}}=��%Ҋ���o�>�s�=����=2�``` �`����ɛ�_2A�v��e`:Y��D���݈�|����o�O���&h��a$]�@�뮻p�m��|н��At	)3�ذa��݋��jH�؏�3338{�,�	&}��p�_�o�c�]c(��dX[���BJ$��H7���&B2	տ� "Umx��urw��8{�,�a1���g�X�e��ڵ+�ϕZr}�����,�)
���n�;�>��mx�� �s꯾'[K [���O!�B!�B�Z�{�E��I��Pt�d����7��$���@��w�upO�;0Sw�&q���]G:(�N�� 4Տ��`� �u�-�~���#Pe�6EQp��E����X������n��D��j���K�o������~;���7��BH���Io�ވ�/MX n* �/��d�
��d[�5��x/x,�JQ�E;��|C���X,���A!��8����q��w�;�@uu���x"���hjj]Ʋ���y�f�ٳUUU� 0::����E�� p��)��τ��)��kdk1d[���I����k�&#	&�I2����x_��W011�`���ř3g��-�D$��j�֭[����Ñ�q-2hhh�7܀����za�ď��&�y��ᱫ�p��M��fKk��O!�B!�B�Z��L�;~��"d���t�j��hka�-d
xOp��D���?�%�E�iob�Չ�#es.��1�U�
#8yJh�n�֦7aX'��?�����ۇ���y�f���JKKQZZ���9���`vv6a�O���p��Ŭ��dYF]]���QTT�ձR���0<<���N2Yq,�������-��؅�@��+1�����R�ҺG�z�?*&a�[ܥ�s���Q��a������v��v��͡���������s��!���c(..Fee%
E�3�s����E��cǎ�O
�ޣre�������&�q�!�Z�cp��iL��򗿌O|�Vl�w�nnnFqqnt�6��hjjB}}=���066���s��fCEE���rb"���zzz�&`΂m�I�!q�L��T�0�PA!�B!�BH6��a�3�k�aކӧO��]!Y��
48AF
����^]B�v�:uj��ݻ�U@��ػDא�iE֋�ߍ�T�K���m�O^1����G����X,�OOO#b�֭0��.yEl6l6"�&&&011�d��\TXX�H$���{II	6n܈��z�5���tbbb"��0X���	�fĆ�%�	��z�5��Q"A�&�$�D��m~4��|�E�o�MOO#���p��l6�p�hkk��� ._����)!���n8p@��K1�Lp8���&y����ݍ����۟{�(N�� �*W�:
l�m<Eh��@�cp�P~ǟ`�Z���5|������2�9��������R��������EMM�N'���1;;��Ze�e��娨�X�YA���~%��$����>���+���X� �ύ�R�B!�B!��I�C�|Ү��+I��(���s�������H���5�I��)����10{��RR��>�S�� $S:::, �p��Vd����Yџ5�7"z�����~�=�:kz�^�:u*����I��ը��������055���Sq�7��W_��j�����塮����9�5�s���)���$�'f*�ӮF����&�`�7�I:�����zg� �+�D,ڄ��pO�j�
��r��FQYY	�N�q$�2����ۍ��>���V��f���e���(++˩n�׋w�O�MZQ<��_����ֵ
��u�\�����D�h�͋oz'$����/����t�M��8�z�*�^/�����t��J������וj�+s�$I(..Fii)JJJr��*���ŋ���M��d0�~���Ҙ����J�,��!�B!�B!��/] 4p�G��Ձ���EH�Pt������V}_�(��"~����=z���fD֐? ��i�$x�I�%�5<Ex�Q�{U�#�A�����-�{g;���l�F�8�<�����а���!��}Æp���a�\� [y�&//555���Ciii�H���0<<�d�}��O��c�'�s; ��!�M�� ��9³È�M����;��Xq��1l�N|I��z��ߏ���Y� 


��ڊ��V���`pp���Ypz<�߿?kϟ
Y�QRR2j��se������v�����O�޶��\T)���Q`s��M!<;��慻�cI~x�/033�{�w����Ix�^lݺf�y�%g��`@UU���1==���)x�^ѥe�$I(,,DYYJJJrb��y�^\�x�@ �>�)�D6�a�}�eK�ڹ�I!�B!�B��)�NC����.#%V��� ~$�B2��ѣ& �]G:���)L�S;���7�.#%V��m ��.����L+�΀������P�~�&�B��2�|����{����e��2��{�n�����͛���32n&1�PXX���B455�����tbvv�gUa�lhmm�/��rg|I�`��QQQ���*�v�0`ddd����z<5a�\@�dCqtM��")�B�Wf.�����]/�������a������"'_�%%%())��]�077���Q���bbbbUo�H����������"�j��t� "�zzz�v$v�\����v�_Bo�W����"
l�E\AhzQo��V�a�݉�>�g�g�>��׎~�gΜ��M�PRR��1��d2ͯ�D0;;��	�Ӊh4*��U3��(..FQQ


r�S���������ĄȼR<�݈�)�ו��CY�M&�B!�B!d��W��3`E�{���c��a��~�s�Z�%G(��K�
����,x$����dc��p�ԩ����,��t�μ&�B�"�Exz �g��l@�}�_��F�z
o��EA�Ӊ�'O���)�I `�Za�ZQSS�h4������ǳt@F%�6m���D�@�^�Gii)����dY��������L:���d\b��p�Q�!$}~)��e�S�^'���2�qI��%wa��(޲�C��'�s���"�n��l�:�
Fss3b����199���)LMM�x5�@ �p�T�I���:����l99	+�˅K�.!'�~��e<qzyw|�ľ�y0����d���M
�2����4|���t��/}	���Q\\<�=����ذaCN���k�ev�v��s�|>����k�d��\b�XPPP �͆����Ze$�h4���^LOO/�_ �
O��a̝�ɿ��tz������O!�B!�BȚ�9������ѕ��'Nl޳g�%х�Z����!-�0x�9�Uh�6�J9���.�mo]J:n;q���={�PҖh��(���ɬ$x'-%B���Fdn2����C\܌��}���/
�D"M� @�e��8��z���|~���Y[[���^8���p�s5�L,���(��%�e����gf�?�@g·��Vt$â�i�g��rc�8��z�V�$���	ws:���������0�N��p�Εn�N�.�k��~���F�0�O�eX,�����X�VM����(���p�}����i���w�XYb���}#����&���n����cٹ�љm���0��C��/~�Ї��Դ`���1��n477#///+udcl~"eUU  
������������!�O����J�L��s�\���A(�Dh]�a�؈�+�?��v&�do�3��G!�B!�BY?{�V��1����DB�j�:u�]Q�}��H��}�@�\��o��'m���$�w��������,�D"�]GZbQ(]gEWAH�d��f2�ڝ�}���/�=o���Ջ����DSS
U�+Sc���G~~���#������p8�h4�H$�H$�v^��C�����L&�F�L&�L&������@��v�G�׋���%?Ac~�È'���4H3�區�&�%p��~D}NՆt�6�qwxNase�sa(B?�v��Η�1.�9������'	�B!�B!x�^����5�N��^���1�Η�̋��x��ӓt�@$�cO>�����єp51���	LG�.֒�ka�h��d8��4��m��o��� ������~�9suuu�����? 0�0�(--�LQ�Eו�Ph�5e$Ik2�N�������ϑן+��;�S}}}]����y8i�+C&(���c0�o�d��DB!�B!�B�~�4�� m����cǎ}��o�]!+����־�����o�Ӡtv@���E���?����l{{���BY�h4�� L��H�r��&$�bAB�W��]39�����8Xu��z�}�� Ν;�Á6h>�
�1�~=�9b� ̇�Ecl�'�{H�S���Ye���b1LNN��r%�I�a�P���,�'(>� L��ɾL[78��H�ɫP��w���ll�ν�;��$<*����1x<8��z������`U�7
�B����?G�b1p������H�N��0f�EA?FGG�Z�����K����0��*W�cL�`��^}���+1�����U׺�V��̑��ҥK����a�X��C����شiӂmZ菉��%~�T���?/��#%I���p�����]��}�\�������ܘ8i(���R �B!�B!�B�-��_��i��R�a������BY�ӧO��b��]G�
��em;�a|d|bLt�|Rt��Dggg�����H�r�5�%��8B㽪��������|���G��M���q��I��̨\��c�ey���d��b��l��6ߞ���r�5�����C__���vC�+[����	�K:�M`���M��߅��E!��8�3���n��%�s�'�y�^\�zN�z]���9GII	 ̟�]��f3,���3�}=��gggq��I���$��r�5<r�݁�)'��������d� 8ڭz�=N_\��?�Sx�\�xq�>��O����PZ�͵,ޕ=�r��dB^^����WZ���h4���^�={v�p�$a�P�Nm�]�=7��me�� �B!�B!d�SN]B�8��W�΄�    IDAT̢� d%b�؟Ac�������24e�~C�%��E��9v�]t��+@��:��9��ߊ���U��0"�X�n�g����/��ի	�	�B���¹s����U�P�c0���5�btt����D����r1wműI#�1��u#v4A2h��M������JLt%  W�n<>��G��̠(
���1<<��kH���0L&M-��U�p�.]�������/[�zû ���u��D�A2(��		���T���a��|㻏�駟��Z_��ԩSp�ń�z���p��I���/��1�F���#�p�M�M@o+���Jt�B!�B!� �c/9��HS��h���"I�k��� �!�u�Ky�עKМ���ZC�c���ɲ���� $.\�2��\t��=]�3S�� d՘l��eZ҉. ��+������O�|�h�`�����ӧ100�X,7�ZPTT�PHl�l9�s8�N\�re���d�C�~�lĸWI����`tl�d�]
ɤ��}Æ�(ߊ��rx��;�z<\�z33391�i�8�(,,]FNP���������d������/�u�����Ѥb�K3��B�jk�+Y�����@t  릛Q����W<�������E���~�={.\��k$�>�χ�g���ŋˮd4g(���f�6�;�&@���PR#�B!�B!�BH��x�e�U��s��������� $�$}�Et��h�X(
���\]�J|�رcբ� $U�@�S �Eב���5D2X`�ؔ3!w0۞?@���+��/'�p��8q���k"�������]�|>���c|||Q�����xʳύX��R���X�:�X��NSŦ�
��1��ё��]܌S������G �<��pyy4�dzz'O�\r�W0ď��(��m�y�� �^�*�3WA���.�dc0�7�L�]���]_E�Ə���/x��'^c����ԩS^��hC$��˗q����;����m���rj�$ ȖBK�D�A!�B!�By��߈.a%�L&��EAH�N�:U	����H]��P�}��~+���0�t��]!����( �)�u�MQ�O�"�
B2J2Xr��; �*a����J���)D"���E"\�r�N���̌�Uj��lN��%``` ����I�cF+��M��D��r+������	���`:��:�E��@��/����]Qx��_C�`���Z��m��Z��K��t�������^�|y��<��%���)L��*V�<Ca��e�l�O�2�΄/��C������9����=�����F��ׇ�������@�\,���0:::066�̿!ÌΎ#��xi�(�&M��l��|���R!�B!�B!o;�@�����رc6�E��X,� �Eב.啗D��Ip_�.������7�����o E��H�t�I!Z��H�<�`,�.�m׽��I<����ܹsIw������©S�0==�b��c���FE��`0���a������'ߑI�5V�q�<?��`$�H�p�l-]
Q�0ٛ �ѥ,��Ko�g��>����^/�^������ݿsQ(BA���D277��g������z�I�s�\x�g/�y�o� X���B�E��� j`L��ЙrgR�\�@�{���S���O�ӄ�}B�z{{q��8�N��tq�1::������-{�������M�`[ו��p���H�v�Y;�s�k�^B��7\(���gB�J�ܨ/q����pcw�%�BV�*D���DG�ʪD����=BR��;�ˬ�	3�P._��8�W���>#�B�s���-�����c%4�T[�J�i��rI��"�B�r���& *����it�!�Й�s/�@���p�/�L�����%;��|>tww������=	�NI�o044���>x<�%��
��6<6R�1O��Lc��P�@��u��096�^�@�P�W���eN$?r�1;;�˗/cbb"'&�,�l���Us:����Dgg'���7dc�����o���{�_\���cE�0U�.���I0�X� ���Q���ߎ/<���ёp?�׋��ϣ�����9�s���1ttt�ʕ+ˮN�tz���3�p�[Eɽ �l)�ɾȱ�c���1��{f�(�N4G�9���N���GQ,�V�#$�=�����g���B�D�Zs�}����>�F��2��g�&�,���kb�1y�(�����?;#�܉��8��F�J�((����Qe�Lc�}������ d)��� ��:������.C��[�R^z^t	+����ɓw����d���W�^*l9�0���]!Y�3�`����E������}�o����~�+D"ɿl�z����BGGFGG��f����/�$�9<��߿db �ތs�|wr3N��� c����4�	� �7�T���$���ܥ��$?�g�*����E���,�\����ɜ���a���$�sLOO����8�<�������x�\��~�w�%'C���j�+D�A`�&GdKn������|?|�$���	ccc	������{���b�k���˗/#.�'fY~�nƯ\5p�r� dk�	JԹ��Ma
�m���7�| ��X���;єÞI��6����r'���;\���� �e�B�D[*#A|`v�ڊ��~�>7N!w�y�(>8;{4 ���>
���۷�n��I��>
�D^!��dY���"I����Ƙ&s����]�f�W6���y%��������� � v���k�ݔ�]�N��]Q�Dױ��/"��]�&}��_�����.��A	���/�b�9�S?�͕{��-ۑ\�ף���k�}=��n���2!���r��t�4�R��O�|�{ӌI:�Й�E��Qs��B���<c��]FB<Ep�J(w�46F�h����*��ғ�c��l())��hT���q�QVV&����D"������(B�в���{0��{0��^��8ci��R�ed���qD�D����y_΅� �#4Շh��|W^����m���w�󓿿��fTVV��p]g=�D"���h�װf�o=\#�K����`(�]IÍ�|�����y��<�Gq"4q��7�ۯ����pI�:��Dr����녙��נ�`P!��>�~=�6�S����n��	K!��9�隘�7�ۯ7`�����r��
!q"��q�|�M�U78������:�^GG��9 �Eג�H�O�𩳊�Z������EhR8����Nt%+Q��o��o��.�����^c0� M�\b?�6����24�Lӝ��!����C�"p�'�)'��7B�mǀT��W^�94�ݞtEQ�v�1::
���^�)7;/��d2��tB^&�.�9� ���166�׻|}I���c����*����9�N-]��Y:{HB������l�Ϋ�0���q3�{�oxqDF�%0�EGD@ň�(�
DEI��$	��d�}����<��:����z�9u�+WX���tw��<G���r<ۓĨ���p�K��Rt٣�!}x��Y稞qJB�I6�ˎB:�{*�T����"��~�E��+��Xu�(3�͢���t���4M�o�ض����Jidd����+�����~��?�����ǿ~�8+���ƷO�B ڼ tq; �}ݾ���l���'K�����N��f6�A�ڿđ1?y�K�=r�/>�M��㠿�G���yH$�u]���1<<��{�b׮]�ԓ�l-�-CM���R�����,��܃���'��M�kcnn/�k���s9
�3�� ����X52?ޓ?�.n �e���L`�7j�O�.n `Yv���n3^�qD�p�� ���x~M�]�Kg���ε�07�����5L>�2n �G������oϐ����W��N�� T�����;�;��{�W�6�B���b�>2=
=�� ��UW]����۟ǤQŹ��+op���!w����T�,��$tFU}��t�Q=甴X�ہW���٧Qɡ���?^J�t:�cǎ����p]�X��wP���L&S�p��>|}}}�d2�g{������ez1~�߄�̌g��f����-Γ��O�x�)sc�쳟��������y4m�(f՝9��mCCC���G.�C$Qr��R��4� �mG������`dd��ˁ����xrh2+/�Q7�Lk�Nіž��g�����Z ^Ƈ�W�h�"Ԯ�x�(��x/�F��x��S��bpp�������㡽��\�űcǰk�.8p ���~��Z�P~:z�g�����v�o�0�稞A���}���_�-n/`�N~v�����;�ٙ��F��gg����_�-n/`�N~�<n �����C$�>V��8��w��+�C� `۶mK������w<4w���e��~G�τ@���!Zg�^2]�֮]�GB� �:;;W	!R L�[������>�=�3����g�}�{TϠi�����p�#���]h8�޲�+V,��ϫ��Ass3���OyZg�>|x��ι\CCCB6;��Whz�l��W�_��Y�E��.��C;~
ϵU�x!jW���g'%�=����e��݋��>�7'y��'��b���AMMMY���㠹�9�#�����>;v���g�h\?~����]u��_��7��A�m	43�7��[`W=㔒��
#Q�z�YكG��;�z�y�Q�m�.��[/� �\r	���N,C[[ZZZ��c鍤���c����3���r0��K�X�1ޗ{!̦0���1����_ƻ�Z�zF��2��͆v�>�\�*�d������m����&@�2��}���pC;���k5
����I �ִaKHo����l�>Qg��ԴA�sb�����7���Y1���J�q��-���]�z�te5M[�f͚U��&�]]]?�R���-�!������|��ވ���� �����~�#�rI)����g����2-���+!T/	,�!�p����?Ǻk/8�����hnnFSSL3���L��y8z��bU)%��,���122�LfjG�=��*lw`߰��y��A�eD�Okc�^��1�z��1i��W��y	��s
�z<Guu5���Kv��m�f����q���Eoo/\w�oxuwwc�+ǰ'q>b��>l ͌�o2�����{q��Ad���J89l�1F;��u+��.��S%��$Z[[+��ɩ9�t�\.7��;�E`$�\���)�@�e�X Ou�qܧ��;��t���^�Ľ��1�W�S �?��0r'��j�^�ȝ�b:q{#w��������� j�`���@p�V|n�ڵoB��1�T1:;;�Eq����|�k�~�Csg�����:D������/NiC�bY�G |J����~�	Ν�U=#����=p���TϘ4wl�]?���\�zՔ#̚�444����d"�/:?~���n�l�t�t���S
4O0�xa0�v;�g��Gj�a6�".�)����#w|��kA��q���X�TŦ�u�i����B2�D"���MEg�.���i����������>��`�/��Y�};��%%ZY|z�іš�`�^L^.�����E�J�6�?�Ѯ�������K���v֟&�@MM��؈X,V����y��Ӄ���)G� p,A�p�bܠ�1	@�Dm]-�_A��}���J3����jӍ���jӍ�$�ն�#wRc&q{#wRi&q{#wR�wq�8��@���K����PGG��#�2uuu��<o���5Q.��T�$����/WC���g��3{���+�șV�e��,���h��}�U�4���p�{�f,rw���L�D`�0PWW���:���"��A��݈F���r�����4l{������1��.� �A9Vs�a."���g���������O�Ds�0w�y\P3��������bH$'�M'x�f��3gΔ^�e2app����f���@:�Ƴ�^��c�-�cɆ,-#وh����`�^lҵ�=��B�rۿ}[��Y�!�����k�N�:�H$��Ѐ��z���冠 ��� ���?�&]�x�W�eo>ˆi�0��d�F ����}f^�&�@�\F�TV��x��!,ˌ���ի���q��`݌K�7Ӹ���;�2Ӹ���;�R�����;�P�����;��׸ ��%����g�D��.����Pe�Rj�T�) oW�e�ܟ?��;U�<���6�mw�~��?;::{�6ώ;�l۶ ,W�e���m�?�	�3��{�5� �� �>�7Տaͪ���6kjjjPSS�d2�d2�������FFF��ߏ��8�3�����~/z���&�C5O��h���g��{�I'�̱��i�S��6}�����5��9� /�"�!�#�!��1�R����w'{����cdd����
�^z�eX���]u.�����BD�"RӢzJY1p/�!{|��~�K����@��ὺ	�.����644L�M�P]]}"vO&�����o����uJ{����C5أ/FF3��'U
�3�ȝʩ�q{A�n�^F�TFŊ��S�+n/`�N�V̸���;�S1��F�TN~��"��Ċ�TϘ�s�\��_<�zU˲�p����y�?򯐯R�$�����醷�ښ7�^2뻺��\�f��zU۶?� �� �>���	D��E����c{u�& D�a�q6�6��R�����f˖,��)��㠯�}}}'��i�H&����B<?�Mu�����FGG��d������L�d��i�H6@���-�@�yD$�z
��0L�g-C�g?������L�c�a���m�%�cǹs�`S�3��"��bp��G���h4�H$�h4z�a��rJ�v)%2�����tR���Çc۫�a��g�;`�m@�H��I��ZA�%UO�0�-���=pxƿ���H6���o����[~Mc���M+�n�:TUU���{������F!���P]]���jTUUM�)�466���Q���bxx���3�ar4�ag��n1=z���v Bh0���HN��(Da�$;��?�ȝJ�q; 4�9��� #w*�b�� `JW�d�NeQ� �w F�Tr���`]z  �Sɕ"n���4��w��;�\�v p�>�`��F"�� \�zU�T*u����;f���¸�Hx�{�����Ӫg��~ =��P�Y��� T�c&���?�o@@?�	�!&%r}�`S�dF���8ԉ��!�?'��ڋ��7�X�i���r��H$�0�iڤO�t]RJ8�۶O�����f��d��df���N�xi�
������║lD�iP�/����r��#�w00���h#�17���X�Z]��p����'����p��D"�|��u�7\3�ˉ��ӱcǰm�k�m7`�u-��yE�g��ǒ��,��А�'����F���@>% ����˿��?��kWc͚5�F�w��X줛'c�؉�a���8�d2;�}� �-���Y/�H�*g��l��`>�&����1%��^<<ɝJ�Tq�D<ɝJ�q�D<ɝJ�q�D<ɝJ�Tq�D<ɝJ�Tq�D<ɝJ)(q; @D>u'��`�$��_k׮���n�7on0M��P����o�r�K�g��"��� �d��3"�xr��ݗ]q���J�*Z*�:_J�,�@�*�ܵ�3O��
���M {|d	_�+ig��f;��(�ƊEsa�fY7h�v�hTJY��h�\a`߀���:t��1�ǋUB��0j�UOQ��{�y�4�����K�br9E��h݅��~,oK"YU�O�t]���i�?�}���u]x�W�k��yسw/^9��~��ͫ	��W�    IDATx�^�i��0��7����t��S�J�����Ȯ���ތV�V,Y�իW����(�|M��D`��I��]�O�v*?�t�ķ@�\��M��W���L��т�E�B�F��A�y!�·j���z5��7��©��/����0r�R)u�^�ȝJ��q{#w*�r���ܩ��0r�RT�>N��2������1S�Rʋ֭[�S�
')��J��g��̄��
�>�zFh0p/"m�[`���T�(�[:::�����>��Y ��2��8�k�����J���2H;���=�i�S�GJ��w�9��c�XҜ����i�4B3�g�x�8$�qT��.Mߤ��"ڼZ�J������\��3�ڰ��!4����HV{ho�-���~688�v���tG#�s.��V=�h���l���o3p/)�x���K��s1��#/?���,nN`�ʕX�tiYObW-��a��Q��$q؜���,Փ�J�H�,Dj�*�F�J�����S1�3n/`�N�V�����;[���F�Tl���S1�3n/`�N�ĸ � ��^���r��+ .���T=��ǲ�O���3e�~3d��3B���gm�ܷb�b�Sf��euutt<�z��ƍ�l6�-!D��v �y�q;��H�Yː�;���kʄ��r�p� lsr�o_A]�fiCX�``����D���ql�Ł���h�@t�2~@�n�4���6��b���tD[C<
��R��7��ՠ?v��  �E��n���I����eF�H)��ۋ��=��DqI.Bdޥ �S��\z�ѦF8��Q@�~�hٞ}�n��6�tT-\����  ݣ�x��o�y�ɑ�h�X�d	�/_�������?��it�U8.1X��%���e�Ǜ&�ffIv����;͘�� ����{��;E��v 0��+�2r��(w� �;�7H3r��R����Q��L���`~.���d�N3ظ lޣ�����^2S�H)�R��"d�ߑJ����#�w̔�g䶭�g�
Op/2m͛a|(���	!.]�v�s��P8�R�/J)�V�c��񣰯���{���������Ӡ�M�Cm�u^��4��f�4�>�]�#�6�e����M��`{��'�Op/?/�F��>x�1�SJNd�Q�>�Z����%<�mi@"��7�]���Ç��3�c}^z�Ȗsa$T�+)!"���'�	<����k#׳N:���8�}�t���ᗑ�A��ZǼy�`���������{zqx0���ze}F+r��
���d#��v-l�8������I�4����x�;͔��}���p_};�E���:����}"��N3�*n��'��L���'�I�4���t��wͭ��̘�sk׮�V�
������~ ��8���K��Pa�^�� �,S=��h�vњ5k��B�fY�u nS����6�{�)�3B��{e���\�8������;|�vj�!$1�:#�:�Ec����:Fy�c;�F���J:Q#�a���#z-�
��'�wE�Dn�58�GCs��dycC��A�ۋw�A�)�PAkK��hYv��������@Fb�10�F1 6�a4/��)���"1D[B��}o��]g���C�
�d.'g��ÿC�g/�c�Q��Q��b@ss3ZZZ��ֆ���,�D?���a �� �/��h+��@�}~ś&+��b�N�ᇸ���;M�긽��;M�긽��;M���F�4~����	��ȝ�(q�8�?��kT�(�ttt|A�
�-[�,�u�Y ���C�z	�Mש�:�K@;-��ܬzF��d��[�?���+�(R��;��? ����n���^����C�� �˧"  �4�� "���0�����DDC��yLC�t]C,j"��U ��� M�'"��W3�����rF5rF�h-22����B?�8�_3�w����=����_|�o�F��l?"��2���"�K�	����]���x,���҃g��z��yFcYR71:�E2�DVD����qdDzm��f���>�i��0�����]-����w,�orL��3��w�<g��� �^gQ�05���i �:�7��qh�뿷mۆm;�(2��2�D�ӑCY=�����W!�'��̂Q��v�Z���x�d�b�^z��i*��0r���K�^�ȝ��/q{#w�*?����i*��0r��S� �4�����Q��< �wtt<�z�eY� ~`��-����1x/�P=#t�sDh��OA���e+UO)��\e]��ёV=��Ų�K���A�v p�&�v�"3������쇓T=G�H�H9 �����:��T���_��5�6΃���4h���bI�看\�!�Ƴ�U�ë�G@@)S^�43�h�|h��?�BL&bm��:��Rz�'����mY�h������v�ߐpO�Ɛ�M��u^+�n�lh��lP=�(ԖdG�O����Y�1n�&7���`�N�ⷸ L����Ӥ�-n��żs�$�-���,�����  ���Y>��E~�Ǹ �Ҹ�� #w:���� �yp~�����%Šx0�J]�v��gT��`ٱcG��8�K)C�˗~˸�D��B�8߹���r� ~�k�.�gI��J�.�(���-� �톷�תg���#��.A�u	4�rHe"4Ѧ���-e�N� 4�������O�( ��Ե!>{�v
�HM�s����E!�x�)�M6n�<���9+��I!r7���;�_���B�^��'���1n/(D��<�NϏq{� ��#xs�0���k�^�.=��<��I��׸���G+�
��P���Ϳ�<�O��bIH)�u��u��Pplڴ)���~(��X�����w�W�"������a�a�thhh�eY<R��*�J�/�|@R��bq����Q)�Z��D�����Q	�֌�&�S��L�%��fc;����O�$b�W�����2��Dy%��f���-E�e��e�#w:������L��0r�3�s�^�ȝ���q{#w:������t�� <�w�^QL5������s��!��eE���F!���R,��_�����������o��T�()� |��;�Igg�*)�����2o˯!_ީzQe��9��^�'�R�i�X>@j]�ǀS�	1��:�k(d��?�O�8qem+o���B�Y7�+�'������%n/`�N������;�J��F�t*A�����J�^P��MF�4.�q�8��Rϩ�QLuB��lݺu��!�_���B�w��R4�,����zE�1p/!�s���W=�خ ��M�6�T!�I�Rk�� ���R4���Y���J3��^�h�<��H3&tfc;�s�e�D�"�����#Q�s(���Ե�	>B��0��+��B�1RȨ���8Q?|i�H5F�T�����;M�����;M�����;M�����;-n/X�K㽌�	���߼��ׂ���=���y��!�?�v����U����G�������0%��p#d�q�3��ϫ����/�a:!�J�UJ�4�P�0�c߃<~T���e�4#>w"um�Gh���T7!>g%"5- On������Y�h�|>�����5d�ρ�t�s�JB3��Z�X�R>���E�&��іE��zM�ȝ��0r' �q{#w��0r' �q{#w
j�^�ȝ*-n y���>�zF��!~�u�֋U!�رcG����� ���-E�����~�;,�J-�����W�������,�V�R/�J]&�|@��ŕ���~���DOh:��9�e����P@�Z�f���4�O�� ������)�&I�&k[�h�>�*��A|���'� :;�Gm������ "�Z��?2r�HA���W� ����p��!��c���A���W������+W���F��������3��VӴ�vuu���!����?_�8�� ���-��|�^ 쏽A����l���N�3J� ~���5_�Rǲ��I) �zK����ዱD~!���н�^��)=�Dl�9��.��T�N�Ծ
��&>��NA���Sg���=�D�#��f$�W�l���Ԅn�l��D�*աzXQh-e�^q��0r�La������;�Ƚ!n/`�^���0r�<a���W�J�� ci8~U��RHz���eYW�B�tvv.��r����;��۹�sϨ�Q����p��`��Eɕ��=�u��u��PyI)Egg�M ���q���g�z���!ڲ�Y�@�	�4���f-��V=�H9�G`6�Gl�
�D'����|*
Q���m�?����O�  ����m��(P�W������+K���F�%Lq{#�������{�[�^�ȽrT|�>�����mU=�L �Y�u����*Lgg�B�� ���Rt�ܯ}	��e�wh��H7�|[��Ri�4m�eY�z���͛�]]]�BܨzKI���|틪W�Y�j�f-C|�2�>[��hbmK���f�mYt"h��I�D�'��9F�A�"�zfc;���!R���+T�)(����a;Q�1r������+C��F�!�q{#��ָ���{��5n/`�~��O���ͨ�Q*�X���M�6�T�����\� ������oB}M����S�������.|ĂŪ��B��[���={�|��+��W���[����=)ehO�w7�����Q�fv�/R=�$���͌K"ֶ^n��Q��}�|;��x"5-����B������a�3���CO�&�i�Q� ������~"�mpFza�dXz�a¨i�Q�̛�B��?P??
���������y�#��P��9n/(D�_kh��H\�*�0���� �$�tİ	{�^�.=  x�vV��V���������v�xA�0n#y�(��> �=�W=�$�﩮�^�e˖����7�U��Jc�ƍ��B\�������'?T=�����Z��l�EKY��B�{  �|¶�����To��,� hQ��T䫿���:�g���z��Z����F�5���A!��=��0��0j[�Ex�w9��)<~BԮ�s�3I���{��ȩDF�Fm+�lQf��n�=t\��SJ.+�6u҃=t��1xNN�*��M@�0��y�E���w?�^��`W4��=D*%n��G7��L%��e5��{�TB�>����6le���Oԙ�c�"��O��L0r��g�i�����+T/)�^ ����3�C���l�Ҩ��� ���-%㹰o�r﫪�T~�/3�g�'�}��2�4;���:To��ظq�nY� �D��vۆs��C�U
͌#ڼ ���a6́f��'�	�@�����`6�g�NTB��l��ļ�m�-�P=�fH��&��D�u	�v�b"����]�X�b��Ջ��D-b��A|�
I>�(�
'��>�*1n^?ɽƇ7���UZ��~�{�=�z
A���@�$��<�����PTb��Or���#�W��W�q;��I�&�Jx������|� �Q���<nY�J)٭��eYo�u�a��x�?¸]^(p7�y �O�X�y޳���7mܸ��w��[��/^��) ��k���� P=���D�"��(:ֶ����M �4���`�ρ�ieD�'4�M��^����T7A��@�"1�sxQ)	=Q�X�R$�B��B7T��)z��6$��M@D��{�Uj�^��=*1n/`���0r�J��֥��\����܃�q��ȃ��>������5�J=��s��U=��OJ�Y�� �0O��R���|gT$�
Hۆ�?�r���!��q��lٲe��14u����k��]J�6�[JM����+U2=^�h���D������M���W��n���f&`6�G�}U�	�}Khz������?�1�%*�¬��D�y�6͇K��D�!����C�u��7LF��g�"�܃����F��V�q{#�`�丽��{�Uz�^��=�*=n/`�\�ۧ�}���^ءzF9\b�N˲�^��:˲�uuu=�� L�{J�rZ__b-���> w���g���t]Ouvv���-49�e5uvv> �x@��=%7<�� ��Ez�Sn�"Q8�=�ȓ�}@FU=b�����#�'`�]�?ս��7��"�V�|$束?�=Z�zQ�Fl�2$殂Y?�7��M�x�E�u1�D- ��=1r"��'c�L��_��=�����{01n?#��a�~2F��ø}<�]���p-�-˺������B@J)R������ ��{!�U=�b��R�}��[�g�K���T*��-[���z��eY�E!�{To)�; �T� �r*D�����&�Z�����`�R6�5km^����mY=Q����g43���y�#>k"�M��zVE�cI���n��-�|GD�����1�\D��xcP�i�����+Ɵl��D�F�܃�q��"�jF��������7b�,��O��{p0n?5F����}�z����+��L�|����[gg�T*�S)�� ԩ�S�ޓ���Q����JR½�`xH����R�M��m�e]�i�&C�zݶm�tvv��F ͪ�������Rϩ�AD*	z�іE����h�|�΀���&D�oB�uI�}�MZ,	s���X��|��x��'��ļ�������f�a��A�����A��<ٽD43�z�>w%"<E��&iiv�a��k��Ϭ����}����Ӌz.�7#w�c�~z�܃�q��1r�?��g���0r�1��3�u��/�zF9�!�,�G�e�S=�^gYV�����B�� �D�������|Q)ƊɁ>8_� �� �b�7H ������;;;?�nݺ��h�7;v쨲m����~HW���䁽p�y��D�#B7`$a$)�eG���ggT�$-���������Ae��_���
 4�:�:� ��ܱA��A�P�E��X5�D-�Do�	*#1U�8%>�F!�7Œ@�\H;737= wl�/�N��Xz�F�����7"
�s�#�o�υÏ��¸}r��,��w�4�c�7�������G�_oh��HE�5���N x��8BCW�V��=��'g��M�Զ�w��0n���1��� �k��������}�+Ж,��ӮzJ9�? .M�R��R���ёV=���R�ˤ��+To)+σ���B�^R���e��\����{����J!�B|`͚5/��RI��"�J��� �W����������a�Sʪ����q��'��,�k.W=��<;ol8&eF yJ�)	݀MB��@��@D��'QI'��N��ˎ������#ͪ�ke-4�o�U��Ư�nv^��ϟ������_/�I�*��E���w?�^���]�$vƒ�g��g��8;�zF`�&��jP=�&h�3�H����h:~�l��F>R�:�t��7�N�����a��GC��Γ���� _����������'m����x��4�����M���6�-�U����-��XGG�B~�ZF۶m[���[�[Tp�s�G��z���h�ko��z��%��wK)o��訬�X�T*�g n�RV�/8σ��fx�:U/);�D�#�l>Hʌ����TORB��d�4�X��P=��|D�6������#N�G�G�ke4	-Z�H��^'=����ax�x�ъ<�]��ke,�'ZP�0p'"""""""�b��]�������R^�nݺ'U	��۷�q�� އ���ǳ�����*�}?2T�q��˟���s��U�Q��R^�������7^x�GT�
˲���R�KToQ�}䡊�ۉ��D$
#�� �{�1x�4�l�=����HZ$͌��h�MDg ���z��  ]'�,\/sc�v&T!��#���f&�G��4":3��x� @z��d6=�9��焦�t�ԢU�"�JYѪ    IDAT~�����������蔼��p�0�wU�a� p���Tj3��׮]���AacYV��ǹ@�>��H7��|�q��0p�9:��"��v��� �B\%��{˲�r王.���QA&�]]]&��0�����n����U� ��	�0�'jO�5��,���7��_cN!��0�|�n&N�G��yDpB7N�8��C��<;ig�9��uӧ1�B�@D�Ќ(D!Ҍ�!t~�MD3$�|����Y)�ٙ�k���{�z�:궞��#�"�[�_'53a������o@[�b�j�S��R^���Χ |zݺu?W�)�,˚'��w)�U ���BLf��l�/ =�z
M 6/k�g]U��?x���Z�gK)�#����/ܮzL�������ػ|�y����<��k!GGTOQ�����q��'��,�k.W=��줓{=�tr���:��:��-�B ���;��#
�0!"Q��ND�"];�,�t�u�.ѵR�yҵ2��t3f��5"�	�n�̝|}�p�,�MC'������G3 �ȉkd� �7HRŹh���֫�ADDDDDDDDaT]��͟�hiS��/��RޞH$Z�reN�� ���\-����!ـ�p��Ix[�z	����!��_�m��oޣz�D��B�ǲ���������`�ҥY������k��y�<66�> �U���!8���踝���p�;b�g�q�8������;(��'4=��� M�c=`j���OD$B��O����� ���	�'��R��F���BL�c�^+�(���C�	hf��?Pz��-��\R�t��� ��>9~��O��g�^ɛ|�����������kx�m7¸�v����5~p������[;;;�B|�����Q~�k׮����_!��v�{���x?�v�b��S������w���'�
!.���ܨ���k֬١z�lܸQ_�p�%B��<��+����l��[ �t�^BD4eB7��ѩ	M
7�(�BD�[B�?��V�|�����#������B���T*����n �tttت���eY��wpp�ͪ�������}���g�i0��1羻ii�X�Z������,�E)�w�xp��ջT+')��J�.� ��œ�IJ8���ʋ��M���N�+`�ۇ��͓iR�?�� �S�ԏ|WJ�D���e��W�w�oQ<Ƿ��Sp��?�g�0p�3ׁ�O���6�9�T��s�7��{�eY[�{���u���T=�,�JH)�&�xW*�� �:w���~�I�"""""""""""""""""����Ys�_����U����#�c�e}O�h6����_<�z\)X�u��������r��=~'��O��z
�w���#p>sc>rohR=��.�R^(���eY��?�4�	M�6�^�z@���J�R+��
� �&������?�#D�����������������(T�|�����D��k�R�5Ms,�J�BJ���utt��z�t=�����m_"�|�� �B@J�z�������F`,�z	�� �=��|�0>�i��Z�s��]q���*�u=˲^B����!6wtt�V=�T6m�K&�k5M��J)/�R�Άi�6����T=����������������������s�`��������E|< X�u�f ��<o���h�%�\�Q��4R����.�!�[r�ܹ ��]�34�ܭ�zU/�I`���`>r��'!�����`��r��� ˲��[ ;4M{QӴ�ozӛ^B��6�M�6�jjjz���yB���`	 �wR͌g=�� �S=��������������������<Ηn�a��V_�zM5� �i���˲v��b��y;5M�544��ỔR�رc��y�=�[�|Ox��5B�g���ط~8ҭz	M�ؼ��%m�hK�����bq�S�*`?�}B�CRʣ z�� z H��8Ú�9��(��B� �y^��@�F)e��EJ�P� ����[U����@ڶ�)���z��Z����F�5���ADDDDDDD4#m�2���z�3����������D"0��	ڪT/	��B��R�}R�c��PJy���i� �y^�}����aT��PJY��@�xS8� �D���U�Ұo��]�������^}��o@䣷 ј�9ap�s&��~��u]�_+��߿[��缋��䮗���I��DDDDDDDDDDDDDDDDDTl��7�����V�R�&�fI)g�xbX���u�����{�jO�ר�r9؟]ϸ=�4�h��+/����@.�z
�o�]/�����1�S�������������������'����f�W�z	�䲰o��坪��40p(���OK����|y'�O]��DDDDDDDDDDDDDDDDDT�ң�o����)'3cp>�r�6�Sh�����pn�02�z
�2�v���xr;U�l�go��ڢz	�2rt�'?����0p8o�.�7r�O����{Ά[�\N�""""""""""""""""""�mþ�Vx[�z
Q��������˪��1p�} �}��U=��l��l��� �Q=�������������������?�?�WO�^BT>�=ȭ�0��{T/�"`��p7����oL� �O�s��sUO!"""""""""""""""""�σs���~�A�K�JN�{�u��n�S�H�����}�!w�TO!*σ��;�~�+��^CDDDDDDDDDDDDDDDDD�_R��������uT�!*	�s;����{\�*"�a������z\�����18n���c�����pn[��UO!**�?�������)Td���s�|�Kp���\S(��^8�|޶N�S��������������������m�������B4sR��ރp��<�NR�C�}�p��,�˪�B4m���������v��BDDDDDDDDDDDDDDDDDX��>�n�ޞ]��M�̌����~�[��P	1p9��_���5��R=�hʼ_?��?
�߫z
Q���½�?�>���%DS&�tù�:x[~�z
��
 _;����ܬz
ѤHۆs��|�v �S=������������������(4�m����ܵ�}��m+���<�O�*�b,�[�>�u��T�!:��^8�|ަ��^BDDDDDDDDDDDDDDDDDZ�3O�^�񣪧���p�0��@���^Ce����~�߾rhP��7�;R�}�j�ݯ��BDDDDDDDDDDDDDDDDDzr�n87|�o�TO!z98 �37�p�
���y�-8�?�u��B�g�p�:����^CDDDDDDDDDDDDDDDDDT1�� �O� ���!m[�" �ܹ�ǯ��|J�R�P=�Ԑ�pn_��ˠ���3�zU(y� �;o����)DDDDDDDDDDDDDDDDDD�IJ�O��o�������^D�ʶ�~�p�>Om�`<���I	����Ŀ3.��+�������������������������@v�}����Q@J�s����pn��f�^�x�;�/7}�WB��w�{�Ғ�����E>:�������������������ol�7��|
ƿ\44�^Da�p���> ض�5��)/����{ �y
��? �p��EFR�����
d�T�!"""""""""""""""""���[�]w��z7�?�k�K%!�s� w��z
�w:�ܿ��B��~�{�HD�$
	y�ν_�|鷪��dd3p�:��s0�w��y�QX�6�G7�}t#�8�א�0p�7�\�?z��,��]m�*Ջ(��m��!"""""""""""""""""����^��k����A���S�>��������w�T����{�����RD;*6D��Kb�(�{�)�?M�%��D�K���Q@�Q��.����r~l4�9��3��,��uq%<�s�����0���Q���(�Q|�AHF�v�~�+9O<U�K�ˑ�kw$ę�����|Z*�nw             @7^��/�P`�B���$�aG�	�J���(�ɇ�a؝1�w�a(�h�K�u�Ew^%$؝
1�(�.���
|���Q              d��&�_�c��r��$G�vGB�ko�����u���bw���9�m�<K����}�9O8Er8�N�c45*�������      �>j�/�Sb�~�,fjٲQ�3���jWXS�?L�0d��ؠ5/���R��z�0^q��Y٪]�@/̰t�,wF��\w�ҏ!S�*_���w^�l�x���Q��oS�C�JN��Z��KT��,�~4?�9�2K�����-�O��?{~Ir�����7(��CԲe��O~L�����KIU��oU��ȕ��q������3�d��T����q�\�iQ]���\��|E��z%�9��q�: d}������7Þ_��		*?I�G�������j+�IȞ�^�wӝJ9�9ݞne3hkUk�VU����翷���p�Ux���:�y���s_]�j>���O���Ú��Mw)���W����Oy<܈�_x��N#c��g>��U_�?�ө�K�)����JM�^6�ϧ���]4_�sߑ��?�v:Ux�8e�|��zEu)_C��|��<����W�\y��^��*}���F�^޹*���hiV��3԰bY��t�g���)���Ժ�T����Z�n�����~�ܭ�C�Y�0�Z�E�3�Q{eyXS$�!�g�z��E�'^�@kk�)�_�hܵ����E��=5�����R�ح<���ժ}W�Z6�W�¹j^�:"�"�+����7�5�Gr]<NJϰ;bP��e�O{B��
�� �8�-طޅ""�����rp��Q����-�^�#55ڝ{���p�c�Mv��Mo���ȋ�     �-#��[�ͻ����C_�@��t�������=��2�=AO{i�Ǭ��n5n�>Bæ�"���e�S�叿{ήV��2�9~��o����s-�/�I�:���J꿿u��6��f�|�ŰN?�/��_�^�p���~l���LH�!/������l��t��>��a|6�p�4l�kJ?|Dؙ$�e�:}y�n��9\.����;��u�>��v<����=����6�����U_��B7�ө��y^�#O�~�WS��~|JX?;\)�:���J�g�N���?պۮ	�f�x4�O�P�.�t͝�>���%�s���ʿ�Ґu_}�>?�Z�Í��������������+�ƯV�5ߠ�?���^v��h^�Fko�Z�%�-Y/V���ߩhܵ��Y=�]��qBX��-o��E��|�|u�a�����+�����o��Zsͥ��dQ�s:<���J=����|�u��'���lG�����|M�Gk难�j}��3Զ����?L������t�]�x~F��z�0��IIߏU�8K�#��y��^kްV%��Q5���w�&=C��/�k�ْ'�7`"��])���2֯�;
��� �O�5+�������v������w^+�̧hn      ��J�U�ޓn���E�'u���7ޱ[s�$]9Q����H�����jn����&X�~��=�<k��%��P��~��G�Q�~��>?������.II���|�q���nnGh�#O���]���|�Q��\�R����G�}~�'���.u<��plxO �=�<˚�%)��:x�r�E~��X��_hys�$�:�b%����=qgd*����L��^*�r�nc�G}o��2���e�풔r�A>�5%��lM��Rӂ��Y!g̙J;���LJV�%��>ߕ�����!���R���V��Qcvkn�:��
y�w��9ݾ��pܵ����}n�}��vI�����=��RՁ�����)wF��q`��z��OV���u�۽'�!~�������4�#l4��[��_�{����7�V��X<_�_\'�ӏ˨�wvj       �P������=B�G����t:�d69��i:�y�	r&%[�!�$��g�^�3J:�����U�>S	k>O^~�Y�w	�w�&gR�ܙYQ��h\�7����ý�s�����!��-w[��캆;�.���Ec�	��|��M�2���Z�u��|��A�׵�'�?��"��q�W�}3SR���p��Ɠ����;���3_o��n�{D�}]���:����z���p4e�<F�g��ľ��+UW�_���w^+��w����D��Q�E�G�$���S�K펃8G�;"�X�����M���F���zX�w]'߿�QYnw$       �Q��[���hnr�\���٣d:�LJR���Y�!�4~��-�6|�\
�6�E�ʝ��ɡ�¼���L�����q�WQ��BiݲQު�Q�?g̙J
�ĸWN�k5�����?�#�,ݐ����LH�|]��l� c������Դfe��O�o��G�	��Pװ;�Y�3�7��߆'�g�:����ؤm[�|5Ֆ�hoW�7�{-�PP��3���P��ü��?��uJ�u�FQ_7!~�ׅ+y�4e6;����?���w]/��se��{�el\'��� �oR`�b[ޫ����c
,�X�{o����;�Q��W���&��{]�;���Gil      �����x扨��s�Yq��]R��B�4(u4�awuK>T�sŖ��^Y���:�k8�����ˣ�Fg��n��~�@k��Qz��ukT��G,mj���i�=wDw�S�W\�5:����T����,]ו����C-]���Fm���hk�l�@{�6��+��j��N�n�� C�6��NZ�-_;��,_��ϫ��n�߱��i��S{yYT��}��Q��n)����W�E�ɕ�fw�}J�����Eu��O	�	.�,y�A���OA�gT����u��/͔l��Q`2V~)���{��
,_Bc;"�{� !kWɷv���<�<�N9S����qvV���k�/xOj�x      ķ��T��u����T��R5~�"��p�\*��*m���Q_+��O1߽����ӵ��Z�&~l���U���?\���=�P�۴��WS���k�k�n+Q���W_v��*{�ʦN����+����w_W�Ѓ����s��Ah�{~oQ��a���z��J?�h����x�+-]}��5h��zU��_��V[y��|��ۿ����U��C�7�G}������U��t%:@�'����J�/wgfE|�X��W�����<�xyr��z|��3)9h|�S����f��zkkT��b��n;ogew�R��oWE}���z�5��X���+%5��\6A�Ǟ4��D�P������'*����+�����&ӯ��Oɻ���|uu�[�D�[6����R���#�QÊeQ_�j�οX��������>�ߦ���'�J��Ŏ�S��#;�ө��j���7g:*w�6����]��>�;5���K�32�1b�z��gr�g��u�)�9�lU�}+1���Z�_�%�[/�u�)r�}�E}쎅.2�^K���2���=�*�b���O���sr�r�ܧ�!�*�;�$����/xW��?e~D]RK�jwE��      ��׮7M#*�}�����[
~v������h���O�c=�� %�֭�,J?�Zѩ�'҆f��^_��S�F��%)�Gg�����"�c���|_4[��pOмv��׮��q	����>o�]î�4�_t�ʦ>iwI���J��O�2w�'�C;��m+Qe'�vzO�Ѵ��|�4��X�O��k����!����h~T��:�Tɤ�]NgT֋U�e;����;ul�%�L�w�<GMkVF:Z�����ܝ��������]�x���龻lL[V,U����-�~r�J��'�j�|�]�V�Tݒ��|^ջohۿѐ��P�q'����_������y_��*��w�_���G'�g�9��}�gt�1*�X��ߓ��J}��=��7^���C�:i��ǜȮ�1Ĩ�R`���Y��    IDAT�-�;�!	���5�;     @��5�oj��+-]�οX�3��;J��RR�>b�^��u�ʦ�ྯ�}�1����h�5*������(@X�λH%�;B#��v������VI��\�iA�i�aCD�3)I���ɏ�%��UZ3�r���8:��`���Jv�W~eC:Ĝ@@��+��c9r��<a��cΖ�tc�ϧ��*�x�_.g�\X�[^`�@@��/������:A��O�
^��?�����{���<Ks;       ĸ�����;F�d�t�����&kԩ�A�H;�p�v��1��%���Sϴ;6gB�
.gw�[.�
/�����ٙ�dqX��ʫ��x��׫��I��6�z���-N�x`T�������
|�����k�el�*ߌ)j�i�|��I�Kin�����1����e��~Y�>��<�D9�;Y��}�ֳ26|������@j��;,Ի�L�}���iH��2      ��ط��N>M5�߳;�^ew�q!��LJV��%ʉ+��OR���[��kU=�-�c a+�l�vL~T��v�� a����*}�!���tYB~�r�8O��|��(QѶc��?xGy�TKz��7�X����HM���c;�
9Rr��U;+�_�T�E�dl�`w�w�c{��/ϒ��Y�7��N-��;Z��?M�O>�QWkw"ؤ��B?���1v���s�       Ĥ�k��Α'�WP����b����T�I�t���De�<A5?�r(X�~�'�8����3�QbQ��m�!�y���#�v�j��R�����R�9h�+�ِ
�Pױ+=C�^���Oِ
��ҭr��J,
��}��=��]��Xn����oC�#��QƢy
,��{���GJ.Z_#��U���*�t�������iw ���kvo�s���O�����b����hqŨ�S`�b��xD��/���_���k4�      @�0��U1�ش�q��J=h�ŉ�&�����|�B�Ic��v)����c�.�
��چD@הϞ�@k�i��ʉ���z޻j-�bZ�}���am  u�.Vӷ�MwE�'��rY���O�3�1-�;T�Gkq ��j�L�=Y�'AO`45*�h�|�/�K�{���#U�_g!���n��s����[��j�����1�w�4��\��������]��?����eT��-��|
�Y)�sS�������
��S�#Cx       ĥ�Y�*��fZ+?��4]�}�i]<����e�F�.^hZ˿�J�RR�t���:�Ϊyg�D	�E'�(P��gMK)CT�1�[Oy�]���W���-NtM��3�on2�����4�1ü�e�c��(�b��O?��[��{�-�?_���+%���x1Ǩ(S����{��_sq�F�o�(c�)��)xN���"�X*ߊ���r:@��s����C��x�i��f�)�v��V�X�Zjo�;        ��U�T��k�u��A��s.P��P��
��]�F���<����ľ��<p�Z6m�v4X��x��F�4���T�.V�L��K V�M����.�������	*�۟lJtN�3���;�J��M�NuK?�!�5��xI����<���jE�S��wmHt���N;_}A��O��9KI���t������0dl�(����k�I.����s谎��L^�X����X�Jƺ52�|#cW�ݩ������UW����Ҋ��KRb�����1� 9����~r��\��M�2J��(�"c�F�����;�       `PV<Ŵ������q*}�AR�YB~�RnZ+��C�����Y������.^��uk�r�AA��qת|�4)�!�9��Uݧ��y�IA��K�k��P��نd@���U��s*�Kp��ӕ�� �l�hC2����S��7�T�8�8�?L�+��!�9e�&���qA��;\.^~������,��Y������`����ؼA���w_�9���c�A=�����+LM�;i��}2ʶw��l��a��Im�v'""�;�ﴵ*��+i���aq���ӿ�S��:~X�*��W���d_���jig�eҶ�2J�(P�E��ew4       �M�V���*��A���&h���h��/�G��ӱ$^�j?�����w���:UeS��"",V>�Y���A�I*{��,�kC*��ʊ��6��3��뼋T��tR�WV<E�W\-�˵{��P���w��'�峞U�kn�311�Vx�Dm��-6�:�u�&�,Z�����/�R��zD��z�EO���\%��S��C��m%2���6�������o?9���;�
�rl
���"���Bڱ����t��K$���x@������瓱u�����J��L)/��ٽW�ٹRZ���RZzG==CJJ�^�@@FC��� 5��hl��e��ʨ���>�?����       �ʊ��6�{rr�w|q��B�}��xݲ��ojT�G�M��G'WJ���Mю��|�y���צ;���D�;b^�¹jټQ��
�]u�*^��ӗ�ڶ��f�\�93���e*}�����ڐ�<5$ny�v���L�n�w�*y�4�"��O1mpw��)��KTV<ņT��JMS����~�h����)�j����������+,�#7O���~´t)-����g=���Z[��GX'56(��񿪩��%�Y���
����t��g�uR}��M�w���@�[��$IIr�ܒ�)��t�%�Gjn��+�������OFSc��,       ���f��j-ݪ�~�jE�'���1�X�LHP��Mk5:��k͗���"�LHPƱ'�f��Q�	kZ[U��t����j�q')��aj�v�ɀN2��|F�����R����u�h�.^`C0��ʋ��6�;�������̿lH=��^���:�� �ʊ��6�;<\6^��?1��/T���JzpP�hܵ*���P�R\p�}����j>�gq��^�K���ۿ�8R�$�[JL�HJ�\��'ڥ�vlv���Qkn����O��V��-Z7o!��5�W�QY.�b���:~�]%c�26���}��c*�e����       ���W��gLk)CT�q'Y�(���'ʕ�jZ������WS�ƕ_��=�Ԩe���g<#�g�4��q�Z��ʗf���h�$�� ]W��c5�YiZ+w�n�ŉ�'!�P#�5��W�Y��Դ��/�ԴVp�x9��,NtM��u�}�+��Y�&�.��}�
.gZ��ש��E���hj����_�dsG��=�kW��ϰb����ĦF�ہN��         T�0S���.;���'�n:޼�[��l�����7?t�7u�\{e���{Ӵ�w����[��@K�*_�mZ�:��p�ŉ��++�b:�PX���ϲ8M�9\.�r�|b�\i�Au��U×�ې�TV<�tܓ����.�8�5;_Q��j�Z���x_�JM�;#�ӿ<9�Jr�
.���^_��W�<��;�����M�  �/��         �0��'hk��A��V���Pێm��$S�*_yNE&;]g�<FɃ��e�z�� ���L�k�����~�~7�"踄��J|�Z6��J>ث��'�w�A�΄\:N�ȆT@�O�c�kW�G�W^�M�_�6ON����A9����>���{q��)��#���zE�������T���6���C�W\��K�*���K�:��LLY�Y��-��M�U�{W�%[����Z��I�|q�d��%���[Z�|�P��������Z�ٚ`�hmU�s��s�mA����S�!����]Ye�c��wWk�f�=��� �y��        ����o���ܳ~��ߐ;#���Aʊ������
��h}�Hr���3��,ܽ��q��j�Yazl�Ic"���q�Wj�b�i��	{lJbAێm���]�Z��L��K�>B���H}��IɃ�D��]��Zb�Q]hoWŜb�Z��#�vؑ'
Vx����2��.� ��������S��[�'A�*���i)e�Pe7��@��'/����ﯜ����9oʓ�gw� 峦��ż���-Nc�@K���y���vG �	�        ~ ��H٧�aw� m�J�ſ��%rge[�hw٧�n:Q�W��>h�[�����Q�F8bIY��qOn�r�>��4@ׅ���II*�x�e9�ԁ�gZ�T_��b�j�-[�Q>{jȧ���dq�`���ʼ[�r��׮��ܰ^�3�o�7����:Fl���*�������\U�?1#�����Xg��Z{�5��L �/4�        �p�g��Ty���d��
���.���L�k�5�y��y��g�)WjZD�!vT���ڶ���z_}��pX�蚆ϗ���/Lk�W\%��cI��~}��O	��j�_�l=D��j���~մ�{�J,�cq��9���2o{EYT�=�M��|�9�Z��S�<h�ŉ�\��d.I�1�I�q�ۣ�K�s��]�MMj-�jw @���        ��_uK?�;�����i�J�Z��p[�X�C��,�~�i-Ԯ���y���2�;)��;�_�s���R���cO�8�u�3�6O�/T�Y?�����\e��u��ojԺۮQӷ�,[ѵ��'$�w��*��*�W��Q�w��f{�>"��x��M�r8Tt�D�!���>�����V}���Lk����3)��D����Ұg_PBQo��  ��         ���z����y����Tb���"�q��i:d�#��4n���[b�T�o�W�����Ԉ�Cl�|~���M����,N=Y'���<���G�|��qA��~M���AM�.��'*9��q���Z�/��W?>E5?��z�N�5�_��i����r��Z��J��v���y�r7������_DtNثm[I�){]p��Y�'�]�Q#u�3�w������t���B�ߟ�2x����f�}�������
���T6m��;;Gy�]dq��J(��~�� �8���         =P�c�e�=hiV�o��UiQ��T����y�<y�A���nЮ�^�<S���L��}"_}]��j�S��#��u��p��.��端��W_P���j٣OW���jٴ��`Tp���?�����ꉗ�~�S!R�W��߭���|�2F��ϖFm}WZ��xÊe����Y���Bވ���l�des|и;#S�����gM�>�:�����k�=�+!��K�:SR�y�I�w�ݦM��λH[��[�"6+�6Y9c�w&%���+�}�}���<e?���RRUx��_x�V�=_��|�t�k���Դ��=hmU��o�^YnQ��T��ڶ�(�o��Z��I�|q�-�ʦMV�˻t�+-]#F*����}>���{�OT��k��	 ��hp        ���e�~��vǈ�@{�*���Mw�҆��#��rCBw8\.e�0ڴjW����S�;�	O(,R��j^�m$""�M���K��B�p������w��'X$8���w�x���_k�e��
�V>g��\w�iW��IQmpw8��ϷǛ���U��}��lQR���jE�'�|N�X�?mmj-����׮Vˆu:hʬ�������Q��U��;��	��/[��5+�z��Z���'d��6$�<gR���|��L���(�jX���<U���U>k��}_P-e�Pe�j?^hy�ƯW���7�|^勳T�?뀿MV��#L���oT����� ث�?�         W>{�mm����,͒~�1rge����|Ҽv��ʶ�ֲN��l�]�[7�f��Z�E�ɝ�eq��I�˗;#3h<y�6�A��j��덗Lk٧�i�4Ĕ@@�3�6-%��Q�Z(rj/y���NɈoe�SL���{ƹ��.O~��a�O�T	���EB{����ӐOH�7@i��8  ��        ��U�T�������϶�y+{���-֩�d�^ϯ]4�|�Q4��t�!ҜI���i�N�2���rY�V6m����K��_eC"�k*_�-C�i�h\�5V��P���݀��V��+��4������DW��%vG@����LkY'���AC,N�}��V���OO�9�,� ��         qjǳO족r�e9B�V��c����I0=?�ȣ�JK�ftج��j^�ڴV4�Z9��]Ӽa��>YdZ���r�gX��S�*_�mZ�<~�Rfq�2y���)�ޮ�9Ŧ��a�*���-N��?U�c�QPV������@�Z�Y���3�%lq @<r�          �i^�F��?Q�1��
.�m��[���GJb��J<Դ�1b�2F�{n�ۣ��F�z�[aρ�W>�|ࡠ��"�~���y݆T@�OV���]�iʿ�Ҏ]ށV6�)����)�c���{n�!�5峧���7˙�T+�p��X��k?^(�}�͝ط��L�%h���Lk&]����r�Fպu�j>�g�d�^�_����Y���uO�gK���s��=��6� ��        �XY��wWZ�z���g<��͚0":��Sip��v������+yr�jE�'����W��<�l�`�iѸk��}讶����rN?;��w�E*y�6���[�KUo��^\T�9�,%�����׮�D��H;��wK��׭����me�SL�[9��Up�Xm������[��tܓ�mq @<r�          ᫞��ZK��֊�]#9��qP��Ӣ:���$�#�k�^��vU�0ô�~��v�ŉ�.2��4obO��O٧�aq ��ʊ͟4�LHP���,N�gǳO��p�p�Tx�U6$:�n�Gj�v�i��ʫ��x,N�}�0/�� �	4�        ĳ@ ���I�������e�{|$%�*P�Euد|�T^�i�pܵ����9��՚֊�M�8�u��?U�7_��
/�J��$�]׼n��-1���J���-NtM��u	���=�<��  `/�        �\�K��o�7���^ce։��LL�����>yL�׀��+�U��릵�3�UbQ�]hmQ勳LkG�T�!�[���Ϙ�{r�w�O,N���x��+-]�\bq�kv����U;Mk�����4��qS�����$ �x�;          ���Ԩʗ�6�g{���QY7{�y�y�捪_n�{枤��Î�:i��O~���!��OQ�y�;\n�c%�@���U4a�����sϢ9����W5�{�����s�����^�ZK�(��~A5�cĺ@{�*����7�TKvh���EK�ࡦ��;+-N �G4�        � e�STx�D9\���3!!�:�u�y�g�P��ӻ<e���i��W��ӏ!wF�|�u]���/հb�ҏ<&��k�������r��!�k� �ޮ������_ո�7��xZ���wA%�că�O���M��x������=�\�Z[�k�  ���          辶����e�;T	E��P�G�5gÊe����;\newRXs"��O�;�-\Èw��*��fw�[*_�-C��1��x�v�����m}o�������E�-N �G4�        �V6Vf�>�t�q��j//kN��W��MkY�Ƅ5'�K�ܷն���@�V,S�W+���[]�]o�lw�[�M��|i��1���M�lw�n�}����ڛLk��z�}���D �xD�;        @Q��5��ʒ��B4��,x�[��,�k:�}�����܈}�߯�YS�]��
V6�)��v��rgdF�������M}R2�c �R6�)~��1��4��F��}jw�.���*���5l��p�}!_co��8O
 t���          V���� ��S�������մ������Ok�����|�;ԴV3��n�]��<~���?����+���jZ�M��	�E�믔:�09���x�3!�t<�O?1w�^�j�^���>���>V�H�|q���t�\)�Q]'g̙p�}J00�9���-�`��b,�  �IDATÝ��~��R�G��+-}��:\.�qgRr�����2U����f<-a卤�w�Ѐ�~���"��N?��lm��5|^�}�H{g�O�7΄���Ve�x��9�{=ޕ�a:>l�+2|�=�뫫U�����S��5���Լ�[�-�X�#O��:΄���W�;�|%���Z�+��l�Zvs�=�=���}�<y�{=>���=]o���7ԫn�bm{�!�����Im�KU3�=�~��Qa�~���--����S˦�>�15|�Yd�Sٴ)�1Җ��<���<�D��m+�n�S�  �w        �OH�/�ʼI�R�ɧi��g���UQY�+v�����y�zDm��Q�����^�����:5��LG7sd��O4���3tȜ����p{��o�^�K�7@�#O�;3Ke�&wk�H���i�+ϩ�����F�Ѓu�?���fW�hpx<V��R8��9:}g����"m}����ϫ��S���_�%bn��N:U�s�����}bW���K�g���y�����~�6�0�8\�^eL�^6mr�����>��&�k�iٴ��5�2���*��˺=Og_��|��9B��_�'ʊ'���y���Wp���h���D�{��w�Z��S���A��U�n��@k�oN  �XN�         �;gB�
�]kwI����bNqT�H;�H����G�)�f����#����� �۲�s�kn�|�Pʊ���N�٣O��=��N8����a(wm�'X�bδ�Kt�C���`�cD]b�in���(eȁ��k�f�\�l���_xi���WS��%Y������g����GX����埪�/펁8�p�Ut��vǐ$~��g=kw��0�^��ō|= ��w        ��de�u����|��*�,s�)����{�p�?$�f�yczW�����7>�rg�سnF��߱���|��:��Z�nR�G��:�3m�Q�{O�;+lY�jv]��G������ՙ/����j�/�un�3d�����ζ��$O�k����a^�2��|&�s;��t�r��և~�#o>1���1}�¿�C���uq4��Hk�:�����$�6w��ׅ��g�������W[��/Q�ܷ� �3�ƿ        DY͢a�ײq�ZK6�W�}'�,ު]����a��757�jkT�tqD�oٴA��?	�zo�h��_�qDv�諸O��kz�����>_*ou�ie�S�>wo��˖�]o�b��vhX�L��k��M��	��3��[6oT���a�)/~ʖ��hjZ��Z���w�hٸN�]���뫭Q㪯�:�f�ܠ���P��=L;_�#C}�������ùQ��|AC��?�ʗf[���Z�mU۶���75����:�f�\~�nc��VՆ�:[�v���-_��h/ۡ��>����6��w�.��ym�KռnM�x�ܷ���o�W��s�>�N�߯�g����eK� �C4�        t�a�|�TU<W��>���<QM���$�ڴ}��x~z�bE�9x�[���?�o@j-ݪoo�@{{��X��U��C~������?T������\[����|�M�������7U�4[��+��-���~ޭLu�,2m���۴f�jZ�2��.|5����?��D}�X�Z�E�K��&��lٸ^��1��+�kǳ�����+�Һ������=g󆵪]�a���s��罫�7]e�׌���Z�!wS�o�N���z��:�~�m�ݯ嫯���h�����j��77��řa��7���/U��;��:ۛ@[�j>��Uc�׶���:1)��;oPێm�-髫Ն�o��jgX�7��Z����g�W�i���Z�5�L�׫�YS�>�j�n��є_]�֭�����h�+��k�`���s*{�ɰ�_w۵j��sIR��]eӟR���݊U>��oB�Z��Y�_�P�?���������  as,Zгn ĕ�����t�C      �M\�Fn
o�7D^�aGʕ�f�Z��]-�wk����JKW��%b�^�}�����Q��
Z[Þߕ��Ă"�l�����[�����Hr�g(e�P9����N۶R�n���c��#gBB����9r������o�C�q&�(e�P����0�+�պycD�.����a7��;#S�̬�uKKX��G����D�SST��c���Q��rg�Du_m�Z6��̍b����7�w�3)Y	��C��Omeۻ����+9:׳����=I��n���'�WT���שy��n���_��,��j#2�31Q	��!�F ���Y��6�0�22-Y��zղiC�7g��+5M�����GJ,�#���޾�R�֖.ϛPP$gBBw�I���V�
+  ��� ��     �'��       ���e                 ��                hp                ��                1�w                @L��                hp                ��                1�w                @L��                hp                ��                1�w                @L��                hp                ��                1�w                @L��                hp                ��                1�w                @L��                hp                ��                1�mw  ��-��N}k6�     �[R��        @��X2���;                 N�                  ��                �4�                b�                ��@�;                 &��                �	4�                b�                ��@�;                 &��                �	4�                b�                ������h_Ԁ�    IEND�B`�PK
     ˡ�Z�+�sz;  z;  /   images/a657ee5f-a898-4bcf-bee9-a045b7cf922a.png�PNG

   IHDR   d   d   p�T   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ;IDATx��}�dU����z�B��=��ff��a� E��~���bXu]W�[]W�.:,b �H�!ϐ����=�=�su����ι�UuU�V�ou�Ztͭ���{���p�S^i���6���-��d~���q����n�%�c)E�Q��m2i�΅��Xi2S,��'m��.�FQ���-���Tm�����b0s�;B�~����e�>'Ax���;hW��������߾Om�P�-����sC�z�C�"�"�ZȐ4]PR
��m����5�������(|��D�>u�
e�ڶi2O]�m��$��0���9@m�������+��XҰд�OP�1,�|��� ��r�:�P�����:駙9E�)�3��5Pn�H��~{����mַ_��|���O[�)�٩����~qme����
`q���eIm�ō��!-o��/@Zє��7�dڶ}�|���m�
��-��!��he��x��u��6�o��~������_�$�.Z|��/LW����yf�!������o���h}/�|s�o5$��`qQ�)^�Z�,�̲��n�V4��8Ǧ=�`���e��J4#f4���`ZNѵ�iM4�h�Ry@��Y��3XL��Ч-F�����k6���,��LW���a:U��!�����
�<�.�0�x��N詔<�Q.�f�dw@���H�t5�C?z�v�f�ॕ�g(x����sYRa��]�^��Π�)�Ѡ�fF�Y�o0��C0��+p!�h�Iv;�H�8]���՗
 ڟ��h�4#��H���A<v����A2ɫe�{��caV(�(�Qiy����X����3�W3��@X��?�EI4c��j!]�"�� ,d}�D׮[涯�xSԥ
�3�2�b.CZrbe,�2i#;}Ƞ6�d5k��x�X�F�`��h�o\i:㼹�o�K/<��4�Mc6�*�Y1�g�b�)�L��E��>y�يܺ�652�=/�P�mWHa���H� M��Z
3�3B�����h'K*Mk1\��cC(?z of���.j�X�d�X/�Y�Ҽ���n��iE���1kD�͊��u'�_Q���n8��c�n0e��ym�à]2��ߊ�T�u��=��,�~O;�;=�K�n�"V�G�VB�zR��GV��D�q�[�Y��[.-n���Y� M���1�%B��Y�R3���������Ĳ&X)��X�X)\N���8��������{~���*��X��4#��j藃B�dY֓�P�6�t�H�����f�̥��>�Į�M<�U?!���|�}˜϶ؙ��<�����6��p҂���nz(CT��>���]���߲����[�D�چD".�a�.�߇v3"�8!iU��[ݼ��4j�9����#�x귏����c�觕o,}~�1��WRʂ܈�4�m���$/Ȑ1�6�������ӏ?��J1ޱ��,�u"1":���L��qO�Ik�Ѯ�!:�PuY1��+#1T66b� �x��)�E�z��P���ebJ�p!�BMQY5�=�@_��y����s1��҃ŭ��՚-�]��}��`�Lc�4�E1�8�hV҇6{F�+aAMezN��J�Lo�$�]]���u%P3,�)�c�D&����&�������D��ٝV�J���54���[`�B��2f�V;m-k5�uz0�?.�d��8M3ᯮ��ӅvR��OΨ�l^����C�3���'�(�Hf��,�o�&�^�n�^y�;_�n5m��F<���*�d�[�8��z`��J�`_��D��;��!��VRן,s���@g��p8PQQ!��O��eg�����)Y(��;��o�.X����ΚfX��0x	����k]#�k!;w#�3�:넥PK�C�`���:�E���=S\\�?���H*�Z���Ls�K&��H�h%h]ؾ�!<���(00�L*-�|1q50	}�82� ���X�N����o~�
�;C��W��";f�A�Ě�O���P�a�>2u�R*QP�c+t{0��|r(�F����f�ʈ�g6�^3܇�ۿV[�\d)n���e������Շ�o�C~4�r��U$���i�%I�T���좉�!��:aŮ#�#��Q�%e�����E���}Q�����<�h����4GؿEE"qv�ˎ3��B �%s�%�/- �3s��lᕖ`+�f=+��i�\f����P�I�ξ6}��-v~:����-�CH�&�|���{&Q�b%�z{�EgY�:����:������m�ɫ:��x�x�w�'���]�ǡ�*�t|�܍k�����F�UR`��K<��[0����o��zW�>QgGR�����'ahC�=�ъZ����Qd"���z��ƞy	�?7	�Q2��C&6������ߠ��sz�p����.���HX�2q~>����Iv�2ы�Ƣ/�'��g��iH�;}U�V�
��t�H��)�����0r3C�0������$��̶<p)�m�o�9hi�HN0>{Y�����E��CB�i|��jH6R}'�����4A�kj�*L���V^)�(��a���O��@�k٢�$��5@'"9������D°R{=Grt �8�d��Zh�{��TYEmbЏ����*�4�3�K�ӥzV�Ok_h�� �B�A�C�n��g�gƆ�coB��Y�����j�7�L�����	�W�L�c�]O���m�.[����u��P򳏣���a)��؝�G���!����|U�y��ct��H�1$b���gP���g2��?���J�$������-����v���'�p=���^��@/��%p�{���;܏�+އT�a��䋯��Ӆ���,�u�QMe]���G����:
^�!=Ǡ���#���,�C�����X�H�UP�e�p����lM`5w�.\.�f
7N:;(�*e�I��I#�JqzR�}�t��S��B�ij�V�DM�O�����]�@�O�~S�Q�-�
_K�*�O��Y/�Eu�?�pԏ�6�c1�%��t�sa<�l)�bvH�woC�?��.+��4�.�i�ҎE�J�5��@Z���"�=��Ϡ�̷kl4�IHU.���v��t�LP^�R� �i�T����5H�hB�:!���	!XH�����-��ό�BO&��0��#6��C���T����a�R����Ӣ��	Ȓ�>Mb��!{�P��nc�)�,>3$2��i�fxኘ�0(Ғ:Ns;q��C!��yU���S�c�7����k"@3 ��4�ii3S�y�Nz�J�X��e	v�"`�;���:�B��
A0-A��;��7"��FJ��H�B%]1y�� ��Ĩ(\OO�c�G���DL��J�[�x&�M0I�F�X�'��oC���n�`�D��L���H��hZ��	�}$@D�т�1��y����|4J$#~��I%��f�"ZS��� >�>��UM����f����v�_Nm��5<��`�D�'�UX���H��~*�#�l��*����C�o<uJ!fRC��0�K�����Y���ob�F����cV��?�=�x��&��e�~��%=
3#��U^�:���ue�8�)"��9�"��b\�~9��������i����7�?D�_nw��M�L/��M��s���s��9;d�P�=�O8V-2Z�du/FN ��_/�ȱ!�0՞v��}���%Bm��ϬϨ�0�zF�N��GF7��r�i[8](�X��uE�������$�����O~�n9c7]������Ӷ#��au�浈%�L�o�Z�E�$&�7�N�Y][��HN[��� 95�W_��	��c,>�N��w�����n�yYhln�燈����k���Mm��a�/&�Y�q=�B�lFt��z�G���0�g��9�^���f��� �iaC����!۬8���9h��=p8��$@�
��h��K������o����VU��uo�R��[i)DШ��d"���
�k4{�f����@����Ց4	�z��ڲ�O�'�E@����MŨM�\�v���k�ꢬ��xt0���T�(!�p�ظ}��CH�;�g�����,����K���Yh���!�ӱ��t� �L"M%�CX�*o>�?��C�y�dt6�����ק����g����eE�>-���/������x�p$f�8����ԑ� ���Ț�!�+��	��ʜv�=Dv����N�|�KA���7�B�1)�ljNQ}�=��;d�!�H���3��=���@s$�K�feD�f�C$FL/ll��;����V�<��7#�XN2�˕v2jB�˝�@�����D��k:��߷dt=Nl�p��\�5&�tQ%{|S��3C�sP� Ms�Éd<1�������d,mY��7�wS�_�wi�w�4��~�~0������Oi�Y4L���%�00HD�&R�F;�s�"����*��;�}���e����v���'F����f�&�_}��}�:�Ēp��������n�IcwN���:�r2����l=��X�픭��２�����׊>؅�������쇢1d����1r�LzA#���(�"�P�u�[�!,���сa������rܰe�	?��r�B;�Ey��a9�t�cU�;ػހ�؎��!A#�$��meY��s�5@����2$�	bH�]2�t�1c����\=�	v�����;��=32$�}n��a��ײ��}q�"��8��
�{��@������1V��@�4'8Dk���o���",;��-ȹz�����:�A~��ާ龳�!|����v�a�/ːI٭�myF�$��bV����b��w����A1CF3Sǿ����
s�'��?%|O�Oe*?v��fq��e3����-4���F{���>���^�f�_�������2�nN&S��=��b�,1�E�����F�B��b��n�Ӥ/��a���r�v�z&^Vp2\�2�'Ơ%�0Ek���ԊL$�����Y��U�����@g�^���#�u��{��뀕���2�#ƭ,J�}Ub�����R�B�׳�a��HRȯ��"���J���$�����
C_�sti��2-9$�)��UX��k��D��vH�D�}��C�"r
e�\���F�H�����.F���_q5��
��m@��qq��K�@���&�x2g��E��h�_��I�\04W)�Vݢ��(�{(�� �~qY��y�~�5(�{ 0=��`��P���pd4��ë��ِrb�x�LJ��W�vHn��gZ���Đ�e5,En��ȁ��\�$¿���h�I�7�#nm?�e�����]t����!�~z?�'3��hVL��(+�'�'�![&�Q�����PgL�f��~��AKP�@.f�Ёي6[��\�~Y��� ��K��ٞ"�'q�z����Bv:Qt�F���?���W��l%2�\3�r*��������)l�횋��&
�b�|6��٢������I�e2��8�W�2)5�XA.dk�������0���,>�\�[�b�W�@:�l�Ӫ�8�!C�.��]P|%P#!�D0�³(�~�����
{0�QKƌQҴI_�@xYhN4�0��� �(%�BɆ�z��"Y��j\ͫ���#��+p4��:�t��u#?���V��?�A��v��(m���b���#(��5��p��'VW��?$¶��8����Dp��g!�櫰U׊	ȓ�VY%Dw��A�ܙ0� ����m�VQE�"7��ar��L�@WS�@FB�Zb$$Y�s��1A�Ǎ�l�8w޿�E37N�1	 �z�D���C��XfxXYXD�XQ��fأ��Ӌ������G&M���`	b�ٽ��	�[��i'��:Խ�dB�GM��ޤ6g	z�{�i��썶��iO�<t@(��Ѐ�<�N#������V�
���;���$���[X:�z�ɈP��(�w͜La1�Ngo#�#@���pVz�a�Y��ٵ���2�cN�هk7��F��wb����U����H��B+�1�� �1%�oG���D�o�V��.�/��s�a�0_�
�e���3�Z����d��ayE3"yi�y�V��AݎǬn4�^��[����E�"�cq?~/��2:;;c�_V���w�Ia��~<m��Q|݇�#�X>�vZ��|�k_�/cC��=�1�G�B7�T,��A��r(ⓗ�gl�ǯ�n�:&,Di#��L�W�G�n���?�{�)���"Z �a�i��amA����Ah4I���'�4��p䅃�R�(�P,L�J�*�|�g�A<V�̄��-�i),�憢-`e��f������^�+.�^"\6��g������><�������L�1�q��V=����i��W�{��N�����&Y]L���$2v��D�B����C��'�Z�] ��
;Rezv�W��-H?|nR��6!nu�%{�T8��=�뗠{Z!�H@=F��ƿ��+�<�V5��	�3*I�S<�[u��ۧ݊+;����DҒ�2�� �ǘ�@~G1�~��P�?���9Kt8S1�w���x�[��~��⋌|�drF[�ۍ�r����b�)fw	�X�f�Kb,��C���aܶE��c/l�r��c>�b����!��C�¦�{�|��HZ�yb��V��p�57N#}L+��9,��}R'��>$��ܷ�����k�M������ʍh��M��'0�ė���-���3O}�8�u�pa8�"1�����%m�`.�p=3���'oڄ"~�9h�h�ӆ�n���>M�L�q�	����$��_R!]��5lw([�>4��<#'�K���6v�JvY�hʆ��
��꩘^6��>J����U��'�)�$%Oޓ"�y�Wx`�bC�V��eZ9�2��-�W^u��\�(Y@��сM��b�E��х�9�f��!M�C����ڇ����a�V�qZ���c�A8�[HIy��@�	B�_�S^J�,C3K�Y�E+��bS eǓm/f�*$�����6��d;_l�r] y!��?!�0����g�M��9�4pk;w ��DG�+~���tE#}�o��+j��	�� �(p�%^C�=.�Sߘ<�@�Y7Ŕߡh�W�ؐ���%
B_��͹�"[�Ղ��}E4�{C|���p�Q�dВ1X\ޜ��=�(j�:�&�XYY)`��~���	/��"�2CfIr���`E� ���F��w���;9����p(�7P7N��,%���ɺ��pVT�}�K-�U�\�>��Ŝ���0;6	�{��%dx}��_b�m/�ɑc�����,8�>I�e���R#1����*w�\(++CMu�	j��̙���ƻW�p�d�$�h�����'�R(�x�ڍ� a�A�rF����ņ���`�ß�{��<�JL�~�= _x"0�
N"�ԣ�#_DQ8���/��D�\9�+#!�]�E�2��.��d���
��p8��H���c�/ Or�I[,EQ���x�C�#�#�%��=�Xk��bt�0c������5t�n�v䈱`��K0U��g&̸'��tc�3��D��|����(��:Ay$�e��хzlJ+�EO���a�H�����pCQ,S[60�i@D�0Y�G��!f��8󯺺5U����#����h����Ç�q��֬�v1��*2��xb���21&���o3�~�, ���֞��}�8�2+�زb/J<L�4<<Hv��N��*n�?X��"�,p��!UUU���LQ$=I�B]�BkɴL�k�	��-R'(��D"�λ�����+�PRչ���l�%.�,���B3���hoG�"C�|[+�o-��V�sX���&e0���{:�%��԰̜?3z�V�ɑQ\�e+"�Q2��ˮ�h_m�ˠ0[U#G��{��̲"]ŵ��7^Ƿ�������[��pS�EL���FaUk�1����ۈ��|I@� [�Ծ��ń�M���[n)@YYg�0������,1��Ċ�8ғC`��۲
�S����E:�B�Dn'��GM3�FY4.�ˍ�d���Uը��Ĭ8���	�&�U���f��b�J7?���d�󷏡`7\֮]+c�I����}xf�s(&��,�l��l�㍞�4�5��e���@g�S"��}Y�#X��0���(��*����`���;	�T��d.I��4��@� ��P��]������8����F�57>�������>E�8�����Lx���!�Z�
M�a=�H�����µRc�#u�PS4�Uh�i-z������/��T���F��~�`��b�ϋ4d`` c��|�=Z׬1|\s0�Y�q�Dx�wX-� A���7�N�I���	T�!�h&O�m��+�*��[s)uj;��Иe�p�Y%%�������8�����~�H@�0S��q>��=�^{F��`k��\B bU�z�n����@U]����
l�Q�����"�W*.���D�*u����&h��D�z���3W��4F:�	x�⢘|ԟe�n����*�X%iى�{�xz8G�*HӺ��j�n���2�/L�"�Yb���8�&�M/̈��^�S�I[�I���ҁ�"SXI��e�S3F:�}�#���	|M9M�O{��]��4S�؞K�еե��|~���9��4�	�zpa�	����:��'�Q�NzM���l������.f�[IR�$�.�����!�zc^��Z�
Ȭ��ŃH��%f�[Ҁ6��Z"^��Ļ�}�S�np�EƲL7��PL6�H&�Ԝn�̭��s��%9����"�W"�����>�n�B�m�&l�&��<Y%�c��/��ƅ$}�<76���ǡ�3��7�� �Ua�I�����~�N6��[�R��a�<�^	��):�O��}8j+B�KAM���(F�:�*m9^�n'n�����p�ھ����Ӄ&E���2�W#zp�'���ߋ��h��ۍ`�	|��# ?��ag�x��Fr'!\'G�n>�p�x��L�-
��FFFP�~-���j�oWz!�IhW0~��aTUV���6��MU��?���M�Aó����7X�В��t�3���>�I��`�-��a��j���c�h.;����a�:Y��e�Wxx?�������=d�0�a8���|�)A�އ{t'A͙��YtG��Q�i"
;;N��|@A�P&��:E�IG�<St�2��|4>��b:A�k@(�0��DC��**��r/!}�z��ć�,Q����O�O���&K}�=��1?�)��p�s������y�#�8A+㹗;e�w;Ĕ���G04�4 Y͹]�*xq��Z��>.ғ\�Z=|P�K�rx9��l�_ºj%��<���ݹ�!|E�D���"��Jp�����&{g��{��9��� w[{��}��dk:�O�'��
�A���A�P19�uB��đ+pP��JJJP[[+���ȉ�jG�E6�<��|���R���&�1*�d����OJ�.H�z�
]$�͟��̨&��!�:Ja8hL~�����;}�L~?�L��3�!��8qa�'w�Y6��#�����_Ax�F��4�������L4�e�턪&V��k��N����Alڸ�_v�ܱ�>�(���66`���@��.�9b�X}%�^?��W�QRQm�(
�$<�.!㩟�ub�h*���j�e���+���#�����\e�����E"�|�>LsJ�M�c/��.,��`I���C�xP�_�au"�X<dHB3�Kl#�"�;���՝��34�Pz9M�Ёɭ�D��Kn�-[�o����.l�$�b����[�ك�^Z���G��P�����=�z��`��M��T�JZ����N$o5:6�[O���}b_���+Ѵ��h�x�U�2����=e;��,�d�`Ög���[C��~�$I݆h �FZ�	}3y�\YfH�~��L��$N�<�#�w=�����Σ����w�p�͂<�椩�oooǦ�N��%�}��b�5]�ޯ�iSv�p=�ů�g�^{�G��}�qU�r,�4�e�d6C��T��6�uB������'D���&�E6���14�M�P�#�1��*���g����fiqĐ�-�səL�����	#���iF�S6�['tF2�p9{���c�Qݼr�V���C���x&����g�_��ݮ���\�"T3��=b�o�8˫q4���چP,�DA�a�l4�W+	\alR��#d9��������:>t@���"�Y٧zc7���jY���Qw�����8����w
Ĕ�;Q���Rz�%����V��N�(Ny��{�J�uv��!v�gl�"�w2��+?���"�/kF�nZF��>�Bg��\�ؽ�m'��ϻ�x�`�F����� j�����
�9=ة{jjs��J7-�GFe@1^8A-i�1x_��&�1-��3�5�l=KlSQL>�4<��F�����M$F,(jY�T_����G2)n�8�H��@O���#�ۀ�@|g���+ϋ�
����!nK�Y&E޸|�����>�gt����Ҟ�獻�%��J��)���g���:Z��Hϓ�i#��X��o�.i�Wu<��,������蓄�톯_2��L���[$sv�M:jz*0�\�;׵""�<>��\,E�[o�,� C=��C����aD��`�!��@"��BǏ�H�y"P7���u?�G��pM ��S�˼�e���Fq�v.Ab�cɮ.���n#��!+���6\�!�^���$&�T1ƤQ�;t�C��=C4=��+���QxRQaq�R�s���=�:'iZ���[�l�d섽�A������u(�����dMK��J2�q�1b^�9����Ȟ�#�W����Қ�:q�
�q��%��O$MM�ά��i���x� ���	z�]n��WP�U���v$����b��P �w���%w<�˗§�IZ(�+T.ݶ��v}��O��b��^MR"J�]�+क�	؊��4{ݰON�E2:v�؎�&��(�B�f�N�׹�T�[OB���H���-kB�d��\�lTo1ĥ��2MԨ��1�Mے͓���0c�o~9p� .��,�P�n$��;O822��=>�.���J�:W�3!r`/�$�#���ZS�T$*�a:[�����!��4�Oı1��/�U�\���~��.x��Ι����v�vثV������?*�Qݼ =|5�����q�kP^���ŞF5F�՗s�#���{ϫ�QG��b�J�J��-^�3���J������*D{���E��R\����)	fV<����N������b�����"$߽[����w�}~�[σ�3���?������>�?R҄�n����)���	f����[�
S,���'1�%��r��r��mr�K<��r�6�S�y���c� 4;$�8X�<��� 0&i���?Ɨ��c��|���ouu��F�ܫp��X�Q���h"�,��+���z߻Cl�)�~´J�6��!!N����9
�(Ь����8c����/�燂�V��Õ��V�E�
����bqó�\A\�j���&�����w�,2��kk���l����ϣ%�%`�d��0�����!>�����y��D'�����w���s��>���p:��M����[��Zojj��3�YGɱ�����[k)�+�ov����Q>6������4����غ��<��X���-JHS'�H����Ŝ5<uޡ.�ϲ`�D;���`ǵ�@��Ni������POn�c~"C�H�ߣ-�{xX�>��?���ċ�}%#����
��8V�g�Y��8�ÿƱ�n|���ओNY�<Ax�d0�ǟ~/��Cv�W�ܣ͒�Ęs��/}5�ӳ;�����5��[��}��nNv��F'o��ྀ̽s�y���H�Q�;=����[}����H)(���o5�!��J��H�1�ɨ�Bh���0"�Bm_%��co�����W�2
�3�g����뱬��'wubt2A"vj�q���"S�"�p������GCC�4�]�������H�h�T%��&5Ǵ�[�DL�N�\V��V��kO�ˌC�/��T��N�J.��.��|1���nCI篰�p�8�)CW���KkE�n!���`�-��Ѩ084�~���wC�"]B�L���g�j��z�2�#�ܗ)ű�w@"�u*�0���7� ����2�f��ĔS��X�j� ��{L��s-湓�D4��]9�jxz�{F0H�т$=��컛&�
p{��Đ�׈�-�rbf�<x�o�ג�'S�֪
�%xxx�ؕ~୅�>H@`�.>���"�S���Hv���a��˅b�/3؉u��u�p�}⁹�����ԥ��V��Hb�}�rk������$#AB���1O5�����n!)Kbq��xN^�Yc0_�����Z*�X���l�t��!��.���^ ����rb�˛��ݐV4s���,^���&^��o=.H�{HR�y�Z��� ���9�u�J7�у��Z�hʐ��م�"ZeV���4�d`n�Ԍ5��3b�F��S��S�� ��E*?G���P������˦��=4�Q�ԧ�:D�w������01/.[�=0:�	������II�e����i!>�ה���5��$�1E3�2��դ�V\',vf}=��+�C]���!5��!J��o����^%^��o�.|}7�)%�'�@�h:�}�=��P�~9;��_A��ԋ[x�X"�X�J�����I!9����O[����@H��,����Ѹ�L$11a����,����pd҄G��IBN���"@F*G�,�XWg�{(,��܌6�y�t���Z-	�$�+��_�u]����Q��J�af�n�b�rb����Kj���̯�f��9V�"� ����@?�À֚��Nf$�)��03Z�u���{8���&ie�=D��_��H�S��Ey�6fF���A��/6�#qw�/g������z���p�l�ĺ�:���rPkYC�@asÝ�Ƥd�hξ`�7CK���O����<j�A2��Vd72�x�&o���k˪�%h�U�S���4.�[`#��&�z��T���*¦�H�z��[@c�j<.�pXr�}�b,	��������mB)zV��.�D��{Ǆ(.�C%=8��Wn9y-�����`Z�����eZ���gosh��R�MZ��!ۀ7�Z��;�$⪞J䗳kO�f����]QPJ��C𰴴T���WI��'�$���Cq+�	11øp�>��9�<���J�-ƓP]�VA�ׂ��W�U�}N�Q'�l�h�NXeS.��"��yC�@Y�?ہq\��f?�z������ET1�.o;k1Ђ�>CY5Ը�W�;V�-�O�<F�W�31�ҿh�2����}�����w��V��Ob��^�$��I7�����Dk��ܲn��د�DVn��n���K8W�&���w�Wހ�<⽯55�Ѽn\�R�߭��O+���B(k��k���r�D�-����)B5Y���G�[i���z�O߄3�p1ڡ����E�YMm%�VTQ8b����X�B*�� ;����I����,�Be^�'z�i����l����al�#��<�.흃�b����q����
�r(�t2t�3���Ca%[G�ض}ݍ��
.!yG�u=#�]����~X)��l��.o�U׊�B�3��S�.e�H�Npr��A��$�O�/Oo�K���P���	G���=�����xd2��[��U)A����C�2��e\���À3������$z��X�:q��d�P^b��t� ��G�f���V"�d��#�ә�+ԔP�)o����K���7�k�"�A��~�zACS���$ho�3�q���.~��KjX~/M��km�E�pޣwuؤ��c�W�V\0u��� ��IؿV>��V��SCp�+��2ـ�᰺G���BmGt�V���ŧ�,��&nk/rQۍh?8�J��S8�����ʋ�9m�� ���D�~"�l��E�E,�~R�c�e�H�ץ�Շ,�ʺ<4B�.#��M��&ɻI�3����Z���v�b�b�c$	4e�eR���5��}�m���~6Ĕ���^�i_���O��Ж��fb�&7y����c�g��$z�Ľ�ޏz��`����#�ȐcCLl�5N���ࣻ����bbV1��Lz��ڲ@R��3�1s[��m9�C�k+e?Sǜۈp�OL"�A"vS��2u�ܘ�D:� ���|.$��䤱?�&�B�L��mMNX/6��2F��ߊ����@5ι/���Ǡ�qz�S`9S�C D;FS���z��&fӜi?��|�-��?�
��m.BUg�h��AB�˃=�q�]x�tG��T�����q�\�I���e��c�i�xz�lgP��|���ݫ������� ��D��s�F��>z�7��Czl����`�&N8�','g�6�"�2��wb��;�hX.z��2V�|H��������>�H�A�h��]$����cF!CL�0��G��,Ѝ��^`�Wel�w?�'N�	[f�s�0C�$�rK�� D@�|Z�i7�9��8�ϫH)�%��a����A"f���B�4r��"��Ldm�=��OT�zf�qĬ,c���}�"�ħ��~3�x�
A�,����Z�U9���.��b?��SH�E<�h���"\��8�%���.�i$#p�*�"��
�E�!�sz�ԣ��	�=���d1QO�W��#�uςl�S�=��Y<�.D2���ȰnO{a�t͖���o�-\b�    IEND�B`�PK
     ˡ�Z�v %� %� /   images/dfc5a72c-0224-4495-b3b7-0d06b4ba9157.png�PNG

   IHDR   �  �   4o�_   gAMA  ���a   	pHYs  t  t�fx  ��IDATx�ܽW�$�u&x�="R�Ң��� � r8�w��3<g���������\j��l��ZVuUwi�:32"�m����#"Ktu�dgV�3�+�+��� ;�s�����L>�gDu]��,�����(�pN��3k�s���=q.��Ϫ��(��Ѩ���W�b�ކ���1�#�����#���7�w����Zٳlͼ��\������8�=;��3�����{���4�iG���Ǆ���֦y��us]'��Q�ȟ��w�Ys�ӏ����QU2׎�8�'����$�I����9my�˙ӗ��"|�kB�@<&^�R���s�n�s��y҂��wN�u�AF�B �^�i��l-��K�|�|<g�9�7~_ǐA�/f�8��>uW��m^��}:�^G[�6#N:򗘏�#�iצ��L���d�"{��Щ����>�:��\�}��1��7_ϣ�3M�����ˣ�uH��;���g��f��:���>U��ʃ���5����;4�D(QB@����*XcWU�-"�$��$�I;����6�v��Q��i�H��׵�ӫ hkM�N��'3j
�O��t�#��3�i1K*>J�q��5�}Oqi͛۽��9AOBS�w6.��9�γ��}7��'��+�&ޯ����6zLc|��H�/l	9����u:��DY�VL���!W -�������EfN"AּT#(8	�$P0��?����>"SO����b26<|T� ������'h!(I���2��A��`L�6�fڦ(:��IS7����/��?I=#��0�h#\���e�s�̟�ָn���G]������K�[Ɨ8I*?IC���̬GA�i����5ϝ���$�4�q�l�G�S��ud�gQ���x��NڈƩ���ko��:k���$� J��|��W�������b~OZ�q5o�0f��o^���I�D��ˉ�LN�K���690
&`/G���|6��w�[F��oڶi�UA�v�t:<Fӂxv�S��9x�Π��� �D{&	�$���Lӎ.㿛��	d��Đ��l��������c"h3w~�S�cB�=�6b���s���|��^s5�ߞ_������U��gD��S��L ��,"
�q0�t�������m&A?m���J^G�'���6��c*�n/ ~���`� `���0jS�h�ű /�g�I?��c�z�^�O'\3�g`��8��qN!u$�b�5��ٴ��jy���p���K��A����������_�y��������|WW�ɐ�}5�#ab�3334;;������}a^���`��ud����a\�ᾃ�0����\|��0�3'��x}�|��x1G�M�d>��j�H^2Ԅ<�2��k�6�Y�i�{�����s�a"�Z�#�/��p�z������L���W�jiP�������P-�׆w8
��������u�kا��E^�~���R:��ƻ�a��^v"S3���iBk�g�v0'����g�;�cû�5���t��iz��7���s��9zmk�L}������4���^X�m%�AX�=:�247mjLW1�ˀ��$DKKK� L�	���XT܃����p.�86�댐���M���\0+�[
/���C㹇����=^D|��mnn��1�d�0��������j2���<�σ�Øq/!�*�_�R��}&"D�����s���>�k.k/�a�m��h�R���3�c��=s{�m����?�<���;ý�w��q~�$dd4fZ<�%���Lm���m�����Q���f�}���=z������St��m��/��,�a�Ϙ�a�y�A����*�^�1S��{��N8�*WWט����0��;v,҉�A��lm��iL�^��_����{���۷xX���FTr�y��&����,9x�F3����fy�gϞ�������ѣH�N�{�sABd�P���Dx)F`+�"��^Ԙ���P����Դi�Ba�Ef1"3��gna����`GU�H��t����hE�
�� ##�"1���m�`f�c�ά6S��i=s琋��@2A�Ə��2ѝ�%�n�������m����Fat	��^D�z���Eemo�З_\Ϟ��E+�As#	%Ҡ�S�e��pT	�f�wc�t��C�y�?~�N�:E���w�\n0u�{����i/Z��g�ӟ�_�7��?�#ݻw��l��Ah{���al��� M
��`���������r�2ݸq#L BL�X�ˈ�-�mL��N�1)������1&I/�E�lD+\����]4K�'��6Z�����Ԧ�s��1�n��m{�m��ؼ��$��Լ�	�f�����OY�w�f89_Xt�m�ߋx=����jB�}#��ϵ��H��m�Ęr04�E`�~@�����,X�ih��ph�ƖO�vM�Ϫ���[�A0W�J���lnm�O��)�?�N�8��=���k����혧Ah��?�J���9����C�x�n�Lmvi���d�+�;U�+)��U�9�3�6-�N�p��A]<ߛ�NP���&a���H%3���dcax&�M��N�y�N!�����~��c��3;Á�0^��g�Ȉ� b1͉���|C
�p?h��HL
&�e���%V�03���F�C7|�u�=�ƻ��l;�||7�	����$�R?�+n��A�����X0�8�g�54]�w�����ߌ��b�Tff�kH�Ü��&BClWPư��9}7Q���v�`FJtΠ�$C�d��Id���)��Q��!?<7�kq�:��t����1~��Û7oя�cVp8.\��tՎ��v���N2[��Çt��e�я~L�`��F�NS�V�$5��IV[���X���Qd��/�42�"Π.�p��g�S������mrf��e/��Q"�\�@�č1���c�:�� |شKK+4;3��ٳ�~.K�Ċ��g��g{{��3��s�r ��L���a���1;�p;.�&��+<Ns虆2����,�)��!4d3��@���{���k����+� ��\��v�_sMg�
�1'{{�aw���r^ΖQ��r�Ѣ�fb��mt�w&�s%�����|9:�#)����0�&~�h3|��5h���<�5	2�
B("�3��/jV�2����������Hb�%��0��`�}���w����c��PP]�9��m��I`��7o�O~���?��v�K�������셔>�̊���B��-g�b|.��A�\�j�:Z�l}}����W �%D(,�cb�Z�T�bp�����s*D��a��\a���!F��[��k���bz51��HB�����T�����MA)K�K�$���cN��5�+3?�|�yj��_��,��L8�1���a����o���<� p��;問����ح>��=x�@�kS�������H�!?Q�[��PƬ�D�DG�A����VQ�i�V�	��_��}Ȏ����;B(�{�e��h�%����$�fSթ_�Eh`���:�� ���FQY���瀆~���5�)�C��؀�7���9��_�5k��>�,�EQ+,��9+�B;��ޠT�R�E�%C����%o��%�1#U#qH8��x����B<���1��ա{�b��8���7��F�"T��� 	�s �u8���$�:�?Ɏ���L�����<�n�s�	'��+\L���kYnF!c�{��5��D�Y���\MM{�4(48���lYW	�v���oƦL-�m���5zҌ��N79?ij^��#�ae�Gd_AЛ���@��5S$O��?�@o[[����%Wv���1��mrH�T�K@XLP\]2��~�=�(������J�j%f�aB8�A�w�ܡ?��?�W^y%C,B3{�df�B"����o���_�ΟA:�x)Tq�r�.4�b�jk`j����\���5"c�i�'%6vcc��1�j���1#4!�J��
�Sۄ���J�L^��Il��\��a������r�_�����1a^�(�!�$�.s���9�S!��3�1�1k�S0�B�9ƚ�c67�l,�=k���r�Y֜�#���*j��H�f��i����L�X+�@J�K��3��wK1g�H�YhRS��w� �P���a��`Ac���vt�m����I�)Jɼ��O��Vv����?�|ς�s�b�$*#��_��A�l1����:�f�6I�`/AC���)ki�W8`�qЏXS���p��4Ư�%xJ��B�����1	 6�س�! l3�$�4[&�EjZ�P��)���1qCB���k�9ar�Z�̤�e�y��6
�LK�Ո�j؃M�4FH}c6f"EM�:]뼚!5�y2g\�7*UI�d2�k�.&��aŷ%���!��hX�9��G��}"m�����4��\L��$�TdN6Ne8��"����	s�'�+���H�/������wm��*�Z���*��j��l��:{43ۣ���`*�����ٝ��-�D����D<؇Cq(4�>&��߈�sG6B��7C�O�f(~����y�N�?����?�s����`W|�72��T��`�]xx�0�e�W�[�+(�ⁱ+��K�9i�Bc˄�c�jv�hT��+Z���W8c��өߑم΄J���G�ڨ�Ϸq��Z�BD���#����*e<��O�_2�R��W[K&����;�d��"�g��-��V�LJ�Ț�����8w�C�""
R�K��
^Oj;�i��k.���1������sd������o� 5�1)gB�Ɯރ�+��&O��97�|
`K��<��*@��6�[��ՕeZ^Z`��u��9���O�)<�#A���f�뾿wH���^_���p_���<
~���?�!kl6/�,��8����/��/�Af^Bɰ�B \73S��|D�D��NGO9sL��A�^��#mrĎ����V���1�}&�$�>���$�4��M�u�U�iXA���0���C.hL��]cZd���NL�9e�(d�u\c�G�l�1;H�e��;�� ���ٖ)F���&(��"��J�mM񷥲&b� ��4Q���1�35oҎbK��,�#͘J_ka׼�o�]�.mBuY���%�rUOH��>����<�]�f�\3sA#s��	f�לq���gf혥����ԋ�Q{A���cC� l�%�-���َU��`w���O�Q]�r38>�P&�}��ٟ��l��{��ށ�	�����O��O��o�͆���d���=ZX�p؀�:V�
I��r��c��|�vw�s�Y{�4��-��Q�9�N��o'�9{��B�j0f"f�S�bly��p�0��Ò�-Lgğs�ɳ����E�����6�� �g���⏅
����4��)4�,�d�R�3{8��1)s�WM�[�ɡ��#&2��.�$��l}�Q�ƙ'�䚓��Ȕ�2����|�/%�%98�BP�24 "_�Z*Nq���+8.y]Z\�?s�?f�G�h> ���9f���Y���i�a��A�ƃ��;�{Ro�����=ۛc�~��m	48,l6���K���:}�{ߓM|x��e���/i��cL50���6�'��:��g�(�q����&���j����olÉ]��xkk�67�i;0w�`�/=1
5^Bzіώ���C�\�ҋlӀg��6?KpV�M>���9a�:J�����{�m���k�����&'LP�؅a���M�O�'16_ո�����T�H|�Ck�i�e�gZ�\^VkH�|*v��T6�Is�S�
�T�o�v�k��S�@긃Pr	IXA�8�F�Ԏ=���.,q?�֏��3�h9����D+++A�.��fů�|��8�H����t/�<z��dS�5��ܦ��]�s�^���"����/P� ��?D<������
���IR����a@H^G�0o *� �`C��|��0����6u��N��k����}��!=z��Z�2AI��Ha��k@o�w�zǈ,?rh�@�3��<�J�H|:7�ؠ��L�I�?3���{s$�PҊMM;}~�}�j�gc�ߖ7��[b:�_K�G�˽�I�`���i��\��k�WEG3ޝ���H�2�G��.��nF1
'	V%~:�)�ufiq>0����?{�.^�D�.�L��Y�?1�D|<(��װd�%
�fz��!p�=|Lׯߠk׮�bfn�5�^��	 t��D� % �ol<Z{��MRC�6o�������a't9�P�K3���2������I:q�4�<y�V׎���T��=������ݻt������˟GHa�'�+<ޢ���3q��i�3J���w�_.}��F���M�|$���*��|�Z���M�C�~�(��S>�����<��hk�'��=�濛±��ڂ6��0��Yd��ؗ��k��B�����iui�N�<M���*�=���-�}\:M�J����,�d�t�f�sj�y�̦����C;�{A8�qt�m]����]Z%��JA�H��Df'��[\�吖آ�Zsa�Ǐ�t�b�Jc�v�2�׉Hm�������j�S�N��������$SE�N��3���r��@[�N���{Oex:����d���yԹ���Oz֤�?k+�i��Y�_��32Ƃ�<���c��t���_�3g�2��3�	��ȇhXˑ�g�$<����|Ĵ]vXS��R���/�5�G^u�rd������E�������ÍVV��ܹt��%:{�|��9?6XZ_��ٶ���	�����L;�t�K�C��C��ˡ_*]|��_�0/'����|�3���f>�ϙ�{���6���T���I��u<Ǔ���q�m��*~���i�3\3l�3��k�qN6h�|2���^��`67�Z .Z�Sv�`�NP�c��I��L���-�/���8A�'{��yz�YK�~��Z�Cˢ��$C5�R8.�x��W9w��}�}�6V��;��Do��	�MjWz�1��۟M�0yҽ���h��~O��G��qL���&T���b�7٧����k���R��-_�7���(8����;��En���qS�Sf�+O7M'梨ܸ���	�������=x���`l�� 3�k|�A���M5�a�� !�aC�18���t� �φ�,󄫑d�!@��1(fgI!Z�N�p0�.8�[���nllĪ�锧_&(����d������(8�<ǋ��ߤv<j�^�8�t���j;��c��x�zos�����89�ĉ���#�u�p����tE�^��-��҆�Z�����}��I�z�p�x��f���G�_HH���s��ו$�d�}��iz�������iqa�=wR�%UQ��oW%UM&pD��X$�#�)�h� ���ʚN�L���Y��QǓ�I��E<��}'�w�t��&�����<�E��v�	�R�6�D����9�y%��6v�[��fC��r9h�\�"Ğ�|8�[��Yo�/��:�����\���J'��_�'�>��:ƨ9}���

:і�!�4���ҹK��g�����A������R��R<�5-���`�R��(�P�T���bk�?fn���-�������ֆ�I�T��s�$��W��Q&A�ؓ��i�Ëd����!x)��F���Ӿ�|R�����=���C��l�7��e�u%	<������a��6��=���+�t<@q<ρd��R/���x�Dl��)أ7~`[F`�_�����Ξ0l��q*�đS��Uk)�
'�fHx�Qf�@��WGY;����ê�}a>m��3ӈeѶ%�Q����Ӯ�����e�?�ьd�~ֱ���g��<�k,��������Zz���#AAK�J��3���� ������<���aufJqcB.��vt���4���nM<�*�=4���2�ۤ��o6\�ki�8���Z8�"�'����(�/cz��2�0Phj��9�-I)�7 ��c	�yŧ���"��񋚶���Q�Q�ݶ9�ss��{B�ٙ���>�g=��Qp����W#S7�WϢş%z�w�d*���l�«L��g!(��Z�Dt���+X�I��㢑�1��yZ��4�T�Ǌ�*N���:����ģd�cنMGw>��rK��4�Ǚ�MW9���Z��	N���ؙ
"��i��R�б��2p<�|��B�"_&�{�ϟ�G8�&	�g�x-�4��/�x�7�6��ay���Χ�x6v�ӌ+ާ5�xN�k_��Ԯn*����`ȶ�������\?�1	ɒ٘�b^���+,����.v�#�pY��4$G�B�K�2�rO��6���Dp�bV��T
�-���5c�k����� >��؎Ҟ�)�s;��I�v��M=�x�D������;�ߤ��Y�����sl{ӟe<�4��%�dГi:�Nv�=rO8��:�B�:}�K�g�.�����㔾��$E��>u��z��b���Ԫ��YWQ���������"W�+��m��K�ћ�505��mi<E�ap�$����7"<�%�:0쓎'������4����q�W�c�3���y��8�;+�4�0�FK�~x�J\C_�a����k-Le}܊"ݓ5sm=�SxK�w@GĨ!Hr����	���#Kvw�?H>G�כ�ݵi���ʖ�V�	�֥KH5��
Ig�1X��/r��=�1��e���U=��Bt����:�b�y�e[�>K8o���}�����"+�.)��f�g?ڠ�@���*Ced^ږ:䛂-��g�#�S�S(/��eX�IZ�웷ǲ#�y��ҒB��8�$�е��u:���q@VO�,7L/*��	��VȔAx��ɵm�ۍ�*h�<��$h���_ԑ����ȓ��,��x�7o^��_U�Q�3+:���n\��[9��l�c�^'V��u�{N�c�����#o���ȍ^�x�k��r����Io�Z��{���O�C���9g,�AZ�.*���G�7�=�*K��[�n����������E�ߍb�_��(=���G��q��rM�<��{�B���v�a�.�r����|�9]���,�L�V�e(L�v��C���t�Ո�������֭����E,��&��b����ͭ�xww�cսN7��	��-��f���&/����>4�R��nv4e�8�����m;u�R��R�������?��~V��&�ǥN��� ���=��s��:��PfR{��J���al��j-��Hi�w����4��N)�DUv�@��ǟ|��$�ZJ�����i��Û��@ܚ�_���8��ˡ4��:�	��A+���A̜cR�"�¨������I+�}L��SH� �yۋ�|Q/V <mH�O�_��~�{�����i�}�����9�4��q���3���P��O0G��(��v^������Wiie�Μ>#�<�s*m�U(����f�J�f8*�D{j�{?~���߸A�Q��-�O4qEڌ�z����������q�������ϻP>
7���֤�����9'�̚�;�dl�#�=�G���	[a!>��� +�K�i�2��Xŝ6d/�����Xi��g9��1�,�L�{�uf��x�$��}R:m�4���!G;�r�|�â$��<g{�W9^��iK_�3.9K��8����Í��A)��r��;ߪ�왳�F�6���]8����«��0������� 沵�M��s�����>�z���R��Qڧؿ���ec�3�����p`�40w~�>��r)��a�^��T��ˊ1�x�hD�k��ݾu��{�����[,��%�Vr�ie'�B�(J��*�w�(���<��I�3K�)��U=ޓ���\?!	�$��d��~�����
��y	e���&��yh7W���xr�J��$R4-��;�A|��}gϞ���G�%��ҥ];���Ƴ�n������_��~����>���p_��h&쌭���M͝?=�vJٓ���ƃn߹C�\z�V���͢�'H��&X�.0���O�\�B_~y����P�.�I�mm�mf�1xg����h����:��Ey��9@q�ͦ��4EL��J�U1`;mV�AOL��*G�O�!��������ܦ���v�t��sC���V� �(l�b�m�$m�R�*�ƈ�{ءO����jO�:)>Vdn�Z���36��իt��K��a-�p��	*������$�n�L9p�]����Ï�� ��ͳ�3�I��R����sc�Wv<+qOCO{�gy^�ަ�������Qٳ��_0��*6�����}񇙎�l�|�m����=�i����v�^}�e�9���c���H=����F/�l[<d�>���a�ʕ+w�n�P��䙄��yI,��7]���(�x��o�ɓ'žƎ��N�9��Rv�`�=��n`�k_\���������������}�������X���j���{L3	�
C���qhn�N��1G�����<O:����$�<�se����7��)A��}��8�=�~�I�ݻ��3��4v�XZ^�X67�e�Sl�s�������h�D����	G'��18�C9����w��և��.]�D�ǎq�*H\�{�%����v�`��0p1�e�Ηu���[<�{�K<������<�G��_�y�̔��� 6@@d��F�����[��}��{�"�'9��K��y3�|]�.}�B��
�>��8�r�*�(0%�1ϰ��;yB�ёb� ��'`z5��6�N�_G��:����8����a��������ӧ�:k=��. �B ���-0lH"��1X8�j]۾q7�nb]M�;��%���O"�g��#��̈́��������� C���)����.G;|�M<o�s�"�l1���φr��\ZJN�H�K�KqC��T%�,�w��N*�,T.��yH�ҝj����"0a>���-�\-��y�ݿ��m����u�v<L���0h���]v�I&L�N	ȳ��$��{�3��6��O6b�~R�QcOe��XyN������g='��S�`'1Jk]e��|9�!��g_�4n�G�"I���!@�('水f���L������Q��� &�����tՈvt����ۜ�71<0�aTi�+�#�0.~��O+�Pc0l�F&ǃL@��d�<��6���D:�fj�
�������$�2��_���fRcL���]`[b#B+�u������<&��q{�o`x�#�cȑ��
�'�wLJI�)�K����bv��=�  \�=�]BNxO��ҝ&�����mn�!o6�a�"�l����{_9u��.C���8Te,�Q�w�����WDY��x�S���-�ޖ�u���W����x8�vޓ4ǋd � ���%ajBh	Gc��,��������(��~���i�?Y"O�3�uJ�c��[���+�ޕ�m.7"<\�ߨ��Ad�y�\���/�۸.v6��M-�o����zv�����)�HHLq�}�f޺ū��7tʶI;&��E �0	 v�1��GO��q&�G��_�<G�u��dǒ����c���/��o'�L�	gc���i�6֣�Ѵ�6��3��Y�Iΰ�ì��L3*-�(��5x������cz�!/)7�bz�ܧ`f�`��u��Q*����3Ǚ)fS��n`��{�ke�I��t�b�هS�n3䒜�M����o@s�'/}B���xB����4Ȥ� G1ۋ��㩼�nʿ_��M���=�ys�1��^{�{����/��u�kchw0!�|Q�2J^�H>jwf
��-�w�1^�2kjH<�v��O����g������Q(�M��s&B��%�RW��b=��[M*�6x���$�U�-�a����i�dN��D癝�����5��=�Z�Ip:/�M_>��&|�)��m"��`h��Z�Ņ:�p�ұckt��q���.mnm��8�U���acg���ZC�y&T-qY��H8k%�1�$��{U>a�O���L���إr�1��l�9��o^KO&�o&��$��t�v�9���6��c�}H�(�|�<��fH����?ICRԞ`N��#O�&���}z��7[Fc�(����� ����߅�Y~ElH踪��h%�y�Ƽn�#��ӜZ g��δ���w����.bt��Ȁ��~�';5I(t2���Ovt�����b�3Mv�g��1=o(jZy^F�6���h{�ӳ������|Ӷ�܊��%���2B�W�\��AC�X�F�P�m������\��6�D��.C�2ܯO;��Q��~[����^��7Զ˓'�r��d�(������!�xO�s\�!�'^���)8�5�� KHr�3��q�U���
GГ�t�1.<<=i
��1G���Zu�-�u2�0�ӌ�h2�v�C�������m�n����p���0hf4N�t�"�0�A�g්C]���_8v�A��eh�����aMs�\�%a��-ϟmZ��
`|�6D�Dff{,U��Tw�D�y�{�"i�����&!j?�Ȝ��E�5c��˽��Y�E���x��-f��}���fs��y	5M�9��Gs'=�y��x��w�{���H���S� /`�t��(� S�3�n`�C�-�|��'���7(4�y�kkk�5evvF�w�]Wx�WF�={ a�A���S|c�˒D�G�>D[��Օ !��DI-���۹�8$���ĥ����͆��x16j"0�&@���Q����S�T�9��U��N
[%��4I3dk6Y��2�0٧p����cn֚RJ��#y�&F5.u�����S��#H�]#e<c���a�SC�	�[o�E����|.R���6�&�P1��Ӳi�1^�^{�e��Khay)(���9gz������5
3Y3H���-kHh��R)hyy�N�<�^<0U� )�H'E�ۡz�+��k�S�J�g�dKO4mk�����j]��;���{��8KYbkk��l?I��>��(�M��G�4O��=œ�9��֢6�42�j.�5.��F,;���#z��ց�V4o}�#��i�){��kD/��yY`sK ��{�׌Bt�!�5�;U]xAp�<��������徥z�����������Z���:�Zc[��/�4�d�I/o�Ϸ����;�ý�{�oܧ���W^y������zV`9��b����Rާ��s�?ds���t��)z��<�H�w�mm> ��O;�b���
���PYȞ=KK,m�� Q���[;4?w�]F9;�KFjU�G�s�2.c|@�
�C�Y��aǜ�c轄v0�c*�ĖC��D�=�y���2����ۡ6�:{iS��ӄ�!C�os�3� �8�MИ�w�S�_�ϡi'{睷��>r��P���s<#�����ټg�Gq^̠.1]�Ƙ���aG䛏�1ˮ��YZY^ �Va����0�3��s^R;��Y��� l���8:q|9��,�Ǜ��xgDF���h��8���0�=>k6�N��fh�b�l��Qжǹ���g�i�`��|�U��?�!oE{�˛�]�cow��p�����,����#n\�J��N����YA`/�����6���S���7;����͜ek�+ap���p��Ժw���Hq��߻O��|���"x�3���<��-��� ��F/2h�X�IPe���)�4�%����A� 2�ԗ�I�s��Ƞ�Ӛ枦kk3'Hg��uy߱���W'�l/I<�ɞ��	QX>�~��dZ�/���e���E�ZT���Ζ2�&Ӧq�iT���ixs�Ւ�Y3fT�s�i�ئ<��F������^'�Z�3����/4��g��&K�u��*�c������7�x�~��ߦ���ho�>��*���?B�ϨN����'�� ]�=�]lm��[��k�MŔ>��ݛaņ}��X?}�'�������uG�n�
FP��"�\/(�����4��GVYp_H�G�V�MNg�v���2�/W���'����Xl��,H���`/c^8�,�܇̘(�"[��H���%I�[Xbÿ�=�01�߽{�sd��|�A����?KO��#�UK��ڧ�QG�tj-�r~Dx�tl�R���M#/1���Y�<�n����Ѥ���s3�*�&{n���ތ��� H�޽C��/��'�~ƍ+���:G,-��}Ɵ�����͜"[w�L#	G&��Q`
 ���91t�}��YZ_CnFĹ���Fph�Q{ij�9���������W��ߠ��N".�9s�����qD��>��(�p��.�5�7a�zZ_Wj���j�Xpd>������|�Y�� /��*7�X���}��.�`��ᮣh��i�eN�ij�ϖڀ病D�����~��8ʸTL�	�b����q0�� a�C��ث�F�}���Z]�x!��� �Nh+�������;��=�H
kz6�7�/�:]|'ۚ�����D�� �I���Pܥ���;��g7���%4 �3�vk���9�G�?D�B��l��xn�N�e����a���
�-Q�
���JubQ�R~�s�s�T�t[�xJ`:�|�T�ՙ ��Fu�5�[{�ˆ�f籧�
uz;䆣|u���#-h�+���ß��筕ц��zҨR��X>6S��_H��'9��+�dh��F��1}���ܓ��ٳ�i��ÝL�Z���%�K�f-�+�hU�\�)e������p����JLʂ@��j�v�h#���/hg@d�Q[e	^
��;8<�=���̦^DS�ހ�-������[?ήz��=~������nۑ6����+�p�l���6]Z:�~��j3�|N�}��L��*�mvn��N;��kT�?s���*�����D��MaN�xge6���k`��FO�K˼����G�F�ޓL�Z|L͹4�F �D�)�l� x}u��@>"*TA��q����x*�l�~w��.�q(�<4��^o�Y��a�y��������"�9*�-��盽�ƚP#����C�]�t!0�Ifj02ƺ��E[pxqٱ �[N�)��w7@��  ����8)P�^P�{�R��]��	�ql�ێu-Ie����[L]3vw%����C�)�����v��	49��A:#Lv��u��]�����8��=�cL�+�����^	6"�䱠��w��B�t+��0&ok����M?]{��9���5�O�
3Z6^[=$ܴ��
���
��F�?8�~�6 ��Z��O�Cֺb��z��9�<�fQ���Pd+�E�������úۅM��t���~��3f:ʂ6@kq:޲i$����$��7�ؠ������������];o޸E�[���|��ܨ�}�0
E'<^k����r���#��6զ�zt	ku�~�^{�F��|��Ѓ��b���fk�cʨ�aG���Lg��Η,�e��`gc��@/��x׀��r��b���2d���6��j����^@����&=v��x�lr�ra9W��������`[���_ҭ۷��p���t�ӄ}�$++����N�
��	�a�Xi�2E1��&�U���h��9�Ĉ��z�N�=Ƶ}�Y>�F��M[;�g8�6ܦ+���=�gϞ���Y����`�l�im�!��K��(@����q�t_�c�v��A�}��Gt��ɴ�}�v\�`Ĵ��GL��B�5�"��I}�q@�������]�u��z�FD3L�B�Z�}��-�j<_��k��+��c�G�I ��`�E�����F��Mp�þ�����857DU���`���-�0���U���M���ž�&!2�H����Z�j�P�g$�t���a����0�0�/�����a�m ��|����Bb! 9 I�WV8y��o�M����=�t��	z�z��7B,����T�ѿݫ��8\�H�Y�S���nG3c���P]"p�����s(
!���(�fL|���t�l\�5��L�i��"u �y� 0��T���g��ٳgiv�Ú��טa��Bh����C��A;U�QVhҼ�^��9D�)\��6ӷ������0�:�%+���@ln�b���$�;��y~��d.3���	�.�ܥ�ΩeL��~Ќ
+��t�����k�q��6�s���]24ɧ�P)i}}���0����̵]p�kڟ���ᝁ���=����'�۝�{CB~#t�1��䖐o/��3���ƍ�t7Hw|���6+ඔQ�`�+ī�ÆU��w��!��eC3��74-�<��������a?�nG6 ��oM<pY#';ܽw����w����#^.�@V��h�u4�ԣ۶�G��*:��eh5Eϱ�'fv�U�؀��b�6��Έ*��	��ԕ΢G�����YA�� �Qҏ���su���k���:�|����{ֻ�j����E=�9�x����=��Z[�H��fii�����c�(��y���n,x˙�����Zcb�{�}�X����P`�Λ鰿�
o����&��.��� �ZT>�;�E8:�g����"(8&;Cb�)�q�����~����9௺}�}����G"���(���^P��A�pl	_�����4��cor	�x��cE%x�k~"k�\�Î[�Ap�@*�f�ֲ��q�'b�K4���l%0���aư����Ǉ~�V���~��Z��m2:�D���(�˞��D�~��v�P�B<���sgGl[@Bc\��
�BI�4u��j��|�C
��'%f���;�0�7XJ�][�Y��=8jJ|��3��4��v�L@��V6��+%�]~x���ݠ��g���r��:c�����Pٷ�bmi�`m���F��K�����wUz(t�1�DV	����^����A+�\v�
τ���g���*����0���������>��
eG:���M�.��1��8R��#]E�Z��يHm�@
)���'�D;:AR�� ,�Y޸~����i!h��z%�����W����56��?`'0֓��<S�"��a��E^��#�@�Ñ�^�BTY��;��K�Ea'���e�N�F���SrA���9�����q��0Y|�{Ab��M��R��]��ms1x�	?HD�L��a���V�h`����BN.w�4aH�L]U����	qɋ�"Jj�zcn5�~������+�ؘ1'&jt���36��嘗J���x,�J�	�AQˎ�"D
fj|�ds�XN0��2���Ƥ��6�0}�l�%yn�Ì��kF���^1��+���J�X��9sʚl�ZWu~$�p��F|c|X���[n�S�6�$9���S!%����@x�7����b����v��3� ��ExF�+=�`
B�Ai���vX/��LF�ͫ�x;���ߧ/���c��\+2B�yss7��}vb�y�n���q�Q`��!��]:�?���tO�@֐�a�'�������0̻cV$<���o�r�BAR��D�8!�<��	�H�l�~��qz��7�&���� ���s_�JCk ��! ր=��9��f'y�7�z9�䥱��ivi�.�t�^��{�ٞ�[�j���j�����
}x���-ș�˅f'�\;+�~�����L�4�7X4oMf3˵u��.]4���ƩG��-���L�y)M��F�;�`}TzSc��au,ĺ���!�nɗp�^�C!cᐾK�G�<Tu������L��
h�������kF�m�n�Vd��u]�#��Y-ξB�_o�� �d��&�Q�y���1O�:�s]]^�?���:��	�l`4�j<��Ń�$d&sbތ�R#����0O�67H+�����KD�Jv~����Q�#�렀:���l�2�g�X'}Ui[*�+DOs7:���d�jnA�Т���&�[�m�����5��c�K�8KK+��;�Az�/F�6�����s�9���N��"��N�Gb�~xY}N���0��+���@A��:}��x�]�t�����?�� ^��I���=���jQ{�T��DMG�9D�d�=�]�Z\<��x�����N~6%b��"�V��LM��I
cl2a@���ί�o�WA��C�5�$��̠��!�f1tRg�!�! _;?,�(p\����Jp�J�y�@��f��Ϥ�O�ϋ�rd�g�ꂬ�(cY��*H3�!£���M��P�����o�n�s�l�dN��%� �ˠ�vf�r͢�v9b��:.����V ��d�1�{�Vں�\�i�=ו�F����t�LI��u��#s��� HS�c�h�b� &9��G#�Ы����D�e�`�cØG��Sg8��]^{M�C �'���6���]l�V������Ȩ�
�IQ��e�Y������|饠�����S#`
<�P �
��f^CMN�DR1$R�473|-��>uj2��C�Bg���xD#�$Fh�yi�k߂*F��U�����JLe	q���J��kA��B��P�o��a��gy&��*��(˓���L�D��f�V��׼�c�ή�UT��@P���TH"�Hމ��*��)��\k�cL�����Y�4�M��C������L��#�����L�@��� o#�O.$-��������Y��@AbgKbH�6t�?�c���:��)�AI�y�l*o�P�M��f����M2��殗F>r�Wx\G�o�]D" ��'��FB���^V�"@���߼y��I�iE�4�E�M�t�!\��������hue�Ο9A��Vh��a=� �����tlm���;4O�+�,�6Q`��F��>J��2�>iC2	�J��
����ؖ��H�_B���,GI��͞l�4���x�(J�|R�f�1�p�ص���J*�i½�k���wd�g$�C�!�M9�Sux[$���=+,�.l|:�B��<�6�!
��3!pZ	Va�x�SqI
'�}���v�-Xų��j�Sp��z@����_	/�����k�~��<zD?���w�G�K���.����f�.y���uV�*�(���;qp�(4�_A��	_��0���У�~���"����-������x�#S�����N�fX�Nb�d��Eb}�e����G?�w�.C?OO�a'����7�AWF;��{K����Q��>��t�����}�^}�%��;�[���M_���\�H�����:���Ck�1A*��^ڤ�%'�ʅ8*]<�)#<򈼩�>B�,�/
ъ�k��q��զv��(/j�����Ǭ+tVDlE&NmJR�*03g�AjpW�W�����>C���<��کf,�n��D�Uyk^�Zږ��زe��y��0b��'mm�S<����R���E >/�%����r��'N�B��_�F��s�74�p�����t��3A����[Ac��Hx91��A�&�W���{��
����aUsH��1���֑�<�B`�ݻ�Bm�j���Mc�m6�<]�mN�;qRt��Ƚ�8*m�*���/�;n��� �����$��yP#�/�jC!��z����4�Exk�~i~�����~��������!���I[0Yq��Z�����>�ʘR�`�,>k�O&K)bG���߽y���f���(B�m�ZmF�	s���.%��ڤ:Ha����'�����������ga fm<��
-�ڗ-��U聴�Yڥ4F�N}2�x������-n�gךc��̋)��Zr5_`2�r��� #��(�+�Y�3��$��-zkN��,.m���
�9{�~��o���������+��76���s]s]K�`��~��tl���޽�n߹CkkǸ����wysI��P�3�$?��F���������M]�!�g{�P��H���a���(�ʒ��/�:+����e��/��S��
S�F�#-��D�v1�.<���ZXZ`�c��a�Dl���Uz�������߹�i��{��wޤ�Z��y9֧}�XR���I�Q�1�ѫ3�B��q1�W��d�L����";2����i��,'��ih
�^��\t�Ʊ<��W{����l�C3�V2M�2ݒ=���4#	L��+\�:��0/�T3��J��*�-�y�L�8S'�ek�vda�8;�4_�f�~C��gnv��2�y���/N�t�1f���3�9;i�o��:����s�!�۷n&��k=0�[o�M��?�:�<���ݻ���<��̬?��?	�o*�.�y��S��%6�������d�����f�da��d�mB¡^�Si�y!kv�s5�8$�*+x���������a?�P�iuk�J��;L0�Ks��?�>�;�_2HZX��҉�e��}cm�.�K��x`�}.����lj�?U%̍��Ü��l?`37�H8�>2ite�
c��vI
ˍ�5�1s�TC%&��m��1Jm�ܲ��&	eg��[����:��C�:�s-�b�V�ND3ŒG;��s1D$f]���Z�]�9ڹ������+����[��(���֍�8/u������b^�*F��.���x�"&�NR���ufD+����8���dd�!f�8;����	5#qb���k����g�fF��'�^a�q��K�_~�8{�QO�4N�A�:���p+y�j�L��xC�"=;˰z~yN��M���0!�\�Vƾ�Z���-�B�ҙ�H5�g��{�$�i��E���=q���
ٗw�u��ɩ!�V<Zuqq�.^�@/�|I�ک��PV7��'���`�nݸJ��!�%��C~y����Wj�U1s��%�b�)����wl�g����O���4�Q�S甁J%t�k1Rt���ڐ2��М����c9" o^a����䝪P��q��[�6_Y6F�n~i"���djj���#��zlL�'�#�p.-�C���/��|潏�Rj�#Yu�1�B��:D#���q��-{ԝ����E�AG&�;D���O���l����>u��̠T�Tsi�]�5z,0�_��%�Z��tG����|ձ�Fi�!�	f��M��~",fg%�CRx6F�)v�ԯ�9:
���k�gK#Ț��G���%�f�ig $�s:��T_K�!���eN� Q ��_jqzt8M���"8#���Ϭ&�;b����a�!+K[^]fFF�&�f��s�1�� �LP%ۼ�	-]dB�N*����	�:e.�j:>�ؙ%�,��=�9L�$	�[칌Z�k�ό})�zga&���(j�R�?�sMH�9b�n�D�Hdv�Z1c3��dk�i����!ʄ�S!���(y||d�C�}��|�fu��%'�P�>���ؗ��
K��%K�ӓ���0H�>(����>�!�y�����
��Y����)�`J�ڭ���ܢ�O?�y�����w�É)����wv8aD6 ���j�:6��'��gA4jK��#��A��0g�5aM-Z��^cLj5��kk�ֈ�5+���pL�vCWj��3g���
���K��E'$W��;I}�kcs���V���d�����h1��`��x+Ѳ�7�攱Kc �e��{Ɛ*��{+��җ�<C4V"�[��� R�����B�A�45��h�k��SMe��,熭�Fќ�άm`��0a��	)R�'L+�I҉ٹd+��/r��3ek]gk�>�퍭g[m�B�uL�sJ��%�ӡ��� �Q���흺�Y����!��~0��q�`@=t�4��D|�!s6.~���	N��z�
���{����5�'\ӓa��~��:wű���K��ó��B�w�o�'q�~B��݁��bv�F�44'5�s�F�q"��ށ�w�lms�^h%Vx�Ћ
�|H��/qWKTy��đ��Š��q�}�{��A�"�$qf}K�L}��	��A������Ew�V�iN� io�n�l��'�9��]��C��Z�J�u볦 �̟T�΍D�\�;n�#^k�t��o��+���������1Sr���S߃vɱ�I����Q�H�#1�H���xL�4�`p��ӂ�"�;�
�@C�5�zp([ߠ����+4�`�l���A���/��CO{����!�M)�A�
ҡ�&��;�	��=�u!��>��N�>�~�{gɼ;�o��m;�(�����
�p�<@:Q,U4k,Iu�Զu&$�ԩ����K���9�f40w�L�Ia��Be_
7�ߝ?.f6,�g�p����R�*/C�z��x!�4��(�DB<׌�lsE���W售
�u��޾A���=�A7H�.._;~��+��&Q����C�9��Mqa�����R�Ѵ�Y�L�3�i������F��5m��Wf� �pФX�#_���y��sc��E�k����x�6�>�n���؆,2s%j�N^�i�
M�^��/��2�ZD�?z��{�ߘ�M3 vT%�yc�p��s!+\Ouj_���/ӛo�I/^����8��yϝ;�]Ty۝j*�9��G��x��C�����c�˨J~"TJ�	oZ	4׏o�yQ�v
n�~l�cn�A�A������'�l�$��!mnls���G�R@�'@G<���0*`p�{�G׮]�{½�x9��g�]��E��\�G�Ѱ_I�h�Ҵ���Zc�0�[�(�oh��9q	��ꥷ�h�!"�IT '����R�%��X�o�D��O�a���Z0�o.<��$[z���&�	C�I@&P\ChJJwq���d���ke�L��0��?�t�k��FqE���-Eө�A�67f���`��全AA'H0��C�`ɉ"�@�\�I�2���;����B?�����Ӽ��a�t9������;�����!��x��
�dkKBW��!l��2?����	(�q)P����׶ �ƃ���� ��xPW��������$�q5zxz��A�+����@t���AcC*A��N�]J��3�ѯ\��L�Eb��p�=��%-��+�"�-�� 	Ɓ*�~��<��0�����
�hޚ�V�A]t{y�)�m�6�8�Ǒ��8טYg�.t�tHm��t��Dl��$&kھ��d7����!���$$ﭙmN��_car�m��8��&�貙C�MX��yӚ��衷�Z�h)vm��`�� ���-;}��)�����z��/p�3|�pH�oޣ��{z$��G 1S�F�)�4�|L���[����ꫯ��ٖ`Vd=�8)I����мm|����Qxl~@k���	͉b�Z��R�,ZF��ɫ��*Mlr��$��y�z#��/Z�Q�����2sC���_^�T �<w���4�.�,"� iF#46�Y���Cw�F4�,��x�Ξ:N�Kab�C����p�b��c3a�k0Rbؗ�`tnE"0qSڮ����p�f̙���{�#��>ښ�)��m^���3��+�M�g@�c�!k������Q���c^�y�v�)I�"�GJ�0�S�Χ�`�gg�Y"���Y8���e�^��}��Í��9�C��<s�]��+k��
zgk�  J��J*�� Þ�A����G�S'���>���xDu �m�-�l,nKO{��Y;��T=�jȒ�W�xM�Q �${�l�Ǩ_J�}_��e�a�{k{��6�8�&9�53����Y�B�� �--Y5�űfj�т���4��q��I:w��~?~��s��y1��;�4N��i�NX�¨;#�H.�p3��:gFy�d���2��7�Ԝ�����8c�
���M����k��J�U>��}ʄ�Gk
�L�8�|FꄬTX�ZC���gW��`��l��t����k���i��;�lxRcm��zM-��8���SJN�r��
!��	4����]���/ѽ��l�P_�%�%W޾}�������?����=�;t��Mz�]�J���UJ��*�A��L�Aլ�f�y6eAqrG�
%�fx�*T�F.*f�a0���!�*x`�����s�ݝ=�ؐl���D\��E���b�.@q�8��,nPo(@�EHMHJ8�҅��#�m�	�Ǐ��5��c�WJ�0h�2�<�]*���Z�2g��d�B�k�f������]ɮsEM�}C"{��y�e&0Syk�j�])Zv*��%A��f3;����y�14����(��U80��K5sp���s�f�1�Ezn]I��"�2��g�oE72*~V��jh�^P|)�r޵�v;��)Lh�V�q���'O���U�u�A`�-��1��������N�#�/����V����n��w�shp�Ƞ_����,��a�h����;��ܚ�����W8���{���J��PБ�0H���=z������-v3��7����G�qnm$ms�y��1��`g ���o��oq��G}ȎR�	� !@���[��H�/�T�T��A�t�`�?$(�Lt�%ע.ɍ����G�x47d�k���:s�(A���9c�n�69�"�F+4�o-y����v#��ހ��h�Y���~oߒ}JM�$�ʩ"��8 �V��}Zi�rF&@:7��ٝy��^�w�&��FTDf���i鱷�UV�'!I 8��t{�y�Y�#"��ۧn��aW��{��>�¢�3�~���z��׎�~! �mM��?��
�j���hbβkf����ís�Y�@��Ѡ�ż�OJv`)L���s���E!M$�d�o<�ͭm��=I>��n�x�X �#�d}� �~����v<׮}Ρ.�'jS��Eo��^{�[Ȃ|G�>Wf�8�F��M:<أ�G��/��i���ى���,�{Ae�d�,[�1���_"�D�9�-P�p^!&/vzp��s�]g�WB5D����^������1Kǡe�>=Z��3w;���p���DcTy�s�)s�5�-(B�{��5��k��>c��ؖ|�(XUas+if�n��i��T���$
ِ����C��A��ɵ �=/.�R;eE�(PQ�7~�h ���Tg��7|��o��|�mz��X@a� ٞ�X�"��ڼ�3qJ<}�w���[`O<�L�g��j0/�D+R�`��$SC���1OdЗ����t;��H>�<<ԅ�j5���DgϞ�49�:�Â��c��V�Î��t�p��>"4N��͛�����-�D�w4+�HB��Q{���ūr�T�Ax���(���g-?ٴ�,�d��P�����iF�m�N�g�u����J�Vܗl��6�<�Ӎ;���"��q�:���p�9�P���4S�i�:3�-6����_ku������f4�"Ap����9�3�̬�;[�Bg�i�c��5��g#u�%�̲�׮iqz�#v��JF����s�@�;��AQiYe����%������e�.�[憈.dd�Ibu�23����
��;�y�G{�a����$)��=� ���g�W_�æ ���/>ଲ˗/3�s��JPl�JH��6�m+�(��K)9>7ː�(d���5�.#V�ߎ���;����(wT�����M��iWO��!fD>�+���!��,�
�9���sa#��<��О�$���3Ɏ�'?a}�w���|��@JQ��b/[!H���六Y_�">��=�n��y��o�ClS����{��QA{ػ=���.k�J��?`�/ =:h�S�ORgA�/^��i9���!7M@�+�E�y86c���7e��hq���]mީT�-�����$������^x�@�5�Z/�A�~���	���?���ܾ���l�#q4x�9��ˮ,�xw%�UE��C-[둄Ђ�fۦ���,$7� �Gu�|`<D�$�I+�����"˱�]�>o:��ᰆ������Z����]f1O�"�%ڨ�O-�����dS�ǘϡ���a�!69峵R�r-���$����P�49�O��hC�B��l��H��Ɓ5�'���2gvac��w��^@�wPٝ�[w�qX�wB���
�����P�z Ñn�rN6�������i�<�X�jI��r���r[����O��Z�*1Kj	iq�Dv��.&�cb��j}�8�%K�=��3�t�߿�聑�i�hO��.ڗ:�R�U�3�o�^
�e�L�`C���(������� �:N�=c�����k�T4��7��&�����#�i]n'[���d�&߀u5��W��=5����?i�J0yӤ��5���{��M�G�]�����|�wf�P~���l�H^mt�"��l��x��f�d�i����Q��w�����6�� Im�m%�|u�r;9����j�{K�=[r� *�������6ǩ�s�A���dހ�;{�̈b����~�3���e���Y&�c�H8��`��S�G��T�.�C6{�;�j� c����*��Pi����]7�
YKM��
,�~�~�
�?��&Ջh����s6�Rhq��S��a� �!�ap���>�r�����
�[��������vX�>ͮ�����Zo�%3De�7�hs;/��&Q5�v�z�y܆�l��ڬ�Op��?�gE�6a��K�j,P�
4�����q4.����ɲ�s����O�y�_��oW��yG�iM��^���>g��P\�>G+��;?+m��M��nb�K�������j�ć-YE<���_�ob����~P�}n��������-���Sq��H9�����L���F	�:��Y8O_�v��Z�'-�3�$CA�>��-��C�C&�Mޝ-�4ܣ�8N҃�0��
n�ZIqx�ۣ����t�@�����zў�!f7r����ǰ�5<rF�Z�ά��b�=xG- �؛���G�*J-��֍�l���91�j-oВ��>������7j*��&M|�����?c�j�:�`�bb��qx�{��mS
Ź���+I*�_�τl��T�����D�3�^��i}��_�lۻ��Lb�lh��s<��((�d+�b�"Ҝ�\��M�;A/��ƄH���ޥ������=�;�������<xZA�Sޫ��� �� ��J����fi�>�2�b~����-��R���D.xQdU}�[��g��گ��^^b��`w--Oˮt3df%����s=�Ζ���G���!�#�mUR(��O}��u%zJ��p�!��5h�4?��)A8T���K���/Ӊc����(��w�n����������ͼ�m�o��-jY��7�I�ʹ	��u��:'mߞzyY?o��q���Q�*��"w��:���-���6��
+��4�$�\vM��:_�8z��߶��g��uK7/�Y1Yp���\F���j��k�����ƕ��*ce:��h&�b(F��#4f�VW�i=���nw�G��O$�C�W�9]��5������j����po���߁�ù��c@���J�&�峢�WY�B�ҫ�Bj��wN'Ն�����r{Zz  1pHˠ��@��Օ�\j`�h(餂�K�:V�'�������^J��j�� 4v���m��s��[���� q�7�:?�	/Cڲ".����0��>R[O{k����Wn�sE�(!����D��I[�&�l^#�(��`��_��¶���~Oy���Ǧy����-<��Әډ2c:ɤg"��h�'��}Թ�A�UZ5]�T1�~^!�6�GG8}|`��
���w�LQ�4����@�gϟ�r��z�����M����h��wnky񈓪:EE�z�[���t��)�a��^��9r+P�g�jS);��O��Ye��e�c��$�u]	���2m�;0��!,��Ն����b��U|��XI!.	 �g��x��Ӿ�L��ι＼�]C���TW�y��?�ܞ�e
��bG�M�BwMM��HË\� �Q{��K���0 z0-�|w����v0������{�I� $>��?Ф�<6�;�ϬF!=`�	�Ao)��ǌ�C3&���C��?|/�:}*�x���?�+	^S&�k�\Ŏ{ٴ�3�'��&>�����
��Ŝ[,g���&J��cY�\�ཎ�l�]�y���M_$����U�?�[����^�����XL��)\3^$�,�𪗭��4ER��tҐ����3�>�R͛И)��5,:ۅ���:z�ܹ�?��Y�{ns�F��siV�^��;}>���?	��>��0ZhM"W�^e��(��`B��{�
��D�p/�Qw���@aĚ`<���s0�\[_u��T�K�&�W��'��m��4�`�v;IHW��n
�
�q�<x����>��ƍ����FW�g����V�0�{{3�� �8�@��$5��Ŕ�i�&m�v��$Â��X^M��M\,DUd�OX�&	�l���y<����-u��>���re�D�߽pvků���|,>���K�-v�-
�@����:�ݿF	��v��Zhn�7�m����s��������%�bcTF 4qTO�ˌ'P�y֫�4R`,y�|;	_E��jЧ�Q`�0���a������77��l�:�~�߰ ͖��DV�c��?i�#\�~�\m�W�Q��B��d�i�T>/�,?ܸ�R"����]��5e3m���m)��!��޽KWe���M�=y��&\dM���x`G��O�1oVW��~�?��I�w��pg;?Xһ4��0:�Y{t��E����Olb��~�gg?	�H���\'�f��U�r��I����,_S�f�����]�Vu!�F
'K���?��ɿ�:Wѽ��7'���3�dY
Į�rx�F}��(��C	�b�$�����i��\ԞS�Jz�SC����&�"�,�]��3Z��5@�A$�tF8���Z8����ǩ�p�8~{�esq����BpG����J��� Cp�!��å5�[]�g�g�PWagE$X_�����F��"�FK�J}�$Se҈�p.�-�B@�������akUK
b�8�=�n�\ ��bV[&��u�$F�� .o<�u����߷�"��lt�]#{�
4�����z<�)O#�Q���V�]3N��NJK�f�_�9Cn�m�7�"��	��K��آͻ��,��_�i_�/
<�RН�B��W0����eF}磤����@Vɛ`�W�}����FĢ�S(�=Ƴ�?��p�Fb��\7���Lrk�Crrk�����ǀqS��Ù�bH������-���t�N�?�S�N��lrD���`�F4��a�yS�̢PE�^�h��7��QHL�����u�X��.D�`��X@��TAG�G}��ĸZ0����a��i�R㍔i��`udm�3cj���Xo,��a���g�Q)�Z�I�Qm�!�f_($E��le"���o��%F
c��6�B�iB�=NH�����#M�8Z�pR����]�ɟ}�������g�O��^����}���W���[O�g�Kh@-��Y�[#�oN�܍�,u��\��֝&)�q���k[a~��1��֢Ё�k������4�'z���~\1(�G� ��ܴ��=UЀZ�̈��hpD�s:)⿑�^G��wK�f`����<:��f�Y^�JT���`1�����̙��ĝ��ҽ0�V�[ڨJC��ER F��%X|���ӟ>��f�a�~ִ���&��Cɤ���+��j�Gmd�ʎ�
r'<c���M��.�ra�����ޅБ��l��D���By�o@�OߕK��]���u���HI8X�c��uN���y�~�K��r]�[����}�K���]�"�Hq���+��|���R�R�)�ك�0%��.fV���˝�$e?�9z��}�U���G�`<����b��o+Z�I�t����-���aA���7���F�HJ&Ű�0`q��� ����Z���dz��kCC{%Ki/_��p�r	�1�ZO \*����]�	p���0lk��Ot5�z�ѯ.X���ǘ����G��~�$�$���>��m��7_3�A֙1J��a3�`�D����Ȭ��p��7�©ե������3�u(��S��z]:n��Ht7o�`���l�;e�9o���J�l���Yr�k/̌gkU����������q��J�̺��&%Onz/ �:��
xWx��me�ye��Ղ�~�@�a�g�:��q���}��	��L�������9��g��˭�h	-��&�밳{����6(�J��L�L��y���#�����!�v�Mz��P<��F�Fl�(�@��|�t|Lk�s`oӠ�+��L��������
��z) F��Ytc��"���~s�'��i}�a�z>|̦6Y%�w!�u��!��.�$��В6�p������K�ہ�tG�ވ�
&[��E�s��x��d��6��ǌ/T�h3��O� �Z֯-�s�ҔK��j���{	C�e�Կe�{K�#z��0�f��!Fk��Rr�3��ԟ��:7N��(��?L��1�tиY\�hq��sJ��g�����K.uW}��;��D����]{�"=Q�n�Ġ�gxZ ;P�i�E�B��(�<�Wq?����2��0FYX�B6
;����j��c0�5���P"������_���pX�ՙsg���_�;M@�I�y��9�PFIi���w|6kk�I���#��s-)Y7Muv�5�k(��%��)���a�Ӥ@ĳ#f�`�^���ASp�80z���Ht�������dE���]��p�g�8Z�1;d�P���G�F�
,uU���z/�=���Fs�}RO�=�OJ��y�/,mv�����3���mj�h����M�MG� ���� 2��6�ֻ^g{�W�@5s�/!���c��=eY% &$�"����I��uO
����ӭ!w���H�)��[�8~�AY:Y���;�vںځ�(z=!}N�E0�`�1��(�l�D�zm9��֛�+���i/{�G�ѣ��x�,�C�VG%\�A0g�phxw�x���0�n����j#�E>I��*!�f��q��R���D�Ek<aoĔ�` '�G�>�L�U��D/�ʱGڹ��E )Ԙ����x��ǰ@��U���<�6���+W�PC]�t)��G�?��4�'� ���������f�h������G�(�?���X��/GY�}�7��<�z����0�W�~n�yn�2���~͵hK[��+�)��&�ٸ��Wf��?B��~�s#�����l����B9�ηd�[�����عK��^�a����ܢdd7n_����@
Ij'LpS��5<�H��$�^_�J������� ������%]V��J�l�%�h������1��=�߳z;�� ž���/�`5?�����{�w��_��B����e�I<}$��phN��������"9}�}b&!J� ���^��3B�
0K�P��c�͋E�	_ll��I����$pU���XEh
�< p"w h0�J[�VL��"4֩�%ֈy�E��5�a�-��BRae�r�y���4n#ܱ�qOĽNdI,{��	0mbxо��f��l�My(�+���7p�J�&=��%����$�D�f��%^e��Z��e������/LVG5
�9�
Fj/�Ժh��0C/�~k=}�Z��#�C�|����)�i�*^�x4�\���MT���(��n<��y� ����s�Ǵv~2��4�4H./����ш��p%<�v�I׻��LE���3r{c�5�*?��@�����Ꮯ}J��n�w�}��.͒3��2�0 +
�8� ��M��bĈfd'c#1�'y[xE��UU$7�6�q�&��M5=��[/wɀ��.�����gvA���d�֓{������15���VW2�R�b(�o7��f������X�ᷮ_�6z�l'���0���,��yh�T��{L�$�י��/����$�P�D�g�I��%f�.�V�煇@�q����In��ۻ/�K[ˢ˂���e'����^a,�ַkۢ����1�rxϨ�ĔB����D����󄓳��:��g�` �'��Z-,�2�mI5|a ʴ�+(����B�v�jt�G�Xm�3q����b��̱�I�ΣD��	�#������ƞ�����V�YI֮14�nm�L����p��'���N�`�Xm$�C����g�n�� �`򐛰Ow���y�ˤI9v�(����
�6������p�H����k�$���������{���|�/��[��)|w�+j�_���!O]����r����p�L7��2�g9pf� 6٢&���6�Sic"�L�Q�"y�XB�)9�4m�XB�kC���4sI,%��Ms�?��غ�E�Xl�d� ��x�F��8��p���o/(�LO��]��ޗ%�f��RnmΦ�Қ̣q�D���Bmc�z	~iBcǀ����mFk�l���{xcB}���p����5�'�*>!��uI+�D�ŋ��Vd�?�Eˏ�$�^RJ�C(yn�
�������2c{q��D)��:(�P���/]��r(����S�)���f�Ad�5�|J��Ǔv�/G�$��Åct�}^;˽�v�+�Fd���zL7��z
�1�b�^9���E��υ">\f�k��rӻ��y�U��f��c5���}SL��_�/�[��_�nk��Цa&7�
U����h���@�-��� P�z�72y�B�R�Fm�	5>�M�s����#�a�� �jV�c�dhA���a�~���L�x<'����B��"1���{6��F+Q�s�z�$�x�N!�8��K(������d�,��v.h��}�$�]��
R�$ΌǷ)��<f�j��|��x=�mB������w�ag���F�aR^��3�5�����N E�~j-|����Ѯ�u6T\���RDF�DX�����lF|Mp�!����z���W��ش/�dǦ�q�[;��8��~�����8��&��VN�l	Z�����fe "�P�l~h��D|��J�(�qq�߸�!�,i�fc�s�M�<cF�4�	-\f@=�c�N����6�\�	yM��O�x�d%A9Cޫ$�p���,�3�K�Ħű`S�H�$i�<�	%�i�߳ѫv-�oŽ��J!�!!	B�I�T�Vu<���$p����7J%�v��XMuQ=_.���r��ӳJ)"�����k�з�Օg3M��>Qh�XE����`nF^���"Y+�mă�y5�a(^�	6nԖY�������� a/A'�%��[o���^l�`�,�i��˄4[*����ZGR�����؛p��=�I�S�d�����IXʘZ�l�(��gl��{�/b���(��Ԥ�)�m��������u�;nYv����s�]�B�����=����w�����j��J�/��ɥ����+����:e��q�������7닥�2��7���c�\�	 �n.Y�$��pjJ� ɅWiC.-�k3�� ��ULmF��Ҏ���>��~��Q��3��a�p.	�P�Ycd��T�� #Y��L�7x:5�,\?)�X���|/�Ġ�L�ن�yբ���ܫ��jTv�τ��u��N�<3��G�Q؏�j^T}�>yʼ��eCN��������);̹F��yf��`#5T���r,���������A�ga�F�KY���*�Z4'�R5��oc�,�C&�JlF�ckj'LŌ�s|���ضf���¹�i� ^���,]��!,6K�8E�),>F��D�� jK�m>��9�U�p�|���0��x��&�7@1L%(*=�DS!' <��a����:�֛}p�g$�a�Ym�~�/!4I��\h��4���D̏8�w��G&��w0b�����A�K�bR���mml�+Q�ڪ}�3��&��x!���!i��C%I$1���뉫��@�~ss#��3*�����MNF��b:���x��8i��n6
g@�ރ���n%�O��跑LOP)�bf������UK��$��][[�h5���+��ϞG7{��<�{G���[���Y�����0���ý�t巶7����zj�
�q����&��`�_�kL����)p�2�f������vM�h8�Yi��*"�Y��1)�V��җ��
���!� 1�db`4o�26e��+����Eh�5��FaT��a���?��,,�e��ߌ���t�X�`�8<y��Q�gK����\��ڗ`��l���˚k�����(%��VG�*U��[F))*A�Q%�3�;������V2�g��m �QN��IB��O�)J�� ��QY�<(����$����]@CP��6mx��F�V�*ytc�_Α�lB�C�� ��l�N�8�����&���g̦l�o���R߸Ƙ�J�����hF�
�**�)�"�&�h������Ћ
iF�`Jw|L& �@�����/�屃(�4^FL`��V�0(2��	�	*k�a���V�DjHȠ
N!��y0�B��b�����	��,n��1?��q��e��o��������U��ӳYj�>HBo��ݼy�����@3�֯�k�ãG��e���`yt8�����4q�u'tTP�n�����7-�Pw��#�_��
��1�wF׉J�iG+�&�9K<T��+�ЅD�]<m���'�|�Ii	9�`�d�?����ӑ�r7�]q��g{v�Y�,9s�2Ո�ד��5�߅b�˒ne~�V�/����6��&���g�<Xv)#���U�N���m{���@���ʏ��7�Z<������ڐl(]�pŸx'&ZXH0�ʢJ��`�auQU���5�GG�QS��`Ƴ]3tR�P(T)��J�H�sR0̗o���q
�˲��!�4�^c
e=Ӏ�y2 3�`#�Z�<�-�m}`�jȌ�D�~�@�YW�����?�o��6���>�b@�$j�It<���ktx���9]dbh1�M�hӢ���!��q\�$���0'������a�Jly 6��������� g�!$�F�Ú͹�:��=N��h��j�gCANת������K�	�JM��<���fM�������B_�j�т\���Č�&�/���}��ݻ'RY�=S��|S(�S�2C���S|�A��a������C�/l�r�mn��謚�}J�t�gă�qZw#^�B�ߍ*(O�>�^ߪ	�j4�^���M�8&�L��1�ʿ�"󊽕�ư�>	a5d�Z���\={(��l�v��{��w�O~��_OM��q������}����;9��r�s[�kyTP�Ϟ�>�୰�Wh��j�}�A�����)������W�,�JH�N�҉���`0捣c��B�<:ZW���Fš�R��!LH@�JJx�bK �����i��k�(-�"S�Iצ��5����^Y�^��|r�+}�[���u^e�sݙ���-�j��0�3��4 �����6��2���Y�Fe/�o��zn�69K�]T�#M]�|� PB[Dw|+�#�%��%����w�����NFG��F޳|�֋d���WJK
�^- <���f���	{�����\��,��^�
�����aś�=���S�obp7�qa��z����������ll�c6����ecH���X��ؔ17�-��˗.�+�.�I�uv��������g���X'uQ�ɭZh/ŰM:Q]�x6��e���KQ�%��T��7[2q���8���bP�%�|_�GRy���Ծ)�?l�[.%����#��?㕡`����4�Vպ��wz "�������y6Vـ��RJJ6���%��	<Z���
�4]��<3�X�R	�ׯ_'�	fA�=w!\��Vx��Yx���V�,$�M�8��Q�8�N��؂0;�p�K}!d�ˣ�ྗ�Z���\S7�B�J���Ŀל���{����fi���˛����9-�n�"���Fr.1ˊY���'$��I�4�r}�$2B����`=;�}�T���
w��ٸ˰�j�E�t�sW�����f�gYSO��}$\���F�Ĳ@��r�ap���M���B�x�u��|RJ� K.\��e�r�"/�Z�nX���u���ۋ�abxbW��݀�Em��ٜ0�:����uH��^׬.�U�%��k?��3ODS�(b��K4B.\���,��J_��������,�t`��=�Ś�� Z�	$E ���J�K#f���C�C�y�}pB��̖�M�rਫ&�܍���Յ�V����[�v�E4�,�>7R��-�x���P ���N��������fe�Џ>�0�=s6~o�xh�tD'Q�/^\;��Ijeu%<|�o�64���>#��on-�6�b�I��*᧍2��qn�/0��a��F��ڤ:o71�C]���{���zyk��%��r���m���z�
�[�"���w��:� �+���EHǎe��Z.��`�v�_[�ד�e�ji=*PF�)T��P�
h`�;�x��_�o}��@b������&����}���h��=F����;I�l	E\�˟�U���GCt���y�����|�5�8`2��2���<�]�m�z*&�PI@趿of���
�b�ī��%-��X`��A�9b3
AoF�M�DPd�����_P�A��������
����XЋ/�Ł����V��q����������SK�-m&W=����9��*ڴD�%k�ؐ诲�;Ϋ�� X�K�(}~�)�u�"O�_���м��w�K�n+gP8���&Rl,	�Oh��*C�㶪�[���Ճ�!�X����E�C�f��H|y%hJ�}6�Y(�^��L1|!���yZϛ��ؔ=&au��� (�D ����8���� 
���g?cu p��� ��νn߾Ů.t#��X���� A�M�����I�^
?�����Ĺ�fvb/ț�24����^r��o�a��b1�Ct$���D؆�Ė͸	�r	>�7n$~3^��"Y��7����ޱ9A���� �07�j�Tv�v%c��}��<7���r�$̻m��ȼ��Ɣ0*&֏,�߼��*5�9+=g}�yf�V�ZO»U^p�E�z:���e5%�^Q�
ˣ��uW��(�6��}�SKB,�'�*6?j� �����),R��4��h�I�m�) ��z�"�^��랤��(����H��
D~O�iIQ�YY;Ø}{g�T٠2By	���R��*\?�kt�������D�.]����)�T2���ө�V� ̮�؋P��p	J�e9���$�C*F�>����FC�e�AR�J��Q�M�p9M��
R��p�� ��_�5�3�N��T`��ؒG=��o�;�K���c�M����"��qt�'�W؆�s���.hƬd�F�P�G1�[X�6�b���t����)w�9ə䦭�ze�7�ײ>��q��-{�Zs1�{\��OtyE��`t<�$�	�߻ƪ#㿡ād�צ2-z��k��Y���A��r���LѮ����1e6�j�j�"d��b�Dx4�H/���upz��P����:�;Q~O-�I1>0����\�^���0 �4�8�ѯ��Ѫ���h$�����#`�~�y�$�Z	�v/Y΢��-j�3�O��ˁ�,�U@�@N�27���㻀$�&��g�����6�ۿ�[s00�t��E��:��2��=jHty�V=�~���H &!�0��q�M^$<��]-+.��N��7t�px���ןb�R4H���n_�k��=7�G�����}Fu�����fLda��TO���哄��7l8�T<�����dF:���,9e����&RF�u�M'-�g.��m�م�^_CA�D�\���ߠ���ג����hC�����0��O�>%�t0Z";	�Y���
w��vv'���N�ri�y����;�򹝦0����V�[�-����9/�%���?K�J:x����*�ڤ�Gq�8��ƫ��:��N�`4O�DK4�W����IBV
B��G�Y_t<���o���10�P+��Ƭ���
�	h��������������E��{1ٌ{P��ѿ,,ݍ��\V��I����Y�e%��8�:���νy��<��+ ��-׃���ˣGUp�ڗ��ߪ�{r�a��b�Wyzѥ�p!*�����|=�o�ЂE���i�Hz����*�X�y���Y�E�i� D#���׆S�d-;Zy��c6�h���S�{��w0/�9D�*xaW߸��~���Uͬ�C)0wei%�~���c��O?��PT(��b�̝Z��VL�����B#�{�o��PS�g�Ss��Jʕ�W�
�ɍ2��~L��^�r-j��x��2�� 82�w�~��Y����W��������(��¨��::[6^l��I�����񿁐z��1[1���۠	�E�Z�#�[箋�M�-z�}��i�t>/�Y�s%�������5���VI'$_D���ǜ2�$�:�w�%�x.�@�gyxt8�������� �J$=��[����>:ō�lQ|�oS`�I�L��\�p��ˊ0��i(*{5�e"�;�Z��Ь_��i�D��\L��O������pd����QVK�"3�6�Qt�G/V�޽�����9��<w����ٛ�o�a�y���F���&�
�b�z9XsSI/��q2���Y'AY���,U���ʢm�!x��jcx,9�X�܍�t��9Z"��Dv�O�{K3�׷�~�����_�"�'�/>�$c���q��������)H����ɹ��,T�=v�Lه]�37F+�/ԋ��EB�x�>��Ǟ;�ctc��߻ǔe�{��$�S�?�ᖠC��n�C͊b��y�?H�
'���Ed�k�b0��e�(mSM��)C�A�~�Z�Ul3Ͻ�����P�B(��3c�I'��u'^�	4��J�Sp�g(������MZ&�ӧף���niy�����V���M��Q��1��x�D��u���������Q߈.�w��#��;�ñS`�a�u��T܏͡v���\��`��>���̙K����bU��F�����+�����$�cͬJǂo4`������.�hr��q0����ޣFG�_��/^l�Ͷ�gT}�WQ��3�G�H��*� ���[o��|�n�t����������o�
�e�O�O/����"�0�v����%�~U��M&F�#7U�S$u�K�-���j	��~JX�r׫�QV�'�7��ؼ�%^�^;╄0�2��1zTD�ֹU^p}���2��M�����	�`��o�X�$��ea�!��!�/_���ƿH����|*��N�*� X3�u�MG�cJ���?	g�����������0�k/T���3��v��j���`����ǽ�G�jH�����;���OvLe��G�@(Q��w6_�F��B��|p|�ƍ��/���G)�@V?ׯ_���#��� P|H��� �������e������B����A�M�ma�+=r��rB�HY�ԪR�8��U���ɍl(}�#��;)��^s1bJ�Q�vbj���D�����F�n���G�J
��w�I�o�l�^'^����p~1���WO��:����jN�b���<s��*�W% �M��kR�JW�ڸ9e��4���f�U���~6e�	����F.��uo��6�'@�]�|-|��_�x����E|���sa��Z�w��ܙg�n8����t�OcD��h_�pu�TL�0b����U�q)cV
<���fIţ9��ϻ���!\&S�enh֤:�u�l�`���=�8������ �6��z�|�I���/�����s�,;�L�nHL�%*@��x��`lD�Q�����Ϯ^~-�Ǡ���b϶VI�Y$K�nZ!/Zaς����w��WJh� �����H�q�ڝC�S��e�`u�Ld��7N�bf�zA�1�"��sǐ@bS"bl���-h���M<��s��Zs�LY���XT�S�Q�E�� )�lH��F�[�ى�Tu"[�T���u��9D�Q�^�Z���m�bV��<3*XU��^�Q/�>���~=��/���N���>�R�k<İuJ?!���;4B�aϾq��s�}�G��r��2����BE{F��R�� ��N�������*^�@����| �wp�����$��l(Sv�(	S3.���%�z==c����s��lNP(�������p|�gϭ�����\�~[V0>��`���?b��\to8���"oVAY{)���8��o����W�ָY`�����ޚ�{��|Ͽ^���K0U�?*�a����b�7(�R�7���=���Y{_��$`^�G#{ƭb�������B?	I(���6�xd�a<ΰ
q�����'c9�u���ɍ�'G��0�����i�kR�y�	��V���kXЗ��C ��1g4T��F�j7��EqĽ�2D��(���vDB#:PQ1��S][e����{�h�᭾��۩y-%��zȹ޳j�xbyR`n�s�#�?�[�&���UBg58��U*Y@��n�&pћQp����[@kqt�������p�q�BC����l����Ov�X�n&���{�-�0n�k�_���*��϶��q[]��*j�~�y���;��@x��uJ(m(�',����NYA���Q��v��yT�����s��qQCh����d\x�h�/-�}� %h�cj�u�\*�e��gR}t�<(��c�y�>=V޻���j>ie1�p�J�GE��9 f(M���0�>j����E]P�@U�C/�̄��2j�*X�g�������z�>�iװ�YY�4��z�I*`@=d\oz��o�Vհǒՙ�����g1��e~ J��0ii�,��e�����O�F�~��	�߽C�(\fo�d�ԘK�ԭv<3ʧ����\��$������l�@C�vW0�2��C��Rk�:!���mLF2@3۰�Gc�0���$�}���������s��Y~Ɋ���p�/��O�)��J�u�)0�I�r�"��
���մy1S���;�Bv�ߜ�V�����ݭ�.*�-*��n��N�<7+�iܪK��:��C{)nV�-�P�/k�(���C�Ye:LY���
�6-No��<������}��˽DmaF�L�HQ^YrhC�5QȢ���
ĩ)YZֈL5a�$ĘqV�U9oC��L93��a�i�'�[Q�O��s�����q��3oDkߧk<L���q��^?���W8�<,��0+�����(��gh����p�D��$�D��!,�P��A�1�f8�*s�̍�ۂ���|I���FL<N�cJp!>�$�M�߇���_��w�)vp�����X��E/���UG[&��7���{��Kr%\+o`ee��9:��S�&�Q�x>��
�	�M1��n��Ⱥ�ͥF	/��wݎ�=qj��j���j���	��+��V�JB�k�*q`��US9�{.�,8�m��%./\��k�؛^�����5X�A�>�\��T��K�����+����{�k:�j�g_%X�(��YqA(��FuHC6�f�L\��
�VV����8��w�<������DD��?p@$^�������=�f�z�y�9$�6��G��[eu��6YRZ�/�������i���dƅ1��<�,\r"���Ҕ>s��E,��1p|�"~�v\Y!aYq�G��U��^��e/��Ǣ#y0���`�[,!K����F�F[ ��M�(�89f�P���Zk�Ip����=�_lݯ��U��P�4�©M�P�C�Qf\�>��@1��TSH[��"�`����c/�~����̼��ҵ���+�iK^a[��<���������6��:��;���_}��x��yt}�Ù��W���L�A�mĉ���w�i�~��_��?x?Z���a�oTt��Ea��ۂ��~�Z"Xh��!7-uU;J��{��D�k�z�����%���o�l)�/ʨjj��ch�`��%�[��93qq��p�0���ک*��j���v�y�7��Ԛ�"A�p����YƒgW�	�\6	�"���͉��E�u�k�u�m�,<OGx}��l�(���ԏ�R���mD��*�w�};��A����r��gh���\��u����w�P�0�>���J������v�b�m;�Efl^Z閼�;ۤF��H@�d�W���=e��X$�4hi͐C@G���o�=�<{���.e��b�$�1����_�T�M�ra�f�Yv=��l�{L�h:EJ�&ӟ�pi]''�!��,y2J�g�	=x i�-���P����}~��^�,�V��1���[q����gFQ�����1V�`Hh������(lv��vw��*ƞ{��'�{�^�� nFw��$�sV�)/���ZZv��k0����5t��:�¼U���8���KJ�T����N�H��� �TJ�x��l�<BR�<=�n���ܹ=��1K��fL@!AU��j�
`Z�F����r�-���,�4��XC��\�f�zm�����u�?~��.^����-{�:s4���2�0"t6x������O�U咐F���M�&��R������@���l�~����y676��� ��Jc�e�O>�=��L�r6���Z���b��i� T���
M��yB�-����o���T�c��%���z�xD�i�y���}��Y��.�h�m�,+&�L�Ka������/��;����-)��:�t<'Yk1�����k�����Z�EJ6�chÎ���V�	F���Q�X�F#F,�
W|+�U�X���Y���É�f�@�h]hu�w�>-�:)�&N��x��Y�ۈ����+�H�k��q����1�ǐ��5�`�T���$�E1of*[Pc�hR-�K}�4mlU��&�V�u���mdm}�Qƹ޺u+������1�!����,ndb���k��5
���o]��Mn��=}��7sGNb�����5i�;��L���+��;|����g�����"��O�OXn����=�����f-�|l�bM&��^�qJ��!m��k��V����N�#�F6��:�;^������]�1�7������KΘj��]��Ȝ�jE�L���s�c��a��'� �y���am}��.Ti�Vv��>�����1���H�Y�π�*���;w��9W_{��V�l:H���ׯ���ݻ�'�i/��f�;iy���f�D��`l�D��x<�����b`�`i�(| !1R`�3�Fh�"!�F�����2
-�@���￿=|b�E|.{�{)�UK�+�6�� ,��x�>���n޾�@�-����U^F떷��<��w����c��w!x��W)/H2u�)��VRE�V��f;^�Ǿ�(|M�P��(2 �-��Z����9x��iB#ʳ����vs�5Ţ�:u���]��:�|� �U�|U��~�<���Y�`��jmu�F���� ���������f�@����G�Rz H�"��?�CܯDW��S?$�x��g�Sz��H��},c��V�`�
�a]8�H���T�y�3�f��e���f<c�д���>e�_d�x!� ��), x�>����ݴ��Cm�+0�U�t��ae+4��-�/xee�"_�U8�=����L�0�:5:]���$�VR�:�zU��@��&��A+���e�!ڨ���Z}^YR�w�B�*�*Q�,0�h��M�1=��ԉsq����uEA�2O�/�]�[צs�W{F�s�#�~)%ɺ��J]gzN4P,�dN��r��k��"��ʹ�8f'|�f*}����R�����i���簂�4:����1F^�>=���1�^ا��U�ձ_<� "���O����)*׳������Y�ʊ-��D�D$)��P�)��~��G\7$��ʒ�����J/5Ǯ����,��S[7.�#R��[�"c���*:mB�J���ΧO�ↁ����&!2��X���W����}x��wO���pat�P��O}��K<-{�ϡ~�*M?hK1^�w�/Y��g��}�&L5K��>�+%!�%5K�fWTᑫ*2GO`X7a�5 4-m,�:Eh��P8�[�q� !��W�S�Xq)#����M�Pݳv�1�Eȸ�J�Rv*�hHAf-	��K7�J�� >�d-q�O�&��{������ +��_#�������Q�G5�Zm��7갹�E��w�k �xO�>!(/�yQ3�gϑ��H�$޲�FkɎ��j��Fc�Fd���* �FEKm5;c��W�aHê�.m��d���� 9�����'"bunX�d�2x]MX��+��^C�\L@�!��+���h�F!1�dA�̦s9�E�]�>7z'NZi)�n\�U��˓ j��PA���_���A��hδ�	��������|�p�UM��<#��m��鮣"�l���P�����WC�c��l)m`������]���������;�Tf��D�T�s�k������ڤ�~��;-π9�O�<��.���N�y"�U9@�x��5�p���c�}�;���<H6��*���ʅv����iy�ejD��%M�0�ą�5�8:��YA𥱖�^%&�ބp&����]h�0g�4u�ŋg�޽xS�~x��r��mXP�ro=˫K���&,9��2��A�b�6�!�3�&��̦'b������z�Z��E�3) �0$$~�����GRl>.��-e���VrL��|�^�5֒�z�:�k��i��"�I7�����Jl�vM�F]���"i}�a���Y��׃&?(�+a)��/zϔH;-Į�������6Rl(	���S+���]�{�����e��?�^�=�:���C�4��N$�`�Q�����Ux���<�~4ڀ�p@Dل^�`C�4�`�lB�{��H*L�C�n�֤��v�8^I�ŀ�a04��fm�b�m�i�������4��K,kg)�p����_��r����=A|c�����$�2g-��OZ�n>c���kMݬ;I��!��WWp}����ݞs �؂�g�%�xiJ�:�<�V�n9?��-�zͬ����/Yn��\۶٦�_j������y�'u�q��+v��޳�H1�B$�����zz�J׭��s��w�G�u�̒附��5$�rJn�P[��h�8�0�c�DWȆ������~���aѦC�oQ�����ýp�[d�y��h�	�m�H�	���	�Y�����Wז)CȀW)�R�Bޟ���GTH(���Hc9Ax�)�i2�F94��YT�ey�������/^�]�����ko�A����#
|��:2|;,u��_�"�gD���K�/����mٲ���)AL.0�Ӵ�x_C���m�*����[5S�Bsނw%��,�56��(�CI��e���œ�Ɋ�n�`�JH%/�/��pi�cJ���յ�����>���7�#�+�y�䭈���,Z)��[J)��9~��A4Y6{�-�6� Ox�1+�kfKH��4L<�n?}�"܊�3Z2��UZ������E;Ί������QXx(�?����3V��?��d�]����ʄr���Z��sg��g�� d����A�g>� �Q��P%�kI�S��SF�ʮ��6�*��-�0|75\�z����_~A8�$nݼMM�� �`]:V����!�P�p?}�������	�F{{?���A��2����IW��C�u�j��Z�������P��F�$\]k��A�i�*k��/�gŝ��RB��H�^�N��xj��wC]�ǌ��^,Щ��9+�'^@N���Fn�nY�$��kM����(7]Ӣ�������M���+��2m��df�<"�5�l�fk��.�����~�����/v؊���F�P����[cӱA���CY�5�2$�a��K���ƨ�*V|�[�S�Ie�n�)�f�ϬGy.)�>k��m���A����9@UZo�2�U@��v������0C�1��^ΒC�a��Ç�yS���/~�(
^̴��	����6��ut��/��܌^�A��W�`/����ˍ����V�z3f�K��%�z�u��E��"�.TB�X	�z2	�bK?�C�E��$�"lD(I$P������y��{�G���!��z
%�:O5�V
��,z厥�֦��#c��2Kx���ΈG�uH/J�us�� �i�N�������t��V�����D��~�)5�[�\jӂ�8C�	�t�F	��e,'�R���GB��{d��l���Oe� e�K����Յ�5����sK`m��܇!�+��2$ט�Wj�~/eݪW[#8,2b�0aa?6RwlLs��53�Ξ9��ãGO� C��m,4gi��@�8�J���VԢ��O�A� ���;�	�P�>؟do��ڊBBv+�Y��dD����EG0�vCe���%>٥c˃�Ɨ����T^��%��u��u��m�d�3-�=�R��yhe�����ȟG��B����,$�-,sڦ�d�j���#*3bl�{�1B
��1J��XѨ)�0��*��H�ژ����P�c��ٳWht D0RO�>��E�L26<���g�8���g����o�-ܸq=���P�766��E��?������K���Y�V��0o 7���V��!�4��A����Y6Vo)��`u�@b1�8Nh�~ξ����=�>O���c�_�|5n�	���q!���i>�Y��A`�0&�;,���&^W��_MX_=�5R���<>�����_|yǨp�`rùXZ���Q�ż0{�筠���l�VU`_?��b���&��o�0�G�i]ІJYd!�t]�<^��2�f���6����E�yw�+�q�X.��##�bOaQ��$�^��L��8JH)�:6<��Ӭ��0�&V�^��B�4�M�	
~a�7�^�|��&e��gԋ�+�d�X;�������{�������M[M��>�q��%��p�w�|<�Oe���{?�Qx�"\}��ph1�M�i�*�rV�q���=v�R
Һ'�>u�C��=�/YS~��R�'F,�T(Ѓ�aR�
��r���T)������3���4?z����[�ƛ|�����;��I��u�(hh��c��^fI-D�^7޼�����[/���l��L����]��6���v]���>i�Dc�9ٶ��rWnf[�/sm
`���״w*�����GJ�ywW�V��kR�^_�\��z�̺JIߓ�������K��"�(� �in�5E��eOBn�x�K��R�.�n����y4�ʠǔ�Deȫ�"ε�
���p��j�=̳g����t���A���{��^3��D��e�&hh���	Z��H�գG�@�	����\� <	 [��D��qj�Ư�2{˞i���F�T���$f�	k],y�A��ϟŃ��!��U��N�A�������$���v�<p5�7������^����G��|�B��A��ъ�k(IuT�+��S�PY�LeB�uݶ�q� ��ػ�&�<m<(n%��H����|	��P�'�� �ʠ��+,�B�4��r�=����\�&���}�W��-w���=�^!�����np�����ږ�w��GW�dA.�G��xF"�����kO��6��κ�H��'�f܇#p���|���t%�h91��!��%I½����&˱vM-g0���"��~�F��M@f�c
,���x:����l�AM��$�LC�����b$�:PYJ-d�H8���x��jcF"~H�%�G���Z$j�xA�捆��&^���&�p���#������Ex n���u�4�#9�7��Ѫ��㠽�&%��=]���c��=���u&-���_������'l0�ꯂ�x�u.��6�����7��X�Z�v0�ߥ�2LK��U��b#|�Bz�c�UoV;#�0P}ϻŢGRbNB�|������'�Kw>i'����&<�Z��S֞��iR>B���
�L��j��3)B[7�;�x=V~��	הC�p��$�.\���~-ƹq�������E���ђ[K\��^DJ(��"z�����ͺ$͐Z��Kk����T�k�t�`�c�ӳ�y�AI�*g
qӻ��t�#\K q*%F�LP�LfA��r�d��$봪24j�{�{��pC���J�� RAj���mY6�4T5�(��x#U8}j>�vwl�B�uP�������WЍ7'�X��Zn�r������M;�Q9ՂQTMZ�K�N%�+����\%�4GpOa�}"��>G�olOܯ��JC9f2����R*��x�N
E���2��$@�T��MJF�7W$�,�T�����m6�7&�- �(S�mA�o.̪5Q$������Ө?��Cb�9�ug��q6��Ϟ�l�V��GF��p-�����y���MAb�5�zȪ����Q8i/bM��o�����P�,ݩ�G���)*~@�A���AƁq�H�׉��q[x��f٥ �pk�*c�P:��5�`c�ϟ?c�A��M��X�}�6#��/w��͍�a?�!�� Iܠ��jҹ$���n�zQ�l�*��PȜ���C3��񞬖\ZS��5t�eVS�,�� �������b#j���ؘ(%�s����%-��@e� ��=
U���s����� �����#�TY��B��r���mD���to�|��ٻ�Oֽi,����|Z��kl��@T$�2��<�a��=��!�O���q��,�u[�8?#��oߺ�~����uh
�9�y��[�lO�A��x&�I�th1��4/����l�Dx�A8�A	{�ω9"��laIC��Jۘ���~i���ԥyҨ8 ��D�ͷB��i�����_���a�u�G������%��؀֫z#^k/��m7B�}��WJ�(;ӵ�zi�y���z�쒬J�,s<-#+jV��g7ӗ�|��gT�i{	V�d^��I���)��3KN	�!�n��%�|���m� V�k�u`�vS�D׬�>+������B��{�s.�4�Kuޒ� �3*B�l��SH�䖄��L&��k��rm�1|����at���xβ�˗���i��ĳ������sO�9��'�5(O���a4���wӞ�c�Z�Y�e��[�pв�KKu�O�m�A���H���U`�;a��%��?�o����M�gsx��A�%���[���Ms�L! -��B(��s�"�?۲��i@�ux�����%���un�/�x�H���n3��KPdA/z������W�j)�[9%�-e�yM]QJ�!*�9�|���[E�u䏛ҡ�<���Y��6]�6�:ϸA]]ޗ�D�����+���ƨ�a�Z�E�p�;�
G�,s��g�?�Ԇ�A���6e�9=�<Bp<z�,�ϭ����ɕ�{���#Rs�!B��sO �`Q-wd�ֵ\X�hf�BHKVW|2�)����5�d8gY��H�ٯ:n�v��q3^JdL�]�T�hke�n�[nN��9����=�g�!�?�`׵�>\�p:Z����gQ�'ai�c�0����p���-��o`k�i��b�`�<�6���Y�5�ǁ��Oy�\��l��vJ9��P¿?Kf�m4%�D1$���e��Dp<�P�R%`�g���
 �����Pg,�_#%��S�u�e��uL%��z�$�B��O�I9t�%/����"�چ.k��Xy��lTzE��V�P���.��p��N�w֏B�ư��oǜ�Q��	�R�������f�eׄ�'��x��6�=�a夏4(C{Ϊ')q��4��V����JkRM�ʮ%���K���bԬ`�%��^ԓ�Fy�.�&=�m��Th  ?�����>���z�F�Ix��<<}\�8�b�=>�����rk�-i���S�{��������t��)��RJ1G\�]�"�UyK�d�5�-H�ئ�`E�õmRl��X���
+$K�c���%�u��.*"H�h��[1��Q	=�� �(V'���\�/��zF]��W�>�h�}�;�kT���.����Me�mD��އ�lm���	q�E�9��� ��������M9����po�s���4��rh����,���i-��۪Px>��][���S+enL];']�c�M���E��E�%��H��4��"��n�e]ȸ��a�%
���15,5,���Qtߑ}? &|:A���Y�2�Q'�	�[X���"kI <
L�%�hDn���F�
����qf���\�[VX/	�2�v�%>��?�T��|l)��$| 0�mslҔ����w󥸚$<j	��*�=�WMǱ���wu�G��mKyZ7�����_�^0��}�P���(�dE�j���T�8�ޘ��R�:������=����?�4�uk�Dj�7 \��;w��Ql���������_���{�@Ҟ�+o�ˡu�+�Cʸ&�����X���t�����"�䓄��2���5�LmK�֍�PN\$C�?����@�~o����+Q�FU8sz%\�r�D��H�£�����l��U�Nx7텱��զŲz�O
������T�S�&WB-VVe,YbY�:�3Y.I�-�v�ɵU�˃]��=���"�4DvY?��M�h
�t�~�������^U����>X�M��H�R0[
]�g*a�� �Խ�:�j�a��3�t��b(��/���.r�+˷��UX"�Z[�M��1�����o�;；JgH/S�~���,w)!I�C����`��su)�MV�g�l��[��~N�U�)%�a.�Z�X�U��gSd�XdÓ�Hn�B��F7�6�&ۜ���kꃨ'�f)�1>G�f�����{��gOqz��AԞ����/�#��ǳ��rs�x�0ю@/��},�M��B(�*Ԗ�'�3�DnR�\�CKH�4�N-.���.dK+W�'f�����l�l�yr�;����݌�
-�Z���h&��)�� 
m�Bn��2�������<u������[���g�Ke5SX-�bI�h/^�D�)�>]�v��92�w~�67�����(4�����p��������x�QdC���x��x?��G�����}g�?尵4���ݐ���i���jϱ��K���`)z.zޕeE-(�&�p���-b�9������vhC���������B���Gnr�%H�ܼ��y2&$Ԅ5�^Q1ۍ���>��s�Xܵեpz}=�1O���A�cW(�޻7�7�������=/�r�E�8JS�>�)_�ѱ�U������%�t,Q=�喵W+��/�xe���vF�K�4���ޛ���0�`To��6�q�?�]k����/�����'L��/D휵�9Q����2%��!2���V��>c�����{$E�^�h9�c|��5z�h�ϭ�JYh�Sx�-��S� �\�����w�OM���	|�����Uٵ��7��m��#*��+4�xl��I'�(��D��F�Mb���kK�+��mN tk���/~��_�as���[�Z�ﯾ�:ܺ�}�)s������u���֊��A�(�S�O_�x&�=�>��a#j�g��c�r`8gS'��7���{���Av���N��R����6��v5�L�u�D��(���5�o?,γ�t����/Y�Pu�Bק����'���k�Z�ϊP��@����m��UnwW��3��P�zF�24���g�U7��z���D�����p�B��؊Fd'�����k�ⳉSV���Ga�����iv����������.�m�CR���bd������5����P��!!"��y8��'�JyR��M����!%SY�o@�ƒO�����E�Խ&3�w�$}�q��o�{^hv���O���.�Vm����$Z��PŸeun��KP[��eS[3�������ڝ%�WlmXo�˽襄�,�,� ��n�r�Q�*RG���Rh$�&iz�D	�����"��[t��x��t��z��筮����X���<+��k������}wѫ��{�V��¯�UPJ�Uf����?Q#G�q��c��f6��% ��`�!xh)F?��P,�Tr~b�������ԽA"!�%����ᑭU`�Y�6܃��e�`Z�
�k���Yf�g	7�d�a���dU�	w�z�fw�ЁM�����y�@�X���ĵA �Fb�y��j8�i��YbV��f �e�Ⱦ	���,���s a��	N
�/���hr�����꭫�xW-[.>p��'��y���%�B텳K¨cw����^:����pro}������՟��U�{\��{�\�����/$E]8��F�)�@ 	�b`'A"3�C#�?w�b|��	 ^J:��� j�_��_�B��y>����m7�����/�0�R�+˚5Z[���0(�tA�.Ϝb��� a���.���X�.	�B�^>�e��>��'O�2���D��'�|�bB����8�?W_{��� �hqP�@�biyH�
YE��q�q��rb,p=mQ�B�7�6YW�w�-��oe������A	�4��pa�}��g�}}ۻ�:�Od��u�����Z��-��~]A�����w.�5i}k�/�XA��* �kֳ4*-��K�I�k�O�6�����,e?y  �p��2�!����R���F aְ;��oo�{ѕ><z�U���_�)�m�o�A�)_RRYc����O�v��l�q	�o?/���!��i�Q�4-��j60�0��v�Dl%3U>�WC�	�v�pΝ;C`;�{�.��Qj�n7�l�F1l��ћ7o�Ђ���7½���M���^�+
r�6�c ^Q`�P��{�;��f����'���E4
;��<VU��<(;��p��xk�7�~���I8�I#Y4e�5MC&*���췟�%���SI0�w�M�����T�C厮����1���UzA.664�׸��2�Mʱ)/�.�&Y�NV��m�L�'���J���
3l)��u�D��V��{�T��d�KAJ]^�Σ�c�S�bG �����+�Iȏ2W�B���bb]�����/]���5z��AbFy���p*�����o���s�҈�R����a�L��P�W���y=6��-��2b��8���搥>w�lX���ּ�t�6M�q�n�A+��p��PX�\�p)��W�1^�^{�*F�6Ƒ]$+?w���}罰�v&̦��/6���OL'G!�6�s M���c�Z��՞{8�OX\	�e@�]�Eɤ�K�-&�%*"��R�«�A���sH��Kx~XV�2��_��׮���쭼6-�t>#�3�]�-��w[��%��ɻ���V���cb�0O��p�w�FKM�zJ��ؿ���y}���VA���$�D����MJa4:�bL�(<�P֜���0����*�M��^<���H� �6������D��mo�E��2Z��U�������|�#֩!GEt�kD�^�_͵�w�b9�ݫh����s���8�������Q���'��������d�<�
7U�Fe��=Xa�j��8�cî,��d0%y�����o���X��Q#}��O��7o�}�������2:Kl�8/R`�/C���=�L?5<&���M�EK��b#���1V��$R�yҏ���cD�xK.<6�Tn�@ yx�a��b�2�Zn��[-~xOH,��*o�%�������(�\$�������ӽ����.x/�m!�д~x��a��W���tPVÑ��*���"� �~��U�f�Z��:%�l�E���=겪h�A��,�:p�S@���Z�!)��PfU&���Ӵ�٢�($ePs�����$�_q�[ �:5�(��4�FM��,�������}K,&�k��~c&���rX�B<c�0����&�O�Am)���4��H<����}�|>+�`�D��e2�h-�N���Q��|�(jk��mbUen{|�(�ÚB�Q��`�?d0�f�M3��n����j��:F��(M} !���p�)-~/[9o�TJjҍ
��$��n�&�5
x�&�VbD	0	��j�Vn��[�|��C��i�X�ɊW�Y�(����wW0.���2�\,	�6����+�_C�}S�P���vS�HH���W<�Jt�1���z�c��r�9͉��y��D|.{��� >ם)�cn^~�ҋ���CA��2�V��6J�^�0��=k.z��V�{��р�{��KZ����n�Yi:�I���:�g�u<�7�|��\�������^�}s�$	V7yo!�C�L�������G�@fI��d�mI6��4�ñ��52qs��%�q�W�(�ܢ/�����&s�[x��T�	��a}]�$(�l!nC.�T��!��u�Չ�$���+��7�S��L&������-Lb�2�,kH.8������U����2�^ ���#PW�6��&��!��t\e�U�4DyN��[\�N�^��S�L����x����1u�B�����N��2A>�3���Y� ��#�n8����`	���3�4��hC��˵�8D:)̖�)gس�:b�[�kk�M�gIJ�/(z�ѷ�y����6����]���������Q���
�4�-�
�ؿ ��!\_;MTڻ��(\8w>�ܦR%���ۤF�]�υau8��뎫�/�k���&������G@�i�aF�����a���k��MS\]d:���hha�qP���?�U��F���o3�{�̋��L�y����n>
8f]��G�F�ƍ���Q�Y7 �$�݌07m���I���qh7#�M-W[n������(\���eYtX>�[I-|O#�p\%��P	��B5���,+�^�tY+��Rxz�RZ1oH�s������'�C�w�Gk�2�t/7�� �1t<����8usH�3Ca�"F)���C��>�R0&n�zhQ���Ĉ�ڬέ�H0!��f/�4d�<��VAiB��0Fgϝ����p�z���F�x�5z���}>�����
��E�k#����XNFf0(�H��p�L@?�������� ܺ}����s:8�9!��9F�\b(%������l_�tP��=�I����isZ�e1Lq�Ym�u��F�{�D���jZ%�;w�p������.�FQ�����x��Ĉա�5����wùs�mjX�C��'��w޲)QC�?{��[������ē��6�B�-s�F�n��/J���]��~mv퍏�g<j-���H	[^�� K��q{>/�{/C�,^��D�J�����x��j�Kh0J���ɽֽc��vثwl��<7d��ǰ�x�0�kq/g)��F��Z��-��Z�0A0Iq��	8�$��}�SZ|�"�,d�G�زN7�F`�c�^�B�tm}-��V��3�Õ�o��`)ܿ�(�� z�8�H&l�Դ���_���Ϟ�o��6���?�'�c�~��A�"��Vygw�
N�����QqV�Nغ�`@UVT�L2���� �%���I���`P~��].d�ͅP��]�C ��m�3�G��f�v~2߭�l���k�^�q�y��/]8�Ae%uT.���ǅq�)�;s:,�,e�S��r���#��[�)��uڿ'K�k��2��6���w�}��^FX�=�	�aɽ2L�T�	���K�׺e����|�<a��3L�F��
�A��a�F���R�z;�t�>j�̪�����eb !�rh�*m�g��RvmA+D����Lt�=J�&���{�G�\�LF����4n��hr��Q��˭6����]����x�A���[ao�k(4�/u�9��\3&�p�DT��U���	@�C����:sh�y�0;��7I�g�¶pzE?:����H
�(�:�̣���O~B����R`�*쭭��M2
���qSAK"��P�;{:��ƿEw���7Ѿވ�bf�!��\��7�6�"a�@w'^�%�ru�lil8	�q�n4�.��I)f�#`=&\I,]���b�}�\&��5)[���L ���������Z�j�XM�IM%�JFb����Z�'�,9�CS�������Y)/5����im4�*"��,ayG�������mF�}V�x|���-w��`���܈t�����^D���K�~0��Z��>�Ƭ�Lm���{z���^�� Z��|�嗄��qQP�(��;^9J�C���]$4b?�rNd��3��͑dW��udH���D�L��MM6�Ә͇����`��N�횭�X�,mIEeU+�Rk���p�}��{��p �7h *�������u�O�Qo/����c�Q)�[;��Uh�-A� 	g�и���U51r�ƍ`u������?� t���w�Ŀ��Pk�:E�A��ڵ����f�?�@��9'ښl�Z�x@�r>�]��.w]S!M�C�rfn�f��!�.�qq��-��|s�n��]n/Sy��c�=>v���k��<�����"�g��p��bt���^D��w���T*�n��
۸�l��`��B�9�K=�*���u�փG>�Ebb�y� �޽��:�O<'�j$�`���6}m�w���d4e�n�U�%.�H�o� GK��P�E�I���v�.Ϝ=+�S3!~H���%A���p���l{{S{_�<��<ܻw�|�P��M!A��3�%�IB���fp���5vgg[]�f�Q��*iOM͈����D���6R�Z?��>ӢTQ,Lg���&��
� u��tm��"����%�~�@O��S��y��}���gC�4զ�Q���8�(��ښW�*�|k�jn�S�'+`��-v��&dll
���N]H��](�^-|�mP/W$���|������X����}*��E�l�,�0q�c�<˜E���#@��;�l����g����6�{������g�u�E��*���/c��BN���u��IEr!���T���?(Ӿz�R�>��}9��%��<}���A��^)W�J��p��U0V��o���AT�$,�
	�3��0���߇�`��i(2�P����M^D�?�k�[�a��Zy�p���>?� i��c-��ꛈc���x}��8Y9��x��K�ч�}B�-�`å��T�#�.]s����u�9K�����g~O��m�(F֘�������e/����+T/=f���Ll�gR�@*詀��Ҏ�T��V�ꚰV=G�r��ͅ�$\9�`���|�ǵ�������xՊ��!���e��bO�F�^��A}y���g�s��I|/�+��<)>v�bHU*��i�)+��ֺ�=��@��lmlʣGOh���[�����`�����[QQ���>H0^�a��:c�)L�Ȕ�����>�z�`i�Z�˘�j�w��Jz�[��[�S7��}h�j�!V
{�%Q;�Рlp�F���� ��������穱�=XX�Fv��C�;�����H�q��n�߿�-3�%A���5�#�C8\9���HS�R�3��c�**�x��8���~��4R�Ә��C��c7-zz]��h�qb��u6N�*�4LI�MYX5eo�[̂��oy�a�,���۹5c@�[J%�lt6�}ށ�^[ZUP4aN��a����{Z�s�(:EFc�
�0TYz������	�F�5�͍��c�!����m��NC�7 Ic�%k���U�gL���kDU0O�Zp�+��.|f����=d�]��=P�<�S?k]M�y��&(~VL�sf�|<O��,9a�bm ߡP��Z�/1#\��4S�&�5�5�+��5i����'��U:}j�cl��Ɗo_�FQ�`�&�3��%U��J��4L_�JD��%�w��7�毓�q�1�����H���t6��IÓ����S��Y�������A����x̬U�ź�,*���O� ��<��D��x�^j){��5$�X�;�:��l��1�(Q���bO�ƸY��������!l4n��b'���@lYni�n֊+v�3WH��mw�=���w뜆5�Nb�~)K��6&��RK(3eRO�)Nɢ7M+�%]��z��)guNp)��P���Q<�A�q��S�㎘���Fl�B[�|�Q*��;�
=���8�$�i�xC��i����{��������:N�[jٛ����C�fHs�+�{: J�!���5UV��撱c�����B�䊅 .�v�1�����
��t/�L�)�F��y���[Y�V��,�b
��ոi�3����|jvQ(G9f�ǧ��^����x�ܲ�;V?�l'B�,�&2�Q��n��+�Җ�ƚC̝�3�)�>�;�4��s�"X��ki��w�ܲ,/���W��2�<۲��-o�ωj�NJ�45�a�.���~nl�%=>�Q�qƄ6��{L�;-q�ӿ5Ļ<��}9���:���ּﾉ��*I�Zy�Ն�|_����ב��}�A�Kۓ>��Oƽ��P&�Ң�VC�٩��/L�8p�M�da;.'�`�h�I9��8�V�E�X�Ga':a���C a��(I��H�h���A��䥷@�hiFh���tBꂷ�Z�,Ѭ����g�j�W�}ulfے�t�S*wR�74�{��Q���W�X�F1W��>����2t�؇r��w�嫭�\��nz�L��N�����[�Ź�����
�so.9�
��Ra=)^N��n����fO��{��#�����\O�e���ʩ���Ecq�rh
�/K핾�P{��z'����5�笟��ʒ��x��=��ե˗d~n6b'������׫kaOd2�7� �S�5wӒe�6����s�O�����g��3��d0rM�����щ2bXwE�u�S����N�w�F0���/m�jը��Eh�Y)@�3j͵���7.��sգG\��B�'�7����g���Vxj�ˮ���u�&d�i��e�\]yC���zd5��ݮ��v|S�D�1K�7�4p3��\��.
�ԟKo�I�/~�˗7B���h
hS`�����v�v�\
V8ɓH��T6����ޤ���D�y�=�6u#�u��]uw�]S�f�{/��{)��N=��k�gX[n����a�6J/��;w�� ��ǁ�N�?��ׯn��~O���s�^�Xg?82�j��C��E��< $�A�:9����C�I�n�iê米���O�����Cz�97��*����C��-ƨ���Jܖg�x@8T�P@
uؙ�ώ#N����6�QPH���(��W�E~��_�ĀL���6�'3ӓr�̢l���V��P8#0�`:}�-t*ؕ%mjެtCxƾ��Ć�WU@uQS��5V~2M��.���I$嘕u�r����O
\���M?�Z���]/��h=�k�c��������\U��9�ލ�]<#"y���K�3	�Q��^�I1�������B�ҫׯ������N�~�&��t�,./���VJǬ�$��ݸA���7�p-7o~!�}w�MI(݂.���+�)a� �N�	�QT��
�):b��~�%��e1���skW�)�+�[�7��@N�iZnҭ��,��BD��D��#��]P���/5j��b��ӫ5o�~��	c$6��B�=y:h�ɖ��3L�X��nKΟn2'j簿#��9�8ܚɠH���h�6(���+��r�R�G��2�RV:��e��Y�6�e�k\8U� �W��2n�t�7�kMK�n�T��ҭv*�i�b�OR��6�D�
FR�O��1�Ք����=q�����{�J�hJeI��8�xdf|��p��:b��>�LjE'�{����w�Blp�v B�&�������ݓ�ѡ���ZA����ˇr����[Vq #�,T��\��?��3Zp��r�	�"�M����]�j����}ƺ�k��|p�}
ΫD���C�`��� ��%���,��ޢ0p�V�	���&)Ȁ��8�ʕ+����O?��Xμ	B6$�ж6�v9���A��$~����\�e����p#h�Uy��%�ϖ��Rg�����2Q�A��1�]UP�Yf.^�1�wE=s�
m*$�h�I��+3έT4�ܓ��ϥBь��n�
~�'��ib%�4~����� N�����d^*;~�x�3�Xm��W����j$UId��f5���v�ͮr��5���%�#�VXeEgt����.[�ۜ$��L-B(�2�Ls��o@s����2/�,/^�P�l�M�}eA�8�Lq��܃�w&���"��b�8jk�+2��+4������Ik)�u�P���*�@{�	@�]�x��/ Pp�F@� `���/(�����tfAۨ�/��˾Z4Ň� ���B����ʵA�uC���K��{�����33�7')w�F/�qO����.{���Ǜ��O��b��ϻ>��H�y�T���a��f�p{/;����^�X�]I��hziҵY��d�?1.4�n}|�E�a�-(�J�V߼yM4��d��sFҍl�؛S����w|�,b���Ӳ\�?��O�X����IP?y�X]��� ���UUX}`��VL���|:'�H{��j�]G�V1ǎ*t��qB6)��	E=��y��5���F�'�{�{Zn����fzz.ZtVق�B)��sP#��H:,/-<�2�mK\�<��8��̜R?hј,n����L�{�'	�I�:��ǤN�����{���=�<jA�r����{����g*8)\4M�5�g��;Mn��E��1�Xy��?�������<��j�jޖ	>�� c����-bﮯm�P��{{h�Y	^� ���<|�TVV�%�*��d�z�0l�����{��qB���; ����3��d7��A��5�N��r��A+�.@�9W^�,qo���u�p"`���<?7\�	� �:��҃Cu�=���}m�[]Y��=^�[���e-��ٱѩ���Ne�X_[#�E��9��C=�c\���l�����Nw��H��vCLE�5��6��xbFj<��Cs~��@�p��\Nگ�8'l�tCUU]�I7�1�v��c�7~*<�8۽�f��C	��k<���IY��pC��@z�Tp��0���^�+���*�apzܤd'i"�^�+ gD��k����:�qrj��zeuS��ǿ��u�~?��������0�.˥���L^\<%3h��'�����Ԅ���d!�� $ަ�{ث��w�u�bo};����b���,�����8��lY6�v�b��8}zɦ��~��~���m�Eܼ�����dC��ڹ��L�皝匭��۞.���h��L���p�����nJmlM��.��cq-�6���ZWg5�i���7q]*����M�J�;n��!}/��5p9I�OV c��|�?�����=~��s6=�Z��5���r^��w��kN�~���F�2���2���\�pnknl�%�Цi19��r�>��w�uѯ~�+Y\:%pF�9�ٰĊ����۷I��6ռk-��8 �әa�`�΅�w�^���)�G��,7�ڶ��il��c=ɵl{$ð�������9Y]�q�S��l���k�z�U:�If����B�W�ȍk�7m7�gL1�U��nu���w(�&�ѣ������k�ph���ZF��I�	��[�@]D1����c���=��c���8�>6clݠ�Y��&O�p��V��eO���n��sM��5���Ͻ��.%r�0�dck=)H�oڴ�i�5��}i�Q�'p���'�b ���G酑�	V�y�a�;ES�p��r��ÇAf$ke�b��ޝ�l7bg���N�>|��5�?{����1�w���	3�L���{��ظ.Ժ������^�[�y9K�(3!3��Z�˫���yQ�s��,d�P�����$-�ܵ������7#��Tt���"���=/�*�}�����Ԇ�N�����xV:b1�{�!
��0\��{OH�^Z� 5:^�a�%�@.h�gY�;ءi���{'��f��HzXh�*�>��O_c0S�Bi
B���Np�S!K����鱎'�ƿ�\G�J�n�a�M��n7��TR���'D� �)��=����T� �\�s�d��ׯ�p.0����_&ׯ]{��_��<�A�,(�a�Vxh�(@�����T߼�9�W<xp_^�~�ڷ�:�w�>����V$���Y��(+��Vs!�:�����I��.{�%g�(#�d�1�_�2@�L"�i-�l�u�>����+W�Q|ċ���^�ƴ>��E�LL�xS8Q!ob�|E���\�#}��2Ln���5��1�Ξ�^��xX�#\?����~���}Zwq��Ub�8;
����M�b8.?�����3��I�j�lR�Kz����ϫI\��k>�����N�ᕒK4ÑT���y�Ú��6 �{���V0TIW�(��m�ce�:�#3�I�.�f�ǟ|�,��g/��,����˟�^0Fw�ܓ��(x I��`��
]��c/~������׍f_���-z�)}3�ᳱWC9����9d���RU�a�$�癃l����8����;�JKh�[[�d� �66��:G8��Q=t���x�@���H�O>�$�Y��A-�醪袀�V�t7�ݓ�������9���<Y+�B<�м��d����ms� �O7J����	$��j\���M�)���6�¶�KqW(���4��ª��)�~3O���b1e�{������b���Μ�+nmZ���I6]GӭnS�+�=�<����K��N���>M���EV=T3���>�NAD�{��pD��G?�)ۻl�x��5�QH�"^pre'V}���)���,j��K�����L��\ga�@?�O3�CG�����a���0��\jБ�v������K��Q(o߮�~p{J>��fWj'���` u�޽#��oɅyRE��L)Ւ�C�������r彫dW�"h'�(��?��>���Ç� /��D9��>s��̾�
�����i?�EG�v�� �q�� A��E��Qō�)q�Ħ�Z��Vſ�twǬ�1�1V�����U�4ѿ�T����{'��M�}�:d\9�=�����������0���b>3UX�f3D������>6�u������*T��yf�g�L��>�\������=������/y��r(ȚN��a��8���}�r	4������M�_�C��
/������S�2\�����;<R:as�tN��a��<h9�F���{���}z�	�����v�F�k�5��O�<��P�LM��9�_���l��������I����qw��ɼ�y \�rV+I!1ǖ��>�Y�i�-�i�'eZ�c?���ҍ|�W���{Cx\+4�.c�>��:-���6�k����>)dh�M�#�$�
=��i�*=g���v��\������vwUp�96v��q-�0G3�4�	��<���c���j���8qdاb�E�o���+<V�����
 R7i��V|��St�[��j���}4��^ƂqK��wu9 ��sy��]#�[�UZ�S��Х��9����
�@�2�x�R�Giu�����/|����轱��t>H'�h�	��6�{�\�9'��>�]��}��tld���ĐD�i��Y�q��]q�:Ǹ�4M�����܉|BG�9�jR( "\��!�tC�e�:k�'nZ��pԂ7^�n~�����@����R�w���&]�]T�q^?wS���iȐ�|c�	�&��	���_C�z�}�JJ{�\����9�$zmd)���Υ��N�zH���H�A�q{��W��0��5���M����1G3��B�T�bNm͝߻��)p�尉�G]�K�uF�ț84dn���(�J�zd�c���)-���f�W!؄��Tr,�F���������L��:\,~_�,���S����Xt����@VW�d��]m�L��޾}bޡ�]\���T&';���0�*q3�	2d4U;�+��a��"PB�:�$939Im,;��Ӱe�\�l�l\�.�Ղ[����N�H��>.Tu)�$�?g��4Vn&�N>}�q��Ins���+���5��M:M���͢�?�4�C*1�tJq/��A8��m���_�F������  ��IDAT���W���!�/�/=�Fz6��@zmnmIA��`+޿������Ν���z����	F�_�e�Ex���VfZy��r(�� o�J�~p\�uB������&.��젏��vw�'�e<d�u�H�Y�% 3�Ò�H4������&qh�_��7D���cT��j� ���EG�hj�����8"�.vav!�9S$��mFS��f���P�G^fQ����������p�V�y��lon��f��{�V��^o?2LHV�H't�Y�	��w	�Ip��?JV5�W����>����Y��"σ�	J��@R˜3�N3y�����i(�L�����D�?�ȝ�ei�����Ypx�����J0�utJ���n�veM����d���,.�ek���y��U�ZJ�9W��G�;���3 A���B�	3M,�=����vVCSlY�.�WJ���ŧ�:=�5ಋ�&*+�d~#1CWv�`�R�"�k�^����
�n��'O����rf��|������&�-��hRFi����t�p@˼���%�
���'�Nh-�A�cJ�)y�'�^����)ؘ�9,;!����}%���I��xzYΜY��p�B��lsK��U��
�)���wnjю��'��n)}�����.,'	v����'��Nr��Ϥ��￫DvR⮩ ��;�{��kRJ]�n%�aIݟ�6f�#�;��B�囯����s�K����L��G�� ���?��<���w��>D�[�(�rJX.���*�2�YA�� ^0��=d1�@T�ʪ�XoRJPA��ᣃ��Ӯ��Pe�`i�{X�PյU�W�:ʝL���X">y��{����(pp���X�s�Aa5�6>�N|wUd�����3nR��#�9�ܐLk�H���ug��:�7-� ��?���uK<X��A�u���.ݣeL>ҹ�Ќ�Y?��O���3ը^��ߤ��2���.�I.�?��b����v*hM�;uc����Vތ��	bU��?��'���(�䋱�\�L	�x&Ȭ���ؽ����k�����k�'m� �i�ɔ6�c8����:��B���~8��8L��<<!�����6�)B�qrUJ,�*9B'&�� �b��{@Vh�;��s>�}����9%�5� �d�(+b�
	�n[I�+ޠј&����D��1A@���,�be�uC["�t,à�֘)|��1�do� �����Lf�3��m���j4~���	�kn��UU��k��A|���Sv|9v�����͊|��}f�A��|Px0J�WD��Δ�řՊO���u� �{���7����<���N*?v*�xU����}���z7ofI"��e�q_k���+��w�V�Y9/j6Q��[���-f|���ña��C�GJ� ��t�\� �|cpTҸ��0H�n}%� `�/M�?֔u!.'x��V]F�t��g}:i��(�V����]o��������˙�4�%���v+-�e}�ߙ�:��.��?��r��}jLND��땷+�<����QМ!��(�x6�=~�PO#U+>L���6d��8q!u��o��x�B��/8�� V�<�[�%0� ��~��ʦ��Y]��<��b�M%�8�!�����Y�B��70oϫ<�g�^PܸpMK��*.ű疤��( 'SB
��u�2f�z�i�Z�8J.�k��̒���N�3��e�,��Z�3C�s�FT_���z}�	�-'<pi�5�E��)������"f�~�8�a%�'����x^߯�eb���W.pN ^���p���}�`Tɵ�F�]�BR�Ĺ����-L(,�͢������`lkGI�d����9�A�0-0����suq����eB�Kak��� :�F7hc}�?8Ѩ,��6;Yt1-ރ� �EF=�Ba�1�y'tG>��|�хp^e����Io�W���ґ�Җ��h�f��7GP� IQL`���6\1�Zx�Ȋ�KA2�2,uYZb��N&e�q�Ut�mK�X<D���ǰ�����{b��� on3Ȥ��1�J��
����)
*�o���:-���JBT�� ���ה2�f&йg��cpeP�����
<�vh]scT�G��a$����@Ն�ʌ�K�bŤ(��M�[��Gn;�L⌽y�X�����/��n�̟�ӻ��_�V��r������K9<�_����y���
H��ک,+z��/t}N�����w�="g?�{������χOC-��mR��l�Ef��H�W�iOt,�����SZk������8���h�����Q�9j�ᆶ:�\����3�>ȌO�'D���pfI>����^ĹB|1�	{�[<��@�-��ɯe�Rf��<���M��2��H,��56����i�[���ۀuKd{j!��vj��,�[��dP�Jc�f]7��2�Ym��m�<
]bJ�<&��ɉr�,V�L�����ii�ϼ�*Z��5p�����׀�xb����R��R���Ee�R��k��"kV��uj��������+���--��B&D�}��ט���ã���������̛�[���mQ���B
����J����}��?4��i��g��^�2�8�XM��l'?4�S/���>�}Qt$�T���HԱ��>	&�5�=�ȭ�M��fT-��q�0\�b���<�
�S���?��?�����dnj&Xo�Ss�r�TK6�^˺'S3ĐҺ���-ć7b:��q�q��d.�.^�Օ�������F��m�Nɕ�Wdvn��ƈM%�*���$�]e�(Uj=>��^͒�XL��a�n����(mOܨI6�2��Ts�D�U�6.�T��3;�V���ײra��a����k���H�ٹ�����Y,SV/o��aTO%�8�v�N3����QZY�?�����p�l�7�]��n+���'����`��=N�?�X`�q����n�*ͩS�$E��z������a��r��9��ʰ�kk�U�jN������^����'�"����Z�t�c��Dǃ�kNQ���B�|�}�=I�	n(�LL�Ị=VA&Ұ�P�wِ}!��-���Zo�&AH�;�3��d�;-˧�z��P?����`��A�f�H�L���U�8�ʩ��+W�I�n"�`H`tC<�v%�µ����ǟ|,��50h`�)�\�B߶��7oࠋ�Z�O��>���l����\�Ud�jT bi_K��C��y��S���¾+ٱ���a8b��Z�ns�D[q����8��x�br�#(�Dw�驘�kL3�̞gz��s������
ǭ���QɊ���Ū��P��e��Ş�L)���76���1���t=�}����4��s��r��� ��Y�E�"�M(��z�8a/�ht�������>59M9dHkpPGqz��	��^pX0�6�j8h����7�c�C��B�;n�a��Fhv�����@�f�RO����=Rn��u|��X7���K[0�v����%�~/���ت�iX�����ϸ`)�c|>��S�?u���ai��s���\�4�0�W�$�y�VT|���=��	���/��и�}��q�3+(����;��'�K7���W�4�/?V��if�ݣ/Q�z.�ݱ2�B�q���+)��F3�[��Wz�Ve�k+�V1�q��2�H��ߔ���zɌ3�I!��,���J���7�����N��[�����v`��Ѷ��A.�w����w�~G~����C����i@��j�I1��VeV�u���&a�*@�[^v�<!�^\Z����͘
inv&��3D���Z���B�o�����@�
��i��Ӣ�~��{�:W�?{��^#�-����u��k=53�5�??����AQ�ۆ�&M��^ V/}�i�G"F\��U:�/g�����3��|�p��n�����-c�p�z{ɧ�7��c�w����N�J� ���Z�+���4�$a�N8nZ�v�N=��?=���cפkڬ�*�_J���b��|�]sL��=���*�Lb{i\k������P���R9kW��n���ˋ��S@������B�xj�,�=Cky�����a���O�j��n>��f�9~V*c��x��%-&���1�5�^��>闒ѵ�_O�WZ�hf 8.p�N��+�-\H�k�r{�G2@��Ssh7��fi�ُoܐkׯ����H�^τ��8��l��dt�A#����rt����З����15s�����Cjr�"$��7��O|C���٢r:
�ou&���J��.2O ���P�]6��O{�V�L�'oF�[cD�Q���L���|̒f��Z�&��f�c��.m��*�F�"�d��J�ﲒzGh\c�(L��\2K��w���d�o������^s�)B��x��<D�n������*��pYȨ�]eeD���:�W$˯j��r�?��`#���_�J��m���|�#���?�_�ҹ\�)y�2��F�ȁK �	Jckk��(3%k�|��p�Az�5u�0v���,)�֧�g���X҂E�,2԰�(Y)�p7l�)j4@ �u�����(�|�Hu��_�pN�����������xZ���4\\e���(_�|�7f�-e!��5���<�W�:��%���B��A�-�Yi��^�ȇ�����\G�8�m�����Ȳ����f����	���FBK?u�H��t]�4ATkӪ�ߋ���pV�
�qg&1��<�/;���L�ƪ(^����gy����M��mi+Z�[`a�,��`̾"k��*8h�l��,5�����V#�pkO��u�3��
��,�g�r:�1$E�����w}Orz`�ٱw(��Cy��,-.�(�m�@.���Y��Q�{�
���n9�Z�	`N��UΡ{�ɓ����Kk���apGѩ85A�W��q<Pd����HQs��Jw��F�!N7`.��81XX�6�������*�A!�i���H2]~�
52�3I�'��Ǐ��	�j�wb�����~)7>� W�,ʨ�'7����\!��r�P��D�G1i����0���n�Z`���(|b���OK�q��U5�H�丞Y�M�\�T3�:�KQNu�E7}�U��V����IpCǘV�(@�+�j	��J]���nY��ϯ�mpE[{�NI�Xj��C�b�<��R��J�k^�fʫ�{��@'?��?WI��yT�y����Y��9��_�����W������!��*��u��u�bT���h��7 K:j�t&ZB��5#^����v�3E�Ȕ�7=އ1W¾sg�Q�|H������4�����E{���	���3���BM��q�&�6!P}��3�)�f����AȼtD_|��x��PJ�K���W��ۿ�
�1�؀ �d�Jf���)dX�q�NY��m��<���69ǁنrҁ�yD�a}&G�V��9�W�+�d8?���EX�Z������~�fE�16���PK�dVg�g"�n�c�� &r	1�ݍPI�le� \�f��[;w�9f
 �.�#�B���˝3L]o_k"XQY��[�0��ڭ��	��-����qJJ���Z!���:��L�!�	hm[�����ٙ99��(����%��ߘ�,w5�G�!}��,�:�Ӯs^�QRx�3��F��̞�l��72�Z��1���sV���rQ�̛ ��s�l�<�<�Y$i�=G���XP�P�:��x�Z���]R��!΅��X�bG��.������bf|�5,0��`5x�d�2=�WJv�T2Gm�d��O��g�Y���\
��a�%O��P�7VQ
]�)5Y.�QeEa�7f+��r��"�1R��1cΡe���_���:���;�����pLК/���_�8*,��'J��%�jK��[��c��l.
[��>��.��[���E�Zf@�dUR<�;�5�T���Y��Jx%�#oK���+�.'�U�U�6����e�WX�������\0ck8w�CFc�jɠ?����:���715˱Sd�!N!gL�=�u8�·��|��-�����p	�/����p�3������U�^���5�H���ady���PO�=w%�k\_��.-ֻLz�W��I[$$�E���v'���I	�~=�[pm�޹��Š%�HX][cY �c�c=$X@oD�!�§f:D�@���
!no���g��ǟ\�m ��H�=]��[��<dƚV�cT�w0R.e�̴<��B̲T��%-Z�6�"E��o�&�2+A�m^1�o���ٹ��9
 ?l�r���f��enl;�I��S79��xn��J��f h#U����Y���6w[*Ǐk)	�m��Q�#��cJ%�04����!�4���m��?W�΅��A,e�x��Z�g�p���)��~�!�BI�9��ea��+�ZCӌ�n�wbۥ���V�-�G�P$��3����'��3y��fSϜ!s����[���m����3d����H2(��327�����K�{0X�ޙ)���]*���O�-��1��#�?���c��_S�g�\� �5)F��$��GA�1���ZtWa��S��$]��DN�`���f��q�y�هr��y�����^�n[����pnL�l˩����J�<�p�YU$���=�PZ&<��@��f�3S,�d�.ni�njVF73e㈵v��A�����(�-�����N��>���Ǫ*[�(Ƶu�����$qa����]us]��g���mcS����Uh��G��������]��%��a��f]s�^�Z1٧���!��SW��wj�Xe�^f?W�BLu'&�`1�'u�r��4�����OOOR�������󗂇8�\�%������9�`=��)�R(@���1 <9w��r���^���>��}��k"y�$������x6��߷z=�zx��7)���Rǯ�{f�!��c�0	���V��Fk��p!�=�F�w�ڵkr6��mAܱ��,���?�� D��[Ig�6\ 1 ���>�����!�B FX�ς+�P���tfQ�[�҈�6�v�������
���T��A7�
��	6��JUV7^8:�]���31�Z'��"i�hY3D��e�8�r���+��z��ٲҥ	�+?���$���^�	r˔���Ѻ�xO���d�0� �Z��\swmTL��ڪ�NA�.te���!�]+�I���� f��I�.qeJ+�k+�sI5,bp4J 硉ٖ�?�6ަg�Ϝ����ŀn-,2�͠���'�5=;#7oޔ�?�e`��l��x��������45��{ �=}&�˧�
��V��Hh�E�	�&��;a1}�^���j��y$��^�C���W�<^�� Qyk���3�2j�͠50z&ߧNq�^�5!{G�M�G^%�p�ןl0!怋˗ߣE���{��~��tM�g1+�E��U�����w�/��L�c�N����to޾y˒���Y�M�u���&��Pg�d4b�~�;&�mk\mB�u\9���Uz����-�;���r���SeUĸ�0�J{d����N�u4��k�NbJ���yÛ��ND�s�i/"���=5aL��K?�+Vh|��N�$٘�2����ZeK�rT�Q��\�(�z<�(1/���ȍA%�eɫN[� $�n`}J��yh� �<G���=͑X��Ɠ�3˴�u�	[8}�J`{oW^�y<�-�NLq �?{G-bO���Dμ�Є+�Jp���}�bX�^���5�ѣem��(���m�uXa�U��7F���e@���͟�Ɔe����O��y�;M=�d�NZ.���H/�+�s� g]P�>|D�����
.��ꆓk�x��	�Z�z��d<��h^vy��pc�����Y�"h�=f�����0��vm2�e�!�]h��Wf�6�	u��,	���2!�B��8}�G�u��Zj��)�&���Fs�d��� ���s��ܚR.�Z�3j4��H^w����ڋ��ǿ���-����ű�hZZ������*(zG�KH�Xi�4��ng"&������x� �Ly�r�?h�2�Q�D{�A�k���!$sgQ�W`
՛�9���yX(+���
����KN���X�)YX<�u@��x�����1���>#�~���"�ʡUW��'��Z�_^ޫ�AH[��P����|�_{��o�e�޲#�<䢡i1z�L�����Ġ�gd'���^���b����r3�mQ����}���x�<߿�����_�/�+Ov��n<�Tʞ��G\/h�͍s��]��8�zii1h�u�r�3�<Mp���8?7CM���w���j1�͐PC�,��NH���&^�q���Bg���Ѩ�	ϙ�WkV�1���-de�εe��!T���y��s�h[L�{�;��%緲l��F�P[}Wi�2e����� �6��*�y�ƶ"����{M��	*߼�VF�0J��l��K�u�%�R;�ʘ�h�<��8֒1��,��3�LP!dC����?Fl�t)��ܕ�_�0����7�� ��S���3�`a�����\��`�I�����\�TDMa�#����$+�gN��>x�z��00����0�x����Y|LH��m�VD_][}�8	$�]�xXQ��hG|��N��8\��Gâ?}"��^�|1X��������ܓ�Ԧ>2�!�(��F�:n�䰕e�v1��;��u��-���yC}j����{��L��ի��1�ښ��_�3.�������Ծ]��M=g��'#uj�XsW<�ݫ܆�WJEb�6#e��Y�Ҳ��X���R�z8/���T���p��F*��?��H!�X�)�J=�N��
M��8)��NmzR:Fã�����m��
��b��,;M�6��8�x����l@(mB 7w����*����v|W^e p�<'Up��Ë�����H�	º�����~p�2F]_ߦFٵ���������H�C��Q���>q�۵� �=��ڵ�e"8�ev0�����{@m�n��B��zzEf��T2\#x̊�Q�_�n��<^�D#OZ�o�mM�M�lz���.�z��r�d�V.I_��p�d��8��r0��r�WV�@bZ>�|�@/_�,7��\�7�s�Sc5Ȑ��
6sp�0rmeM��SX�J���	�n���%��������w�ᆧ��sȡ��+}�rMvv�YsDC�k�Jr�5�RZ`\�5a�;a=�~G�N�����	7�5l�dw� e%Ɉ�	""�a������\!�,z�@��@2�AC=\C���?_.���PT#��p�������}1c�
m|S�ꀇ����w�X"����,��8Iؤ���(fM�Yւ����3nī�R ��R��舀�4�otϡ�YJ�@��;����^�Ƞ��V�Z*��Oؽ@vY��d!m�8������o1x���AA�g��klg�����E��Yb<{x4���pm���k\J7�B�W7�q��{$�[{a�=��w��KV��q#2��W�@�W����3Oku���`�t:UT�r��	m΋�\lm�p���h�D��� 5���˭�VQS��G���۔5����I�E*�\�<���� ��Id8۳��b��
Bq��{r��5��r���$�3l����.�W}\�YN͘�h+�r"�[b����l<� ,���q�fp����k��p ��XY$x���_�dP�����mfy�j�[\�x $��G�>7�&���|��7h"P�������r ����#ZE�`��S���|VivP�:�n0%m? ID�=Ae{��kTTT#�C��Xo{�^N/���K)��~�-em�
�a�R��2b���P?@�gJ��׉���{��pT
����a�,I('H9�����Ua�F�&�t�	Gݠt�㷶�8v/xvY[��:h�癙S�0�9̮,�-wBk�hO��eb�3��5
B���r*(�
>�m��7K��9��J��P��@R�[0��feC���[{ޢ��Τ��������J���@T1K�����v{oo�.�z��Ѐ,��e��ڊ`��ڀJ��q�c�i8��#�!`���i"+��enme����2�5��],q��K��&������&Go�'�|�n�㪸UT�늬!��HPsOt�����h�X�2b�י�˨���B�?xʸ
�4�&)��ᕕ�`�{,#��k��7��W�C��~� d��g�����L��s��+����{��H�/��B��:����~����m���k)�2�4B;�2��,)�sA�0yQK����#V1\w��y�s�^cS�M4
f��#B�ik��k�Xp���LZ'��p��l;��=<���˓�OujDr�j���L儃�6����|35�H�b@p���<�I��Z�8�o۸��.�ˎ��3a��`Tz}�AG�ʖe� -�7_���74h� �u���Td�y�╅-9{�ܸq���%������u��NMJ��/���*d�;߆}�oH�6�s����|?�~y-��y��b�����$��0���]��Z�@���d��|0�g@{���qR�&�^�j$�]�隮�������ƴ�D�L!�r ot�p!�Zy���2u�5�"D+m���ݝ{���fz�!d�q�����d�]�Q���w̴��A����s�K��+���nS�sj_���ͤ��3�!��7�zrh X/�;;T�9(���F~�� &`Ӑ^5V��⡅�t��*�{�+\��:�vo�0+f������X�3�u��)㟃e�+�>ފ�n $uQ6\[��tp{� �*Z,wؚh���D�9</�Z9�Y����y�X�"�`^��V�6gtr�FBq�T��
<"np�k����VZ�q��"	vC�H+�R~<&�Dl
K;&�N�ϗea�<FV��&�[�F�=/�p��_3�����׃�{J5��߂G��?����eFxt�;��f�K�:�:�otj��P��j2�V�g�&(�DS,�$�{e��VYi�E�Y�ts0�N(#�]ݍ ��>�5CW�$G�&Frռ��D2nzfR.]z���x���\�Q��T
�'�r��C�� �!y��r���~�~�=C�)dvz���(��[�l���tURq���3���)�V�����:ԙb��JT5�L+�%�u2����:����a���&�#��9��ʷ�):��s�`.�b%���08�S�-oe]ZLo�d��Q;Xi�OW�e�$�ƑXYL]o�����Qn�#� v4��&WJa�)$� HA�E�{�-Yh�����^/�gts(F-�k�����#L���
m&R������ۏ�^���%Ƴ,5MNQ9�΍���p��ܩs���P�U	4�T����Xx�n��\c����y��dM�S���Kݦ'y}�DP�'�`���0o �SX	�-�ӈ�h|{��0A=Y���8}�k�(V���qR����T����2�N�x��έoT[ذ��\��aB�0�crbZ�S#��P5۬�]m6oPi}������]C�kdN1����:��Z��+���ų��CZl�3�Kl�zq� l�����ʁ�о�t�F���9c���!�p��E��{�d��D7玼z����K��ᓜ������;ա5�v����-�^0ra˨k}�x�ٳ��uf�KȦ>`q�9@@��7d-�������
8So�m0�݃}y���h_.�����(�S���a=��L�{���td��Ϝ	�L��G�a	Wh���7oW��Dh��3��XW���w�8�ackK�̎f��z��:j��0�vvmػ&�Jc<�N��̄Jť��ro@!H$�]]b.|��̃�*��B�)��ͯ�Lp��$�܂VOZb����-��o9���-���oֻ�7˦m�/��[�\j�N��I�g��%b���@L|���ooߦuF�۩��p@F�Q�.,Q�<>%�G�`�Q[u�S@�)�xfX@jp�Y���e�DE��-9Y�im:�j�5�C /������>
7�pO멜<����ѣ'�~�����TD$�B�e���^\��:���f~��5�Hͭ��͊��e�!�E7V���C> �}]�9кw4��f�rp!���9�,��_��T	'X��Ü0 ���ɜ�� ���l�A���
+=�Rg;!dBu 2�Zȕ��R�B�b�s�"�;{�D�z=�=�z~P��zl�̓m���Ӳ|�|d_E��$�$����~x& T �G�HF7(ҋD(�B�K��.��h�T�k�y��N$� }U�����Ӑ �fF�`$>�UX\��(�y�k=J��I��%Ǟ���9��pO���?�׿�-'�:���E�!���>R����`��D°,fy\d��3�_�\"�wR��[kluZڪ��Ļ���jMQ���*�p�'�˽��qF5���Μә�T #�y���L��E�����͂F�gvv!\�!#��%�aXDJ[�9� ��Eft�Պ�!X��@��iɡC`���>k�K�:��s�.6�qj��Hm�Y���e/X��U--�5;�F��mo�«7o�&3�K��TXCKU��������08O2��;ړ�։CZ[�byd���|H2=l�/h> � I��  C�^
�B���F̊{�����A��{��/�6d��s A����N�����n��-;�f�5C��aOg�e����$���
V��"����}�������NX�.ׄ=�2�ǔV��=7?��j��иZXJ�,����ղ�Q���9���\a��ޓ��EK�rUX�P���,B+�u�*C�=���0���.(�%*<�o����)�8�
%7T�X- �v;�����a��gJ�=$���1�+^�`�����eh1�4�@QHg"g�%ԭ����oB��\,�d���o����d>�$X�W!��:J��Wʎ�Q�hFpn.�c���#� �bh����2�l2i�1�&��|к��`���=zPd�>� (��(�L�Pfj�c�].�۷�Ud�*+.��{V��.�fp�q��7Ȁ��=Q��g8ҡ����=���y�m+(�Αr@�l�oS�!#!��efvR�,�� �6`���{�0�ȓ���Y\:C�����������5�c�Z��a�P��3f���H\�t�����L���Jk�|�2Kd�AY�^3QL��+勺Į��'Cwwgk��HB��ǟ��BJ\<�V?(�]�J|v~��¡�)*#�Ğ,F�4��4�CHb/�b�t��O�M �.��/�Ve�d3>O�w�ne8)�꼻-��a�^�KfE�V[�c�5!��Y����'�x9����Ms���<a�PVB)���\h�8�y�,�Zn����7o^'��q�(?�����x�|�/\
�9(��m��g�˅ά}�0@>�b��x�	49�8�3�@k�%�k�<�����;2�*�5���o`�!�8>��C��A�,��	%\�� �`���a3�j�9{^~������R�c�1H ����2�Ϗ�Lj	|�����}3�gY~��_�׷n��w;�w����f�/n�����Νoy\lp���/90B��K�����7�����������[�kA@O<J3O=�;���������ܽ�P�YW���e���M�����G��w'��g��s*���_1l��xqR�����M��7���`�φkC#γ�O��J�s!��" W
.��{W��h %JxHB��?���DC8�٩�� _��mޠ��i�h��Āw*�Q!�_����9�9�z���'� t���A��6K�8N�������PI�8���~+?>�0ڊRDNI�,n��(P����$�XY�:yj���(Q|���aQE˂i�h8P��Ԡ� �%VԖ���~���߅U�s��8�M�'��'�Eb�����A�X��#G�wXǇj��&�^ ��[�+%i@8��	P:�;j��7�����ɱ���t7�cT�gJq�� �<ʺ�g�k�2h�'�9]@P]��� P��������Ϟ>U�s���}�ׯ_
k(/_=��!��y������,��B����ާ�� qx�Q'EbI�[��e���a��_~��@�J
�L������K����t�昘�����G\׍�?"ON� ��]�6P�~��gTP[�rj�t8Ǘ$���*Zk}]^��}����G�q��*xT�����G��g(�������э�壏?!cɣ�Ϙ4EH����R�q=g@;�6W�O�� ��@�(����1Ðx��h��[���~UW�2�3��.�!j�{��sX�@��ÇyLM�N�1�r���^W�g�y�-!���2�9���J�SϪ����pAh��:JSZ0�R�������}���׃F���xh:�2?��Ϙǃ��!�T�����HS��
!~�, j�����{��{�t��"��"��+�,n ֡�}`�; 1��^��3烠^a����B<�g"iL����$Xu��6��C|������QQ��2N���Ѫ@؈�[�^8-/��[h�E��8��9��N�1�L�����F"�����ΰ��,�ֻ��f��N�via�Pa�#���0kL4���ameu@e
�ƍ�ȇ^'�N��f��+�L8�d
��̥���R�ֈ곲y�:�r&X-<�+������H�B�B��{X(\���!���_�J��c�<�?��O�����d� f��v�i�ouHw�c5b� ��P[��5�{y�|
���ು�<=s���#�p��%933'�����D����T"��-�,)J�Њq�+���F����`� ��Z�Wh`C��$���H���l�Z�^������{�����$��@���f6Z����,�T<�ȷ�&��/�y�%sC~)�\�Q�(��y���q�HL�4�&��2a� (+6EEz䮜Z�1)�l��(�`9�lonm�ɥE��`)�B�q��D
�n;�%�w����H�`��K��zmule~!�T�j(��sa�/WV�,���j2��P8ǹ��c�^�����Ef��pYW�;����pG����uCi369�rP���/b�D�/�[�( ݙv,MBI]nk?l:x"�/^
¾@�F0�P=)(E��>��3%ӫ*��r�C��͙�1�Fa&f��0��^�WW�������8k�^gvW/�S�����Q��z�a�$K:��>���݃迆b���I4�:<�C��j�%IF��1���	'
9���g�&��q8�㿩�9bC��aX:���0����Xkf�ȒNzS�QqS!��r:̻ �������h���_n	�&f���S�׵"����<��YQ� ���B1�����WC�yv	+f��[J�c�ݒnrw�elzԯl� �a-}Ч�=lt�G�>�G34~4XK�
��lʈ���!C����Yն����ȝy�ਡ[��&����(�}�b
��'�Z�ĴS�`��,A:G�9�\Pt��|�J��:-��R�u��W�}R��y�{Q?F�
�9�)-�X\Z��Z���*��X���7�������.fi���o�&�,�Z4{�م5�K��h�8p�}-@�D��*��q$���<d!�A�ͼ�ɔZo�����?`��N����!_����?�T~�O���&������(d4`:�U��p,�!` z�G��l��)8� 3�d�B�$�O p5�T�w0!H�c,j�T���"�;dQ�i������W�1Y6ў�����c�s��eܛ���+#/оi��7�-m#c����4�#��m�9)[b�Lxb�������83�ա�@H�1�0hK|g>X��e�,"���i��Y�0ff�٥����aw�~b�VUiYpscK�V7�BAj��f��x��"����3�����T�POGI
VB�:	���N�V�E�6ﵫ���o$a�x6�=������U�O��L�t�R�⠯����gPm#���VO6����A/3�*[��M#��2�� �G���Wũ�!��c�o����B!dB"Е�5�8�����׬�z���튯 �H��`hl?�V�hY�Uד�O�CU��`�����g��tt����w��W����&�#(]�Q���?��"�w�d07No��E� ��B@=7�0õ Ll3n��8^�n����`ۛ���{�{�ɉ�L'��_8L؄L$����7�X1��܍�Y����tۄ?*� DiY�ɢ��AG�P�=��->;��Ĵa�$;+'�S�K�lK��� �78�[Мx�Qr�zB)��8�d��2�
�0�+���6���(a�X2�[cn�H�?C��E~���&�TZ`i��V���ۛ�zC�"c
��$�(����BX���O
kmsC2�6(r*c��%�2΄�����n*�fL�g����q1�
���gO����6����6�5�2�_0��ڢ���xc�b�<�r�{��A1!\Z�
IDf�3�/�E�Q�?Ne�U�UB�b���Fc��������ש��p��'z!\����� (S�J���\/�s�XBO�BP�ǽ?8�c��#/ �J��l��EI{H��]�z=kU�w�F��8���͙R���@�E�=n%�Y9Hku�$�~R ���N��</A��S��gf	�T���m2bY���U�Ff���f��Î��pH+��p:%鉄H41�"xa�;j�ڤNW43����OĻ� ��zi���L������6�5��_����q|���@I�7�����;�����(���f�D�:��.[+��!��Jnِ�_���?�'O�FH$]x�����g@�����~���Lp?{���A^ �$�!��Qu��ْ�`����Z���P�=W��_0������
����
����[Z<����Ņ�,��W�o�l�&6;+k���>O�v������q��E�ݸ�%,wǑhC����y��~�	+3�dI�b�{��}��y�O��۬`@@UIl�Y�\�d��^`�����(��Y��I��`k�Ю9�ݧ�UKz�{=��:KZ�
YۧF%�\�ps�]�6��ͷ��&/�6O���뤏�<��� ��I
@I����93Qot%6V63�b��ǙJ5�No<�CE׿,�;�tl*�v�?ik�r^c���U�U�a�&������|�R�~G#+�i�';�pV_�bϡ�6����N����A�\4X�v[g����y��� 8n�^1�5lx ���#qWx%��w�~��z����<E�V�o]Y� �o�R�e��� X+��S�rH��"�&�P� }.Ё���s�@��8�7�	�$\���!;Lda8^d�z�*�o7\�����XA��q^O$�x.�e��Sw�{��ȰSY�
�K�r��t>��	��y�G)�|J������}��El�j�(�jeH=Y��W|G�Pq\[92�a"
�2���f~Bہ�m�8L��f
�_:��]�]�^PdJZ h<�~oD@=<(�`1Ю������ ��g��믿�F�����_��l��5��e��a���Y'�Rմ�l�Ub�V�v�>�����NG�m<^�S-k+M�9�ܽx���������j8��}_�z-�����A�.6��Ȕ"EH���ku!;�!.W0b��p\��6������e�iM��y����������=a_`�����OW6ę�����	Y�� �G!8�f�Lk�^��o�N��Y���=�u�U����Ѩy�z����?on�jx��l)�oH����
�,�"+k������!.���`�q�^�~K����Y�Ճ?������ap)�����_0�Т0���?����ڔ�>g��ɳ��n�AQE!�P�7G
Yǘ׋�.�S-�&�\��8X���QT���������%ek�8x���ҺR�������N��z�P�T�h=?�h�n
�*r�7�2���5h/�%�A���J�=����(h���C�����iM��hH��7�(\y�+%l�F,6�o0P��̀^��t�Ee�!����K]2����z]iv��qD��>:�)3K_jcG��V���y�.�D	� zpRݽ��������@2���9|<l���B��[��wH��( l<�'�[N7C|����$��� Dbx�,!;��(аĜTu�<7����36±���zb^$���P!F\�8Z3�%q�X#����￷,�I��º�5����p�A�p���deA"m�x.߅���24H)��kol&���b�G(DxsE�%��&�[���f��H��v���d�;VqwY����L)���濱��C
3���d�Y�0�-B�)�V���A��"Ja�`~�i�m���D+�P����\�`������D�3o�TR�6��������]ie�Ԧ�����3�2��Lw�S�?��}�+j���yA�����r���w�$xq~�e�=��cdl7n|$.���l z�IM��'
��1.����)Jx;�-�~���I�op�ʄ��Y�1�y��Ν{�dz|����l��.h^�F�v	��C��m���P������&yZ6�!�`�ra%wvs�*A�6MM�šjy��A�N�,�HͫŦ��t�ԅ���"��L�ϷPr	�H�r�f���g���Vn	���x�Pf�̗����IN�~��@�ZS��b��t!@CkS�j���<S���T�����s�Y�R�G�^�Ն�On5��!��~!ZC�ñ�v�Z�eF�������L9$��4�e8�wV}4��j(6$��o�`E�9�32q��z���z������V��� 3$�n�nѤA�p ���G#���M��$L'E2����=�������!N|��Ñ�4�$I�5���PJ�)W�Lo��Rb��X���t�1=yV�Z�Eэز�'^�(�"��<�j�����u��W���q�G����!B���ϡ%B�1�i|���Z��ٽ�����U��a;�<�$JeGCu5�:6Li��) �1�6&亁Gv���*�����}|m�]B�P+z��C�F��}��V�׶$�f����������rc�`Qr�ƽ.���I�C+)-S@u6۟��KJ�[Z�g�%U�bs��̧����?9��on�3@(bC�����i�Z���1$��!�9�o?�G�+;k~�Y���������ɮ�EP
�:ǿ5eQ�
 6(���ե��#fZ� {?��=J�.Ȭ��k�\�7JM��th���Eyi����)}Ͷ�4WDˍ�M�Y\'I
��:�ho�/>�ؼ��7?r΋�w�Ҝ��;֌�=M:6�	�Ý��I:�(ډ��6Eˈ�_��I��=���SUP��o#�jkG��\Uk�4F���movP��B��IW&���`���,���хV8t��D�������Y�\xų�T8ui��>.x��+���E�+(���MU����5A��c���q:Ҏ8p^W�d#)n���N{����Y�xDbX��P'a6�liCG�Mok�дYKYY��j4�2�\:�zG������ж�=-� ���]Y&qvP�9ER��PP��53�E����jG���s1S]�8#�i�Z�>|���8G5n�z�vK|�7��"�dn�ܑ)c!�Az�[����e�������Q��0{E&���b��P�q�Q(��%9|��@��a�AZx���~�����T����'t��Ȭ$�eYT��ĒS���g��*��Ey���|$^�P��Zm�OU�P���e�����VzI9����.&���F���+&^E	��z67�/-4A]ݯա�z��M�P�-	��RZ��[��^��Ȉ;�+ʑe����[X�o��"J�M[���ˢ��vU���	5���5�Qe ���P�c�M�����kɭW���tC��5ue%)J�']k1߰~�e���-YX[^�����a��$Gv�}��2]� t�{oϙ!G�(�ZQ
���x����n�~�wM�"V\���D��x`0�����n�+��{Ϲ'3���hbШ�ʼ����ל��]�2��`��N1�h,Jc�'�j4В�;�rS]��ފ[!�Z����#6R��\��5�?gn�u�eiD����)�\L)���B(�]�tl��.{��H�WJ5J%!!P%�<�����=��T�����,u5�|N���`8LYm���ࠊ�+K���
j?�.�C��^� ��Y�nF�e4� �Ti?Z��
T�Kߙ�a�"�=���Se�=�༠8�p+���/����U?.��jY�nT��,���ځk4<έS�wG*|ߘ��,pKT�~�/�v�Qp�1��=L���J`J��x�$��ƿX��{���c��5�����4[py᠋�k�]g")���J������wW��x H�HpY9U�����c!	��q,Vg���+�v�ܲ�"���MI�\��o	v�rQTn���:�<�FӨY�-�(��0��Y7���H{�D֜V�ӧN��jA��������.�H�Y"�t9!�.�,`����4p04ʚ�	u:7�OiyMӂ6w�BT��R�cE��EB����u�F���OՋ .�VRʅ3붃��Zr��HVS���䖇D�d�t�y �'�)�{�)������?l�|��L�����\*�ͬ��3M7���У��V��z�����:r��=j7�.y�K�>��ۅ����b\�n���'�+�w9FX��Y��$��I����y> �I� ���ì[�~_d�D�#�T��rO�g���f�����Uv�y���|�:63���[8��A�� ��e� ^-M�j?ƅݵYc!h-,�F���ՙC�c�t���wB,)(\�5�m�Fk�i���Q�����ՖkyH�y�QY�q%�f��h�0:����˿�Jr�j#�N'$�>�2���a��@��ǎ՚�(Pb�D���9�|%��H�\
knn{��������ߗ֓2�%)۵��(�oۖ�nT�%�# ��D�ߑRT�\��\{�0�H��Ř�e��8[B�ئ�z�C�=�I��6cIl����zB���ۻw��� ��U��]w!\	T7J����/_�d�d�J�{��)��Jp(�����ښG��U'��,f\2H�[FO��c�����>%؊�E�RH`3��&���0�-�.��=;�h����Ѹ�����i�"q%��[2��4Z'��{�iC7Ұ6�̧	�.�d��x���[����5bD/91EÔj�����|>u+]u��D�$�ė����l�*���W_�{��J��\)c�u�?Z������d���3ƺ@: �e����rEd��4�a���ӟ�y�`��ԗ._ҽw˦����"�0�O��L�L�{y[������C��I��o�� �#��<Ux��s��<O#my^��_�QkƓeEs���FB8op��w�4*�췄�`sI9��EC�I��&$ �+��*�R�X#e+�Ax����T)�'��^�����1�h�����HװG9q3�;���S��W_���GF��ay�z�8S�*6D2}�����q�q��676@I��b�2t��W��a�<����g�n�M޸~SM޶�=�[[�ݻv���ǎY��:���7�Sա�.�|��n6���2t3yik�Z��%�
�ł������^���W�AS%c�/E��������1�g\���l��yEA�5V������#�d�:���D��+��%G�;����G��s�{�<�U���x�\��@9@� w<�>�h�7��|��.]���r��;!���Q�Th�r\ۃ���f~���p��w�^�2�F	_�gm��H�:/��O�>)c�Vpb2߂r�ߣ��?��<�����믽.%�,@ȝp��0�j.Z�����¹�;�C��͆��C����L	�g��%:`��5DU��xX�� g6�	���g2�d�Ц��\ߞ�T�m�d���,^]�8Y~s�#4�\&F���A|	L��C�V(#���dûȜm�8���w��2�g��6�%���~�J0n��?��ͯUs�AH�3`��lTl�n� ���f��7�J���F�f�aN�'�"��w'7q��j��?�۷o�~�Y`��Z�e��]��z�ڵ��������Ԅ���%ȳC,�=�9��~>��)�N��t���fd
:�P:�����?����>L�:�:�4Kb�V���ޕ�ź ����ˋ�&����2N��1���K�AP��=��'���V�)5��z+"�v۩�%���6��������p*�hy\�
MA��]J/J�Ϲ�oM)Lc�=��S$���z�Q_�����w�|9�]4�\BY��_z ~e��\���H�Y&;��'MhY�/�6����q�2�rC	+ZU�/}�m��mAF�fZ�[�����8p0���<c���;x-�_Ob�5�K��K�aa�a�{�NJ������fb���kf��L�������3�~i>���i��ZUNj$�g5%7R�u����TK8a5�O��֭�a9* Pu>j��������F�x�fb|���Jwm��e�˲�UKjo�XS�ןǵؔ+k �`��xm����;�,2A�:~~m}U.*{�=��Κ�沯���[��ըL(Gc��k����6��r�3���\2<?�2��gϲ�}�WS�6�}R�
án�^���9?����S��z�C�8��_�v�
>P��D�@Pэ}����G�wĐ���ca�;��|���b����F��A�a�=�h9�Bg���Yz'�_z�$~7F,o��j���D!ҷ��S�n	R#�ȢW�T�?��(^�h5�w\��j�ʼ��x2�I}�WK�D;+g�E�w\��q�/ñ�|l�z�hƛ[	ϵ�\g�&;��t��W^~ET.�Wae/]��z?���u�.�����lf�҈'���.�<_6��t d�5m��0Y�m���kNe���qT����ơ��"�3���f6��kk�F��\�)u(�X�$c��Db�l��$%l�V:�ٍ�bMB�w9zX,�9�ס�<'k��d��2��,��������~�:�<�:��$��ΔVP.����p�����ů�F�	�#u��k77�M�gV^�6����B�`����s�>�5^~���	0W���X�O>�L�/UUү�K^�O( <����ރQ@�~�M�ݍ�MF@|jL�h�u�)?qN��&��r�g�|x�����^׺"�����%������5|���&
�;�R􌖢��W_������:��|bJ��2�H�|e	a�a�[����y'��%گtN����oWɺ���y��]JPP3��/W�23�I<��7��5L4G���D{�}�p	Z<@$��:�˟��\X6��&YP6xM�^�f#D ��	���}Po�]oܸ�<^��2�Ⓟ�N6��LI
X�	Zآ����e]�_\��_�z����50�08$Ǐ�T�2���~)����Dp(G�E�������}���{{�X���SK��x��S,.�x�?܌n�	���X�{�T0� ���O4aTS$5��&?`m���~��?�)��1 � \/��U��8��gbL�)��G�0�8y,
������&��"�����f��X<��u8`��O��n�����D{�Ν;��7Ռb��ݻ���Fb	�,]�P+�۲D�-8�9��$��H��3c�G�)C�Л�������y?q���ӧ���xOtR�����?���+l$�N+�F����)(�y4:$w�/>�[���?�J񞔵2�YCn>�_;���"�ج%�-���SJ��2�g�R�b�� �m*��R�J�������I�Gc�R���'HDv�B6jaᑴI�jq7?����9/��vI�3�>Y�ۮ�אU���!9�'O��G7�$���D�wgF܏�>D�3��Ӳz�MB+����	S3���pA�uv�\ط���頜�L|:�%Ҝ�k��߽g�f%q_I*��P��?��?���oD7|�j��G���?�sm�&X���]bJ�!�C9��kذr�׶pf�Kw�M����	@��\R]cYE��q��->�	��o�.���/�3ٸ C�YIoϞ�Q���Çe�&ĕ5�$&�+�^�}�����}��A1����E�?k���I�Pt-�<����ĵd�!
aB�h�dkG�_�Y�~/�`�2� ���Q�����㺋$#��'��x�=�J��)9,{ڝ�hq6
w7>Ͼx6,9�nu��R����ԟ��x���Sw߾�N�
�#��,1�Q�64��F�1�A��� rH.ɒ�ؚ��:ұ�j-<z$�jnA;��������XZ�'xC-y�Y;���!/mJ_OԵh>Dq�>��3����(�{���5W�֪����5�pu�"f&�m��V�4㺰���i�QsR�%�,���pG�^y-:rBY]b͙���H�>�VBj�ES�52(kH�1'�С��9��&h��p�0X*'r��s�}��K �Nc��4�>>׸g��P��L��M�{ơd"���>z�{b�9J�� �}��	�J��/>{*mi↾����~�{ql����M�a̘��[��Q��ޒj��GR��FR�U���R"L� �&��p�n�e�5����#�����!�<udOh:�Ī(��neR.�J�B�4�}����C7XED�+���ZYyF-Ie�g�q$8��D`0�ׄa<r����q��m���6ۖ�Tu���O�St:���V�h���*eϽ[O�Ƀ�x����y�"њhtL=�s0$a�)v�j�*�����u#S�I���'%����H�-�I����-~�<��W���ynɝ��[֮����Q�I����f��2�j�R���z�sg\���E�m.z,��:�B�9�Pgq�^�+�-��Ǐb�����OnQܔ���J��!#3�j04ks���p/
�>���e����1J��%\��e ���]d�{ᦒ1e�(�)�$p�H��"%5�&Z��(��a\��P\��Dn7�pߏ��g�����F,����	K6�/C�e��6�������D�����
IP�|ᄗ�pu.�
��M�� �w�J���D���X���*ip=�jڔ7����\��[�`�\�v��wzNB#�5����?A�R� <}�$�{�}���*;vX�aH@����l3§�坙����C��ǎ��1$A��:yFI��o2-��mL&¶kǌ�;�8�����W�/e7���d	�
��7�B�|�y�n�)��աR6�[������3fC�﵍�����G���SV��}Ϟ9��r�}�P@I���geۅ�Z��V��,��֛��m�~��8�,-n�?y: 
X4�b`�CԾ�(�hy�W�gV���(��*r�p���ʹ��V����������~�[;&�Z�P��,oS!��_|����0el�6��7���sC��p�<�YB�1���o���L�>=>��nY}^�9�O�.���ϖ�w3�T.���s�S�܇�QQ��De5.��aI0��@������k=�V:	�o��>��3D|>��:|້{�"�+Q����FJ�wc<��ά*���mCZ�����A��3HF�2#�PzR:1x��~٢�5���C�=z���0�2W�{��Pl��Ǐ����b`�9�
�m����i;��({SO����k��;f� �	��w��z=S�g<,���Tg^>UUp����=�Ps}G:���׭�d��sa���J�Ɣ�$P��1��pd�U�Q�Z�n(ciBc���T�Z��븉s�:L���-]TYBf�X]oU+�w,w��qB5�>����7�vBu�u���)?u�h%����N��p�?�=�"z���tT�%�F�O���f� $,[�#�}�3^|�(
MSV�{9�o_�
2�������+�4�׺�Kj�\��^�A�3�Ƌ��8yR�xq��@�%�!ѝxX����`�[�(zQgN����AYB<�Q*I>�k�"{�dQD�0�[�wF���2/���� ������`He��dX�W��a~nW�r���t�=.��/�v9����"��ǁ��.&q�*��x�m"��$TR)I�5�J2�qG��p������_��sc������q�)W�`t.�A#��5XX�!Ŋ��| 9����_SD�5�?�Jv�P�j��L\�ڃ�rq��Q���L�%�D��B��'J�M1�N���P�mm�is��֩��DѵZwj�����r�}��gp�YːT^��$�r1$EM�6�U�a-�7�y��1���Ri��o��_����@���;E*7��RVu>�e{�kL�P��oݺ>����(ƍ�rV�%�v���F�2^uVL �hzH��ħъ-=c�����+돥��t��AhXH��Z��ܱmFmk i���wZX�����LY�/u�1"�����E11RF�4?fi���ƞ( N1��5w?�����i��1�P����iie�.��Z��h��
+J�1�^Mx�Ȓ5�&<y�dIzsݨuP"��Μ>������4�&*�]�<��̏��S�tn�B��iF��^��1�}��u~~{��{�'��-t��́z���K�T$�<=�e���w��D�_�ڄ96�j3�-�����X]6��pbJ�/��Z��\8z����Jt���LNv�m��-��r���x����?]��c=��dV� ��o"z������X_#��SB����fhD���<�����=kY��_փa=y�t)�֭�026�q�B��.����P��bAD+Bl���^Q��A��Y�8���4��,8Qz��zp`�����Zı�Dhd\jbH\^� pɋe�)�㡱����BT�ܹ7ƀ����,�� ��H����w�m�.�x�ȑC�a��& �QB�7l^���kY}����I�^�n߳�qj�kX�"(�=dL��4���B�ڕ�KJ�9���ϮS�6Y�j<�­���c7nv��ob�)�}�����O�j|.�'2Ӑ$�Ņ��a�ܲ.���KF�юn�u=_'uXi<Nj���vP�̡xG��$e��	�<ٝ��C�B�H֟3b��i��3GA���P���B��M<�W\c!��U�z;�w�1�ؾ��:r��:E/�"�g|��8�q�F����ߋ���Jr��4��؀5^��,�g���� �[���~{=@4q��FC�B;��qo��O��ӔN�[`��>k�V�f8Fu��l�����lkϬ2V̐bM.��R�A�(j`��3�d���NL���R�*X]�{ǖ'ɼ^mxc�X � �q�)��U%YB�K�je��2��q�[�MʭߚÅ���I��kr���
@>补�g:�DH���u,˷�dP�Cѵ%�B�x"�sȊ��Pg�ki�#�A#ADC
���׉E�|�T��û��{	@�:hr��m�ݹS�uOY�cx�$����\B1�@��[m|˦��QhX� ��I8�A�e�v����i���!���Yt�����>�J����q�=� G���>�}<t0��l��ʑa �%�L[�B|����
�y%O��?��s�+�U�慅4v)�{���A�����F���s�����L�4�����I�\nɸ*9aG�
�@�U6s`�M���ߘ!3�8�"e[�����Qyޅ�c�_B���,��Dg����}jk$zS\m��b�=l6VY���M%�����V.Q�zm�o�9�.$K�:҆H�?�x�BE�2/6�������?���r�aUy6R��"j��hi#�V����x8��31y�L���o��W�����,A�����Q�&FEȢ1�=^��2j�"��{��%F'þ�W��d���� �Eo�r�p��
l8%�^Bp�hlbc�#N���L��%\�?��� ވ������^:�rJ���7�=z(����>y���!��:�z�]Y�e75y'>�v	��S'�=3z�=�D���ǌB�����q���g����8'#�	�4U�0L�h������5%8��ߛ=Т�v�)Ƭ3��٪z��� 4����<);2xl�pJ�>��ͱ���_� ��k��rOt[
!1߾c�)/��İ�|�ݼh����&�k��ԏ�Δ7@�D�P�i��/�������J����Vd�\˼A `�	2����Ô���ғ�d��z�J��7̀�_�� �~����`m������5̲�Ѭ����p�S�7�s��Y2�u�X�g������X=����A�N���p<*>����0��%<��f>ۚ��]յͫh��YG39�߭�Zcۨ��Y3�C�g�k�*��椈�޺)�s���I�JhwF��
�4�0z%X%&`�ޏ�Ɔя?Gc<�ګ�u��c��z;z.������o/��Q�pw�&����K֓��bU�=&%��L֍Rk5?�';q<�8yZ��q�X;��F$����m3e[�o��~��<l�J!k7��U>��V�l@�g,A�}wn�_s)��ޱ��|@��K���Ɗ��'쀗K?Q�Q��Jf�s��:ކ��&yI�̅JbA�Þ2��5��ƍ�Jf�L`;��А��Y)c�U��{��w��?y�(/	D&��4YE"1t<���I.����,��[�Y�:�pE�5����"X��֥�\/�\k8pa�z�%|���$�$D�I�ǻ��#�y�+~%ˢW��Vف��c�|��w�P�(2CqS�kԱ�M�ĕm�X���E;�ٻ��V�:�pKc-r��*fl���2��MͮZ�.괵�Mes9	m%s�։ب�E-�;
�eb�3�+��?~��f��A:Y�.��)؅��Z��X�w-���Pa�s���	�d�q�GEE5b[�&��]s�%�����f��{�ғ� ��pC�i�Vzz�2��x���Y\t�|�M����i�H���AB�]yk$��A�u��w�ltç����e�7V���ｯ���3e�6���?���C(9� �!��E[\)yh��0�R��lj�L����nRl"$[sK�p݄�������+����Y#$��������*�B�m��1�;�J�G�Ͽ�LC���� �#ku��g�k�Y[�O7�5���m���s���V)��Y�JI�"��
Y'	q��2�ʱ�k���|�6�xa�9A�F��1�x�4���ּa=���`�8��.X=��YO��x!S|����s�7�]B�:oʮ#���� �@cNN[�:��il:B�s��u�D������֎xvaa1��qs�չ��N�>k��>�w��q5�#�X�_�F�|�UZ��捛*�x-��h��O��������^U�{�j���0*by��J������|���D����_ͤy����zF�R���u8<�˗�H �������O�w�JSe8�j�!	(��A2���K�9x���<_]��-e�����*��%W}��䛩��=��H��BIB�$SK�?V����G^�'����~�#	��dW<�݉n�K1S�h
���H�ìng[Q^(��v�L���e~�0���S�&D&z��RW�.~��~��!�a&FZ3���%II.��k��cj$v��e9���Y����(�e�-�t����f��Dm�P�hp���9�
!h���&�\��|!C�<Ω����	j�àx�r� .d�o�4�ƠW־5Q2����%���q��i�����<}�)�MC\�mS��$]�7YV�������0��M	*��~��9R��d���jD�����G�E��.�����Q�hvf{�AO�xR��(��� ~�f{r�&l&M�s�}?;����]ZL�������7R�ĳ�4;�L#�A�s���=%��%�%�lM֣��r���͔=�:;�0��o�<���,�D��n:=�Q"jmu#M���}��z�+U�=s�jj�!e��v[�wjbJpd�QF�qꏶ\�+,v�F�ڤ��#��@E���H'�EO�r0���m]ss�Z�&Ϯ�$a�����[��Q��wFUAC
4R:�5����I'>ō�����W�y[6E��i�Uu�2KD9`^��Yt��u���O�g�}V�U���F��>ޮ��pױ��){�@�r����[�0�Be�	t��������Ȍ�(�Fv�G��A�̐fL\ �f�@�\x睷����a���oJ�"�U�U�`Hm�F�qQ���Yp�({0��.%�P&ɵ���J ��{�^�"E�� Y�e�y%�7�~��F��̾�N9ʓ�?��{,��q3����5%��DW�x�ٱ���=����1,GO��/�ӳx�G����kYUL:6O�X���@s��4�1
F�2Ʉ��m$��=�b_=�݄ɷÍ'�����4��#�9=��	�����燵v���ű�� ��;F�R��,��+αaⷷA�W�^�(_�
�PÑz
�/<�B�$`��d��Ҽ������(
>0(��.kun�Yo%�ԕyqȈ��tF.���;6٠pU[��&�*�KY/~����g�T�
տ��T�0�b@ppXOl�Wf��69AGUf�0f_y^�"�-qrB�K�ivR�^�$!K�F|���j)$�N2���މ�k"k�`F��f!ln��qCn�pX��&u��J<���Է��v�[�2S��&�����P�V��eE�*����N�Ο2�@,��M��*_gk�H$�Y�g�E(@s�z������X��O8�L�et��ϖh��Z]z�,+/ڪ��Oh�_���Rj6'�!r���Z�������~pb�y���A��?��ro��$�|4��Qq=���&sJ ��7�3嶅���+�W�2x%Y|)N��^~��]��%^���bύ�85#ey�y�`ّQ�<sF˒��x�r�X�ܑ˚ר룖�PY�����{�a� ��A�F�A�-�ڇ���M3�IIL��Uyr�YKŋF�����e�b�+�hl0n8�ˇn$�ѕT?6�SqDa�_ȟ�޸����t��t�}����vS;PF�;%�V"�[ӆ0N�Ɛ�	he���K�{���\xJ�D�d���d֣˼�<(��V$X�D!E��ۢ�|���wuZ�|��+ѝ���1S�f[ �����kH;�"^��X���x��3�y������ѪO�n��_�ϫ�;$��{6�F�y�ηf8�lx)�攸XC�Z�]#R�����.�4�T��g�)�gO�v���LV�<���]JN�-�k��%Q���0��W_yEg��7Eü'�j���r\�Y��gNK�%���8?"r�J��Q��s:w��Cj�T�{��T���6c/�5�nn��6r��4��)>4�#���Ƚ+r��8qܥ�&�y)[x���FTyI�^ƪ�V��=J?C��{�ZֆeQ_����C^�rma"�JC�a^�Tw�K��$���S�z��%�r%�Hx�;wN�ȏ>�HpQ�g����r���}R&"�M!����GTas�і�F3�A���N�Z�Jp��56Ԡ���l�It�I���߾c��O ����S��0��QцG,̽g)i��@�F�?�F�7�co�S���p~d�Q��ɇϴ.��ė��J��0�Y���y������A�_��a�䎸�Gi�ol��_�t�l�ڰU�G(�#�A�C����O�ݷ�B'���
M�E1Wg�(;�ī��:Cd�j�!�݈�ZG'����)aH���϶�"n�Q�^4����S�	����f�94�Ol��2�q3J�0t�ɓ���֪�����&�Ю�Lyf�E<�U��3��V^�'s� )K�^���XDۉ�Ψ�F�^۹�=d��<���Un�$�_�Y$A@vK��3��x��ap�db�<m�"\H�c��'�3[]�X>��v�X�m�{��� G��:��C#jK���4M-�P���i��eec�<�Cud�5T������2�f���y� ��&74ML�bY��MAR)KM�ǃ2�Mn�a���*}��Ph�g1�!`RX�B�"�ܗπ9\B��tej����i3�
����+1��'Z%�	��GO�7T�kE�5#����߇˗FQ�����v���2����_��))��I��D�@7n7�x��c���5k����ǎ�{k弣GN)�����S���c���ְ�M��0��@��wg��fG7�wѫA�߾u����hZO�p�QN(]s�G�4��H�܎J��4�\�ج�H"��'�O��`�����;��P����l5ye�%0�+u��lȟS��޲*Ҩp-���777��r��ȁѩb�F��4����vd��`��[u-��iD_֗M��,6��=,ʱcG��Ɗ�w�+kZ�MƵ�?�E7���G�p�� 'S�ZD$�7�#���C��Q��i>΋�/J!l�{�m�S�����K���7?�/^
7o�$�ȑ}a:
̳�5	�J��	7���K� �dt'~Ft9Mk������;�X7�g�77��1=|p/Z�ը�ۚ��o9ޛ�C!74.��5��i��#�~�t!|�ŧZ�#��F���sm�fS]c7�t��d#z{��߲�B�}��G���Tx,g��"s�9jJ��ɟ�~Tzp��h�W�dѻX� �\ߌ��p���s��n�u:��O§�~.V=��j�%x�4�A��[?0z p�`~��G�~䬁c�#V����'������$��~c�Y��u��7z��+1����Ouf!�@�{�F�d(� �j�m�� � ���U5-F�k�r9I9�܀��'�S�MH�!$l��>x� �k߫jS������Ď	�F1J��X'�	�%�I�g�� �3�KKD�Q��\�MAƦ�ܹ+?~\��l0�
������?~�&t�k�=�C�Eg�.��fq�fh&��k��H���]d�x�f���ݸ	Y!ט���\8w�lx=ntgjB�(�4%�2G$���Z����*G�;@���2�p>��{@TI4;�2ڗ��ltQ�X�n��DC���7^���o� �L�I�䄕:�N=s���^�X����2�1�L�V[]q�����ޱ���Ϟ:'����y "eh�홋����C��[��sٻo���]x��76�����>쏱is��(�1�ύW�� ��")�8��V�Y)	pWovn޸���K/ݏ!�c�7R�� ��~?y{�/��MҔ����!kMGՓ���&�6H8���\5�}��mZ���+H7�v��Sf�QxC�a��=�L����HT �Q���(2B-\q��r#���i6���Ki&&Q��+��,L��u������e)Գ	[�fb �G\HkLM��9�	�R�� ��_~M`�3>s�\9���/����X�g/s���e61F��`,��F��@<S��h��<�����_w��+�53E��|�5�S�Aw�U�bok�T&� �n*���ڻ�{������3�����z�/��EeOO�ʥ���[o��gOu�L
���'���������dY�,Fy��A��=�O��WM��v��p5���������QL��wn����1(�K �.~}Q�g����T���g��^�inn�0��a���ƭ;�'��֥^�ϰ�w������������{����ﰞM�۲>�.^��߳�FO�����c�.'��>"�k�ֆ�.���a��rY!�����E��NTN���p���� d���7X+rX����{;z�X8}�*XP,�M���c^�x'r(�w�����o�Yu�l�>�=�ׂ�ܕ�W��}.�����
X��;����Q��c�p�xV���.yr�(��R���6NY��ye/���|���B7��0�F58��U�TB��D{��y;A
�x)j��T���#w��>��J�Ɖȡ�t�	��#tpm�Y������![I���ƢJgh�+��\xI)�m7�?h%���T;^�����TH�#m��RpG�;㡼wA��3Y�x=r$�A4)�|���!��,��X:<(������F�G����`�U��<�4j喬{65e�uF0Q��v�Ϻ�|2G��(�������_>|�XܿU+�4�������໣�C
z��z����a�-�y�䓏��6Ä�47������j�!����|e#h������_F��y�f��$�qOVf�@C�(����;Las�V"�(qF	������x�E����� �܎9�I;%��`��BK��o��r�:��Z�\S��ϠL�x�<J�j+��0� ]�(d�sӉ��W��(�po��r�V7YS�3(o�D������j���ٰ��>{�ck�	&o���?~��1�)8l"PB~G�i1n�j��8�|@�֒���$ì�(>}�8�q�'��kăݨaЃ)��1�r�H��K����5Z����w�3���HM��
�|�m%�RAZ�i�Qv����C�x�t9Lܾ�6�&�'�j�w|���A!�X[+k�S�b"����`��)�v����Q��]^ֳ�J p����l%4 �c'��L�u�^�~������[���37��N��bFX���[��s�aXZݔ#~���va��Z�67/���>��W�S	�?&1��w%܏�C�rh���������7�|=LL�����39���ܨ(�G��I��m�P!�I:�Kqm:�=�ꈹ���? ��rk6,�C�f��2��{������( ;{������*�B.G��Ĝ!I��hOIeB�GQ�<�!��t��������߫c��1�T�rp��x>�Iqza��J����*�ʬ(%�b�j�ޞ�ቲ�}�QP��v�e'�����,�Q��	���B�@a
�'��|#���i0g�,�^܋f����R��Vok4�񶎦�����'���;p�qOD��Н�%��˸��r���׼�ѣ��5~g���G��#1�ƃ��{��1Ձ[��;�PV�"w����l������;jV�?t��{!$|4N����0H�,-�*�u��	�����o�H��$�p���X����ǃ{XҊ`��5�
ao����i*!ѵ+
��w���j�U6	g��C�ë�� |����Ջ. Q<��m�;�=�<�R8|�T�\�	�:���6� ���� �˝׈�x��_yE�.�3�l���'���SN�WՃ����>n�F�4�`$�%Hdn~�j�KgN[�u�y�6�#��mXv�ݼ�~�ih"Yl	N�x���r�ɜ?��)�w�otm���t��w�,]y�=G���p���j��F(��s�AW�^�6P�{WcL���]o���KU��l3�Fmd(���rw��(���iY�~}ls�zEe��=Ԏ����D�5̓�N��=aְ�7ާF������i�y\�����7�x����{���m0Z�u��vt����V/ӳ�x�^J��)ixo�Å��#V���0C�Ó�PGa�p1�`��UF���C�Y[:��}�6@�L����9r��ֈ��yf��Xr$������Xʛ��x{���KhJ�5gѰ�hQ9���|��?��vT�|�M�=lW<�3B�1�m+������R�M��U6Ʃ�>L�WVO��̢m�I�M@�K��� �ʰ�����8�M�Z�y'�-��5�[k��;�X[���)2��-��l5�8�����|�Mߜ5�^|v<�\����&oS=q��,>QV�}�w�H=���苫Z3/�O/Y!��P���
k�Z^�	Y8m�0"Έ�K�cY���T��V!W�L-|�P݊�nQ֋�i��,MHp�v��0a��n�	0���H5C8�Q�V��QnaA�����gg���U�1�R\/n�a�iM��>4�1�����O��m�+��)�p�V�3,*CC�A;���	��!��)�@)l��F��$�f�!��u+��̯%�&d�}��H�͢V�:����T7a��U�� 
�i��^�����������$��.�R���)�x @QP�A0(���<,;/j�Mք�E���r�0��}��W<bd����S�v�����˘D�������&��އ��h� :��f	�����Ž9����{���yO�>y���f٫�-1�B��ő�R@���$J�_��_(Yf�������Hz��%��@���e�}������r�1���w�e����0	T�}�����]%��S��7n�>�Rb�g|P�a�:�
b��GJo�#D�~�+ԏ��J�+Ӓ5��_����>��W_��a��&fiڥQ����j�8��tA�e2�Ȭ]
���jg�M��>��0u@�6�+~�o��o�>���%��6��9�B*�5��t���i�2ٲ��^������5�kVuf]@6�!+���,�Rz.�hV�/�Tw!]�o�4�k��_I�a�7?RBQ�P:�}F0`Ⱦ�ϱ�SO88ƕ	����P�W�zn�i���S�����l_�J^a}�=���=FN�C�q>.�=c�	e���T���eTXh�x��rp���Ξ��5�#H�ݸy3|��'f��PsQ�	���¯�+�^^�w0�Y�"��rʍ�i(�7�����!E�^a�Y{7kQ�����hŷ�z�bjou�z�xp�Yˢ2�M�4��l���0גCG�ss�\q �b��7,�luj�æ���P�H+w["�<q͙j6�!BqV��L-���
ֵ�BꧡoSj4,���`c)
�`�ޮȡ�X�Q��YP�4K�JBx��P.��5('^Z9¦M��c�O�yKd�&����3�ڧY��ƈ�z>'0��b��!p�v�m �)=/V�-��VH>�Ar�a|�n�A�԰1He0]�^�]wU��UJ�ɒyo�!5���6�_5Z�u�栍�.+��c����}���b�uo� �;�31|ց���S��u��y��A�ێn)�3۪��S��FgZC��d�y�_~>x���%l������5k?��ܱa9���U�GB���@;s����3ゎp'�`;�8�2�vq��4^t	�
��� ��6&��D��l2m~�n��8�l8��h�F�d�,�T߄�4N%�Bm����2#ng��E��?,;Z`��B+59��FR�c=N,���{��wL��{�.�6��r�ˏ�-�p���u��+�O���o$��hnI�)�2k�2�y�d%.�k�kJ�Bv�G[PE��u��%F��ZX����t*�R�un��gW�x4L�'�d����p's� <t���K�������h���:�����,v5�J�U���qX��q��r=)�0$�ŦX�Ŭ�(��gZ%u�.�����̳����Z΃���G�ªNǒ��&#�'�\�
�ڳ�����g�QF|��F���š���_pC	����<~xY%�N{M��K���j�Fc�H��\M�j��V?1Zc���=���*��*~<�=����%[e��'ʚ�P˨i}ܧQn<�:����뤜���S�J��SAI�_�%�����!/]?×�q%�@�1��i*�	�;�6���ע�{�����5��60���+�Hv�KG�Z�y5��y�\��y�|�]x�1-�iJ�fc�B0/�8�T�<\q���*�j�	,Kßf9�'�x�qyR>��=��YpB{�$w��~5�4���2K
t �	�=}�x9BT
eVŚ%~�������~��2!k]�y�f�ޘ`fT��Z��4�-i�z�B?]�ff�i>ó�Xl<�85<J�������c���}pfl��F�p�8L>�����h�7�u��r���`�%5!�����.���*q#@qɉ�A��=��ío:�`��X��9]�b[�%�SI)s^�tS	�3ʪ����p�}&�<,L���
(��%KYآ<duaq���=z"J�¹۬�ۚ/
W�Zd��|�����Ou8����z)��F�`W3�2�p;J��ߔ"$�u��a�'+͵��wjY�w�Z{����[[k���,�ݕu�ʪ����FB湰�j��/�$(k9�5G���8�,�Y+cN\L���o~=[|VZ/��n�xY���4���L�V��r#��<Ӡ�W��~M'��P��b4����E(A��Â��=�f��Kcr��S�g�
���#̬�Wn�%���B<V{8��\_���Ts��R�1����6�,��H��K�|�k׮[WK�����w����NP(>���l���z��bj���5��nt�`���{����VJFS�X���7�c[.�x��S�<ock�w����40��0&�O��	. �L=IK-/��*��=��.�=M�M�H ���c��*��3�F40���l'o�,������F"��ux������n;��-�'Ό̯9��c�	���p_�ݽ�s�p<��=�ooTp�D��R:k���R�g����������<�%�cF�llq�DK�}����^��y8A#�γq��Kª�ѝ���a3�%O�<u��FF2�tV����S=\@��GM%IBOf��˝��W;��y�O7j�k�Hqw��O���) �\�f��K߄��U���A��xϊ̼dgF����C��E�m�c,i���,�ŬA�	���x�eOV�z�9TB�%�R�Z�Wy'��#�F�n/W6$-W�����F���`�E�iz���7j��~����ˋqF)�FP����E����4׼���a��$��ci�*�=>�Kq���f�^{�5Y��`�Wbk�hUl7�_!8ʯ�jYW����!��Zc��E���:z��?���9W���L�S���s�9�Oc����\f�J<��&؜C�����ap&);�XS�i	�	y����o�5��WZY0#�����0��H	�kdI^k=�j���xEY��e������R����m���C�]�z�"�b�dn�V��\1�|2���zh0�ܨtʰB���2�Y�4�]�γ�f���B��P�Y�;h���H�
K�	�c�b�\<Y��F��v��2���	�DMlCٍ�H����y��X��O?!�4�R�Z��1��&z��!�H	A�h������e�2���aA�|���;���o��~x��t��!r�u�#?,��YrЩ�,�Y�3�\a�!��0�9 +#u��7�Bi=9>��==�v�е���X.wG#{(/�T!���ae?|��?��?*��,���(F����%C�P`��V�qcҹ"wS�0ͪ�"��,��N*;WT��Št�-�Ѭ)Ԣ���^�|������,��`vqck�{l6Nᡬ�Y�Ia-bP����"�[Z���s�Ψ^ǋ^l6�C.jM_TT)5v¸�gS9x/�t6>r8x-ۓ���{�Bk��5U?�3"�+R�T��io,���l����sr�ē\��D�>���;�%��S�c'$�x!������{O
�!�� �$������)�ҳ�<?���������s�����b��Gb�"���9�ܷq�+C����wS�_�v`+�l\.�NE;u�])b��'��T����K.�����)D"�,�Hq�'Y�,Qk���}�;οt.�4�?$��04�䢳�`��ۓ�nx<�Ȱ��u�m�^J��������8�B)��k4������`�݈����2Ao�ʼ���:J��I7%�����d�����&��4�mJ|�U��9�,iT2^4<��t�J��~�*G�f��5�|��E�JXE{y]3ǂ��q���z�s
x���ꗇ����0�B�c35��U��*�E��jUn�Z�tK�bԝ	V˅�V��ܠ�x���Z�y[��q����?g���@��(FB�h��V����%��О��Q�)��Ǣ�m%��O���t����ɓ'�y��W��D��|Tl��V4�u�J��<�����l�
u��Ec������G!cR&�۬e��5:�Y��f'9C����۱���o�.�VF�V���c�ݻ�H�<|1G����5X�+W�-�CGV��斅�'غ�.n}-1�N���-q���'klY/�Ļ����d[B`�ČAgT�o���?dZ�P-��C�C�mS.\`��hk�6�n��~��ji��b^���Z��u�B��]�������~2z�pP���0h^b_0�h}�Ei8μ���!5��"� 5ʤ\�v�j���8���Y=�l�P3^�Z�!�5s؄�K( ���,�1��e�F���Ut -1���6��5O��2�-F�f����\K��_��z�������E+�����3ə������7�����T�&��,%!�t�Lb����)9j��aڗ,)k�m6�� ζ<W�O�co������M{E	Bx�8�_@�;wnˊ�>i�]*>��+i�j𖘑	4��`��LIeֺm�}�8�ѐ9�~U�����[U]��Ή�V��db�j���؊���8�_�$��vj�$�Xa��v�Rc��ݢ���A|NI�����;q����f��e"%�Q�Nq�B��6kPn���x�j��r�qO����i(�y?4�O��)��	��bA�JV��|'h9B�lq�Ŵ�T�eӈ��]��*���^��ł@�ϡ"3���e���"��j�MQ��,_�>����5+����o^�-����"l��뀡J	�q�u+���ͳ�>� ���<D�?��F�pFO/K�A�l�`�	e��SC�|�V%��"<}�?�pJ�d��7b|rAT�W��L���-�ǚ�J3������*єX(�y�Vg��@�	X�[c���=.1�n�aY�Z��^��Ƣk�6}B��)y��~�$6��:B��=���a󺣻�حC���B�����P4�-3+��e�.>/5��G�k<`>G�L.@z�8�,%�n`�>R7���hx��<�B��0K��N׳$�%�8b�L�:|���4mr��J�僴���<�M�9�kDR�����@��Q��H��@Z,�͛��#�5N�:t4�|Rɦ+�.+ׅF�pa�`a�������J�YM����-�7�Π�6m�"�4���g\6�xI���*�+�eK��ʷW­�7�9��������T�3E�#�{�Z��0��豣��˗�-�7.��0|EnPd�7�W���L3�|��G�?4\A��!6��-k���_o�t:��hm��t�J�(�fad��h�M�8#�r�fC-t�KVC�V0���L+���q�e��?�X��Hk� ��.�ܯ�}��:x(ދ�j�ݻO�⍸����$�a*y�U������DSw��#��[�z��b+R�PN,4�#�6R�QR�X������tWt��Vr�ʎ"�n%'�f$.T�.�a3�ݽ_v@y6�$�+���B���`��9+v���5L��<0��"e���ץ�=��ｙ:���?U|nՋ��6e,�<R��q(G~Or�~��U���6�� �D���x��Q$σG�����[�e�*Ù���\Q�Y�wv�QH#raX���y��uX�$�/{$�`J.��Z��gIƦ��g��zB��Z�By�n�.IrԚ��6;��ƿ=����^iy�1�ߌv�!c�A��KjccVP�el�(-7���&�h�Z�w��K�pOl�������D|p��q;�˴�b��KYr�)]�Z�cæ'��N��h	��<�skd�������;�&E OD�=~�3͟�CA[���=��)NiՖ�"��&ҳa)Ʋ���f�cǏ���tQ(.�����w9>.��%	/v�a-/C%M/�l��r�-��B��i�\�x�7�V�Zi��!�D�ѲJ���Ҵz�j�����!��KK�ρX�����g�S�0��c��<)T��'S5�*]˫4K<|��)P�����AU���.��a�կ~���m�:Z���Z�o�/fNr3tU��J��D�2�2�l����f�JV�Џ:�R����:�,ʟ���c[q�8
�n[*��?�T	��i�ms.j-��}K3"d����ƥ��:h¡��ڭ��fP"��zbFѬ*����&\�i����m�p�i��Z4�đ]�B�uBwz[��f�$�b6�����TV[n���C�x�G� x���A�X,+��;�)����g�����R�:���S��B���)M�$S��O��0�%�H�h�T/N��.��&�ajg��E�J-gw�0�:����L0����%Q�#)%���ɪ�ߌ���'�SX�yT�q��e�,��)�eA
�&�����ݻ��O>�}�e�(�:/�V��V��|/��~��ۿUR�V^����{����7W�]p�(��6B���d�`h�O���g�,�J�����ځ�\��ط�9v��ɰ�lY��ʅ��#)���{���7J�"���D<�A`9����p�r�� �����I�dp�A�(����I���I'p��Q'L7ϳ�|UpS��6M� ���Z����m���ڭ��M��/��t��:'�]h}���妘;���xUM!�����/D����^}�5@��W�V�7deL��j~���n����G��J0��؞�	%���k g<�d�8�.�P6�s�~+��,�D��h��H]](�ۆKD��,���f��2���l�Пկ+���A���z�!a�gZ��Q��e�[�w�44è{z#Y�T�[�r3e��;���u=x耆�s�&�'ٛ����Sd�|�UI?T�{���g�E��uѬ�x��q�b��Ϳ���ɩ��S�H�:x��4��^�Mp|��׸����E([�9��FA��E��������xg\�������cdM�(J;�{��������9f���x��U*�Gp��̈́~�A�F��IY�a^`�Q��w�їs��3�2ge�b.��fZ���7�-�~�?Fpڌ���㛵l$�#�#������ܿ�����g��9��'M�X&���l��ڥ�HC�l�M���J <�m�Q&)�vG���q����'�8�S�5|>�v;��&V�y�]��=�Gx�w�@,+��s=1F.�R������$:|ΰS�t���7�����C�s��CE��T&�ϕ^VTS0��Y��OQA8��V�����?�:~�B�B�͙̇�����qy���+_������)��+��l(� �x9��@��$��t���럩�|<q�x�bn�}�����3g���=Ԡ�1,��y��?Ao�E���kΤ���,3��������~8-����5L�'�(t��3���P��G��P�8eI�����h��ik�&.0"����� 9��M���i.Ք����r�n�8A�B%�߀�U�Zy-��MռjK,m�A-�yb%�x�oh=���4JTSA_���*Yl�&x�6B����G�(5�FCK��i����ҡ�QÆ��g^�y�+w����Lfe_�=���uS�G'5pŲM����cG��}��p��%9�8u����%��5-	�j�gW��NE�?[I!���y��DZKw�Wu�P�-u���Z��<�)x�9p@��!�
a�]�V�q�i�wU�I��=�&~��4�%T5w�EL��s���Qj'R1�D!�ʐ�iioQ���b)�=�FMhr���p5*&�d�y?%5��S��~	IL��4���G�K�4���q���>�+1y���n
��2U�ҳ��>��+kl�f�
Bu5[*O��M�IBjS!�.��_�m��ۙz��[4��X������cmg��T!L���Ͱ⺒S}�C�?Ma�����EP
#�:~�xXz��$�B\�a��H�Z�up����r��==.��i���t/z'��n+������vN��k
+��l:��l����P���>�W�5���*�K!o�-0ţBÅ*n���|�Ő���e~��IY�C1>��:3#����W�����k����<>�J}����ϣH4оg�[j��+�[��z����Z �Z���bԉ�����i���
�0匤�O}CJ/��viI٣2�1*D{%���/�f&�q�Bƃ�3@��;g<�Y��;�$zo�S;���F�]��:/�-�V
����j���K��Xa��IY�\�^}�>fPܞ={Et_��I�'L6u�3�~8^DY�gYEg���m$�``�<sȇ�M������"�̩3��n�����r���5-�,6oY������/���D�R9٢��L]4ܱ:t��t�gr=GP�%� ~���bБăs��ɂ�(���IX������)�ք�j8�%���U!@e.�p���;Q1>+�	�t/Z��QPh�����/y����!��|�4B�������[���HQ9���b�݋���Z�P���R�4�y�~כ$�ڹ7���֢\f��ZG�4Oؙ��i���2^'���\���4������;Ｃ�9���aw��(�����Q�>��ҕc�Y�)�P[n���-Qܦ�f����':[�.�]��\���@��Ň�#	��'Ҫ�y�n�V���[w�>֡����:�Ǻc�u�J(��D��lMi^�7(��	�z$���C��$^n1�-ZQ4#���P�s��_#|��������o���Ol�<��BJ���]���77���a��S�ޚ([C��/�VE�,x^���"�{���5tc`��Z`���F�B���8q����㸟M��Pf�	��]Z/p/�h��r��J��'��cc_*7������1���\~w�]��78�p����L�2J�9,���@��H���UG����<*Ij-���X7�_�L��֚$��E�6M#5Td�z #���SolBK�wC�;�gE��7��N2�y�G��ox"�Co �T4"�F{U>3r^�"<k�./�b\p��掓!u9�;4�!�M�.�yɅ���F�,���20�� �*�h�+��i������$��+H�k5/Qq�a��n�u���F%���Z�2Mtؽ[	,3/,l/��p�0���ۀ{�(7���x��6������=S>��6�/V�z���D�ǁ�dYOV	7�ȡÆ�p�u4uԡ���q���߷�z���l�|E�"k��gXo4�2tf}QVz�ZD�\-.�v�H�ls�x��[����Jg�Ex8�tH��<�[U��K78�}]Y���O�`gcB�����meG���TI�5��x�g��38��e]m�oݹ�<��Wz=�!��gq�ܹ���>�;��� ������OT`?�A$9ʳy(r&�`����(C�C��
 ���w�[&���	�JZC���5�(1�ܺG������)�J+�+�����o譨�D?�W��f�隂���5U�.Hˀ�����ҍ�Gv�,���VB��a���P�����&26b<yJ�����>�M�q��;����}��
]�M}D-�f��Q�_s�(���L�Yr�6��޾u3��,�y�����7��q�d=�U�%&{ʾ�o��EQZ)OFq��6U�����;��,q��<��ӎZ�6V˶Ak�f�k�^�U�{�}$
�d*g��<Qq�y��B�f
�u�US�((� >��6��F��M���_�B{�W@~o�%N]�С�sw����|���;չl(��t��3�,Q|��u%N%���<3��#G�
�FV�ϒyF��LLh-��{v6�a,��<%͜&����k�ϴF)��"�	��w��S��ӧɒO
��(�<>t��g@�:s6����Z$��r�$z�G��&����<��i�2Ȝ�elN}>�q�*����-��8y�x8u�D�E?m���)��������|R��X���_|qUn�ǁ���U�*�[{�)il�.�O�WFRX���1Nϩv;���:��e��X��R��!	�(z=�(9R)�C�"!��a�;�8�2?6 a�d��'��1wWY�K&ߵ=JwF�`H�Ɔ��[7�/^�_n��_�x��Y,KJ8R�������Ң�eI�Y��O�W�rmo��й���l���g���e)��g^X��+���9��������PV��ʧm(I���krS�Ǘ_}�Q��#k�����G�<�x�Qb���	z������}bj�BIIe��Ė����0[B�)s��c?y��B�,W���m�(���Y�=�XI��7�ES�
+�a�y�-�5)�HS|Vi����Oe�N7����tk�Vی��N2�h��7�!\Rk���Ͻ�Q� ^��`��\�ْ�*�߷?>Z?\��R�x.�4�`'|r�խ�JR`%�|��ګ�).��.�8�l��	���@h��J�AO�KC	3�'��ѣ'������b��zz.^w����c[zM�Xv�;'�3���'J ���'�� A69Hl��b嬻���*1��{+�[e���/k���:m�(�G��Nǵ?�y���7?��2&w���;w6��\ٮԜ`�*4�4���?��QE\/f�R���xɁ h^��ؾ�3�H�7���od��䦍gjG�y'�����sM���7��AA}z}����V�h0��w��|<��]�:��x��v���}	5h��+�^�t���D�i�=��R�" @���J��͊���P���4j�q����kkh/F��O�(��C"���ν�:h����<O�MV�(�T|�TB`��2��0é$e�{m%����6���{�}.>^��m{��ǝ|�豬4n�&��5tf��U���,�#�,O�e�:�g����[*uqX�n���S��S� �G/�>���=^�3bIWC_�=�S�JI�`J�̴�k�Xg��:�w/�#��g�c�ܒ�0�9<�WhE���⹝>,��V��v4�sdOx8�Gڛ�gN�3�΄�x6�|S�$Yfސa����	�8*]no�0��L9��,;�0��U�T�d����ɗ�V�_��Y@�*�͍�p ��0���U*������y����Okcpa��Laɫ�#����q�c������l��KK��ᕫa!Zȧ� ���1���#Mn������+f�n�Ԇ�вU�-�� ���}�����i��Ǭ%,0<���0t��i������m2�M�hI���S�����I���y0w(T�[_�+�Br��?dXr��g��D��>gȶUC9um����ƃ���&�����Պ[���k�Y�`g��8ɪW�0�k�Uv٧]4je�F	(�5�O����v���>5�ﮈ�gG��{�d��KK�!0?YR�j�e\G��l�?*��ϗ��������W�����H�4y���X���_�q\%V�X\���x��{u�6H#�x��?�j��fb��e��Zk�% �4������E]Mi��x�(of\�3.k;?7/�W_yU�{gϝ����@X��jh��`�?CmE&yf���z����&~�/�A�³h�1[bb��-:��L�v���֣tV�c����X�����"{I��7	���OJuыa:��(a���1��z$�����0���C��g���ii94��7��@|>�-�
��V?�T| ��(]`�O������Yпq�"H������ʄ�[K5
Da��p���_yn�k���^���&��|� �6�`��E-��!$��� ��}
e������M8q��ǂ�7�ni�Tf�2�3XQx��2�ߔ�޷�x���1�����1m;�T�r�s�so���,
���2"�sC[�O���Ҿ|Ɓ0����kU�#z��C�zI���C	Wu�^ˇ�iщ!q��.A��z�̅`�^i�!R�\d���L#ǿ��_�PĜ?z�G!K�fJ������7����|��P���?����ŋ_K����Gᛊ^š��<���j�v�ĉ��{�/�٠_�n6��j \;��[)��<-q�졃��ykD P��iXz3%GP���+�7�JcK�tSMY���ꝷ���܊JȬ+SF9��D���M%Y���?! !���/���7�,ȋ�9"��s���d��\@h�����s8��%��I(Q	�؊����R���XǱ�G���VB������qʄW�Z=�VWua��xd���H?p�Y"�ƍ��$_ ����tZ�T6N�P�ԕ���9n�+�|��p��]y(���WJgT�|m!���̊R��;���i��(����eg���J`ʧ��z���EÑ�9'�#�3ټ���L�{l������q]׵�>M�o�w�ث��H�e�q2FrG����v߇{�e�8��lK�$K�D��H�$@ z��BU�s�s����B�R��q�@�ꜽ���n#��y��g�����BZ-�J�k:�	 ��b�p�o޼ɱ�`���/�̑��%+�y���f�M�a��ڵ�[��кt�e���!�N?}���;8�0�0�8�񟉸		;�%KlT���@��G�JH0I����f��	��C�	�C�
	G��Ul)�v�o����x�u�Z��]N�.�k�*��M���mo�7��>�:jVN;�\8���������7֍�eY�X
=��F�A��{�\���R��
��^��4�q��b�A�w�^�s,#=ȹ�| ����85km�5u�÷s���-�P���д���̫���n�[o�ſ�ٰ���^q�L��=������ˑ�Fl�(��Sb�����$A9��66�B�:�܂%����g�"-q;p�O�-cv�8�S$�%��7�05�S	n��l�� ���m��ߜ;Id=�ΰF�w)�=d��fv���+����r�A&$r��q�%�.�?��C����ݾs�$��P�~�ѧ�%2�s@��|�Z���@�r�"�ƍ�P<'^gL�C�Ђ6W���+�؆�弻��!�h]��K�C&qs&t�x��BѾ99%���,�MsB���!X{ے�)����A�0�-XN(Os�rٺ�Z��q��������/lN�E�D9XBʺ�"�$b���*�4Q'�z�ݶQ4�L9�P���2p�LN�\�J2�i��J����P����W�b����������K���1&�JB>r��� ò�<��)�u/�}*Q!�ST: i1�T��������������2���ln5j~]-ee;��l�(s
�Lw���
�It�@X�I� 3�*�dDi�u�Fj4��F�=� L������BT_8������ 8�K� �Է����m�����y���d����$�@�y)#i%&�f���Ƈ,u��N�8�s���x��x8l�R�O�X�0�e=17�T��8)���cl�����E�;Ƶ8xA��0�|���;�K�}���x��IV<��k�*܇]��nl����!?S�R��L`�n�'ߛ��X��k�i�2M>Z�#��&\�煖�RF���!���Y-D��`�	Z`��=�)yK�ЇE��%�MC�*L@e&ٟ�M��u��<2��x!�!��4��;\��̤٠i�A'w��6�'
K��yn�-%C+I!�#,8�0���T��d�˱ <1���KZ[h9�]V�� �G�a'Ԫgҵ�1K��+���6bjQJl�g�����Z���EY-D��3�U�Z\ݐi����r�'cg�ec���=/�^�ڇ����ڭ$
@���x�=�sMM�0�&|*�Z ����&q@3c3$�]JýW"2���}LJ�����E���V}���ٻ?s���ן�jr�WL����@�}��Iw��&(9�*�k�Ji���Vڨ<7���2�8�%�� �۹,X�Tpb"s�,�2�����h�xUM(M�.=���L+ܫ�Q�Y̘�=����a��~=�ZYbap����դ��2n�{ �����W�@����u���ns�g�+	�1
�T�zއ���8��둨�͵���[�B��<�C=$*�ڻ�|.]�����c�/
�s �	�K/���X��x<k�Ӳ��L<*��$�d"K����Ah,�W�~(3��.���L!�U�o�|�Cq3xh�h��qT(*D��z�ݒ������X�j�.�9p� ��]4
3%&��
���X#�n��W4~���� ���??y��]2+�\���$��A|��L希�AM��j�ȁd���;L�@��n����pQ�fX]sr|�
���P������[����ך��rC�5���~��J��]��U)`d�]Ν5�'+��,�
�)\���o�G�!��Mf�`&o��#y+�)>?�,�^+UR9g���f�Et�xٚ���{���J9;����2�94��I.�6�8�kwc���='�ʍ�X�������8M�D��g��%|>��3��'��ݝ6�:�=U���c"ԣ��iއ�I��;p�y.�U�zJ�贼UZ���9�TzJ�^WS�����f��!����Gn
����B�b �����p(|��Mo�WCb�6� �r(�����Ó	̒�rWM`2^�4�hw�؆e�ΒoC��q���G���1.���6غ�Ȩ+�F^�DF,:Jq���uo��ݵ�z���?`>2�޲C�;��@�p��c�IX0�!ƶqC�U��X�%f��X�:��/Nt}ߕe��ߔ�)�(�1��;	���j�S���\H�-�l}��i��u]�_�{c���L2Ö�&���h�U��C��l�L�^w��.k�?r/��(���M�K"r�+���N��:���mc�k���q�ж	����:S�������7a�����I,
^ep��i���� ����a�h���*iR��H���A&u|G40����>��m\ꬱ�r�24�!�� �����-IN�a�J�Ja�,�,N���M�0�* ��v ��a\:l����a�z͋�d�����I=���s���'˜�Ŷ��-�eC��]��,Bp׷���v6:����
��[��"�w��x�}-�����6�)��:���	JkU�ҏ���� �mQj\-��JQ�J	��VU�I�vnE����feY��t$j��+T�y��L�AzNCn���QI;���!Y�9�uKKO�]!+�d��㵒�ZX\P(u�*u����s���rD�D��묅��(�W	M$�}&�D�k����%�H!�%cg�[��ԍ" |���#C80 :�-�y1��p7qZ�1o0����jXd҅�����.g|��/���? hH]Ll�LfSR=+}��&aA�M��I�_��ὂ+���C��P���H����)ڹ�/劺�;Ye��?�%!Ep]�.I1WǪi������x�%������x�J�i��r�]V�{FΡ���1�%�p���VS�PD�@�3et�;*�[�gE����2Ö�lr�N����m�r<t͜��^�S]�{��~��H��c���L�H)(|&>��!��B����P%%�DY�������2ˢ{*/(�6H�4G2m�fr
��1v���]�k��$���#��7�y#�?��ϼ1�4�� \8�_�e��$��T��+��঱� �KL�H]�Q�z=�xv�݀��U�,�Ki��f������+iJ(�C�]�Ǒ	/�F����E�h����4�\�z��O�8��<u�}���	(�$�gAy^ɼ�HO�391�<��8�ͥsV�����t�a���ӟQ�q��T��;5%TA@�Ɂ�F�P [�Z���
��uB<��0�� ͖����b��B*�$d�F�t_�*	�l_�R@L��2�j�r��vX��lM{m2��wX��t�v{�1���q~�*K� �?S-��dL��K-l��=G�1�`팲A��J�dE��/��-��LcA�H�����L"�Boll����+R�p�S>�aMy���c�{���\$D����X��e�� ژ�-���Ӏ�	$)u�Ɍ)J�Y��P)TY��D)�M�C9Kˍx��K9��Ȣ"&�_��k��{�w��I����*��k��x��6��$���S�eR����_�u���NS;I�-�λW^y�ޙe�����a�����n
~Y�?X�'���fZӇyw��j`�����u�42�؝*2s��``|�'>r�[kh��Y1��%fIS\��u�y�$a+D��?��37?�PEl���O�7��m���ߘ��;z�}�U Q�φR�%ǚ	�A�ބ�m�PSyKI��}!�8���Ǚ���B��	���l^1��p-X_���͒���1��v�ە �±��ɠ>'�!ۄ�&<,�hI�&I�������!�1n�,�."kNOƸ�Zl�m��eRq�(�b������	)�a�>�ob\�~������m�(�D���ȞAB<0��wy��C��矻GѢ��/j���U2I\"%T|6{>K���;֎E1�A/��Fr��?�y�A���*M|Ȼ��ƛ<' �:l�},K���;��mXZZ&���P�_|�%���X���˯��88ޟ/#�#�.�E %�0�?S�|� �6@��u�z��0+$�A�2���k){�����H���?/�Pj8�;�C��K���I�ឱVss�>�2˺��-�zĩ+!�L����*`�%�t��z��X�V��,�#�=����(��W^e|��[�a|p��%UgZ���Nfi�u��lU�B��h��ЈR�[`�ބޒi�lԽ�n�(0��z�^xQCE��ن����lskݭ�>a2�� ���kk[-x˵�f�����{��06-'�7:"�j���▱�dG��o����Wcqdy����0�awW�TF�g<Z�`�0��bG�>��p��x/(��h�/�>����Q�Yc�{	�^�WW�Q����^�3�9�����)l��w���l�m��!�.�>��Ӳ�ՉqI�G�]��i�߫y"� ����k���n�o�;�r�������L����$2p�P[�xj�7½/�����u�a�|�#G8Ǩ%�/�*���x�׮_s�׿v�O��G�x��Nql�|�T��pŃOk�Z���P�C";)?XV�	��H�@\�IM�hi���{n6�S�`�!�'�t�3�[�>t(4t�&^_F�{��Xs~�Gw��Ur�]�~ŝ=s��esx:r�`&�[�'fݩg��Y!� �im=�R����!.�X˔��h�3B~G(�`��:�=��c�+iG��pI�h��&qa;Ąp-Q��!�
�,�xzcw�{����M
��)-k�(���/��X�' ��j��xO>�I����}��Ϧ��~|4���0�$�;�Br�'�x�Q�=������޸~��n��ܹ�-�V$��0k� "g��8/K�̀a��~�	%�C�m+`�	G`}�=�T��#���95��8@Ҳ8+$D�3�,��Õ�)���"�^Ƀ����i��}B_�߰c��>'b <�� �-��9�6"VZ�H��Q�㲒	�I)�S<C��K��&����c�����:�|p�羻���������w���v)ػ;{�3��'��vW^�.Y]�����cnlC�D��4���X*����p7�dV�OX���C�=�ӟ�Da�0�����QCK�a���77��p!�a��@��1�����@I��ʀ��`tX�*x�Рa�
���c��ăϲ����{@1,�/<p:�B�lU��n\LR����k���"�9o���t{{��VP��W�D���m��F�a�=aM���FkmmM�p#l��;j�O[�4�Xpk�U�&t�:����]�X�5�<k1EopM2G����%��7wi�7��Å� ����% ��7՟�x�[g8e�c��4k��l�y���]�SI;���{l�g���n�%�vP�[�R�1F���vEi6��a���f�����6����/��sa֭{w�����@� ��������ڟ?�����'7 �ݸrL��]p�]����^�(�3����AF3M]op��yA��:�B[,�;�`�@�k�4!� v�{`��b���P�KXv���n!TVX8<� @���b��y0(F��JXr�+A������Gy5�M �9�*�p����n�ٺW��1I�������&[���}
5�˚7�n�mV�c��ǁ:q�$���%��ߙG$�U��g>�)I���Cj&cS(�C�ĸ���،q2,�l�y3�x0�lt�X~��+�_{�5%E��7��!e��V)5Iau���$�7���$G
�*e��_:z��9Q�z���z�X�#4Ҵ��õ8�rҽt��A95����f�r�e�'��E����k���n{m�=�%���q���� ���/���'�]1�b���N�k�+J����6��h5zQ��y���s��ƣEB����	-�c���ͯ�^P��\$�^��!s��G�p[��	0��� ' �7>�DH!;�\C�ah,Ă����P�Z�L`��0������Qj*Y�T�eOz��� qy�{��|L�����$ �#lų��4�Z���X1���x�8�lj�?�Sz#�!Ǹ�KhP,�XK�9Í�<ddW�)]�ޖ�."а�x�6'vpQq�n\��M� Z��x�K�.1Q&����ś�N�D�	�Ƅ�u��%�A}��֞2I��Ĩ3
����g��83�:�3-Qȑo�cȟ+��g��R\ݢ�w6nh;	#���Ӝ:y�愛��?3[��~�}vj�B=39�_}�ݽ��{��=��K��ܼ�#7��U��2��N�Z��{EK(s���%l%)�;a'-G_
��k�����>>H�7��b�	V�
�|�R���V�P�R({��0�zᬢ��{�̘;o�0��!{��.�e�\�=f�q�j�=�){�С���y#���O1wB���(�_��'���{�5��6 ��I�px�*�֨��R���3��fR0�����a��B(��p[Q�'�0�dvpl �{��w�ds�'m��b� �Ǳ�����p��O�� �1\� �r���3���CK� y�)R��#e�\]�:`��-=�Z �C2¦�
�(�Sە�P[W B��Lw���I��'H�L���ioa����������r��6V3��k��ɪ[_��Ϲ�&2/�P��A�٘;6?�*���=Y�g��n'��R�H��{����L��EA4Jeŷ��G�Q梐�,�c!N�X�գ``��	��I��-����|FfYi�)5Q'��f@�"�*��1���M��F��bpB�=�g��e���w��@�C$�x`�>��O�[X�����?��������b0ײ�$��Ωs=��11��v��#|���s���12� F����� ]%�_�)}B:�w��Cf%�@-^!���P��Q����/JK��[��48ţW��m�sJ�35��$�A�&�0�E=����wW��&m�
�_x��f����\O���u�C�����L� ������3�Ի�C����qc������6��Ʋ߸��⬔!k;��1�B����6N\�����E5����>�L?����H������6V7̚���ҳe��r���!	j�!�'�(4h���lo�
���䑍�1A6V��;�,��5gs�q�p����ɳ����F�s�a��n�����&��Xa~W>�&�T�JG-�C���
4�8�	�+y�cK�3�$�l܂�!b�j���w�����)��̖�^�H$W�{H`�"(�����!XCR���8��CJ�~���ӧ�0�kM���!��!�T2������8!� {��!���l����;� ��ѿђXV��d&�xx�ӧ�{a��m��`ݭ>y���Ã�3*w��e�ګ��K>�9<�������Sc�ݭ5����ݲw�<)rPʺ	���˚�^N��
S~D����E�d�cB0�P�{Z&�\KcY�n>|���R��#��cv[�ѸU��$
�G+X��Nk�ːc�}7k�3�"M��}����"\��0����U(X<�͚).��!C��C�a�{�Δ��Q�29U��̄σ�G����$���SO�%<H-I-#��C|hI�<vp�;������ ��?��1-�ڒH�<!�f-��&rbM4h4 �W�\q�Ο��E:��;hU㿖.���$N���g��	�93ta�8K�yWS=���B�ɥ��!��>Y~�r�[�m7�����_�͵w�آ[ ��WV׮\v��z�+���8힮<s�|�ƒ�1L�,���VX���i����0��$`�.�:��y4|x�e����g�z���R
[m�đ�t���`��U����� �G�����e��"0����+��2(#|BN?@b���l��"�$&�������+G	��P�wd����c����a
 ^�o�K�$!�0�@�����[���o^�!�J�~��B�{�b#����~�´�e�#�S���_6ԍi����lȲ��QƍPjb>�YD��^���{睷ݥ�_�" ŋN��nbj�q*�ö��135���	w��1��l���U(�=yb�%�q��D����d69�ύ�q��|Pƀ]�/����ݾy��L`�9srΝ;����W�5���[�h����ao����{��ʡ_�G���N���cnsk�MMc��	���P�B�{X(��esڇ'�(�Y=�5�Q���R����j[�"e�1+"�݈���+m5�nޘK�.���p؃����
c{Vr��6XF%�>�{�Ur\�HΜ>붶7�c�4�2��c��<NVնcd�?���l�eו��E� !;��ƤK�u����򠴰V�x=��ޫ8���c��1��zØ���3E�IHJ�Q��q\����
4;�Z��*�S�g���Ƹ-j&<T]�X�iF��5Zj���`��1�{l�^�v�z/8�fa���d�@�*J;k^�o�\��kd�ۛ�����p{�4G=ؐq�
I虆k����}M� ��.��lŬz2;{n渿�)�./�ӧN���Y?��~������[�|F����I�����2v,=E����|¹��]6���*���M%�^;�T�����/B�^��(����{*��Fa�)����c�X4�	n�H�^����k°d�|f�����όcn
����������}�kb1 �d�ij�s�% �z�o���a�9����� ����1��d�e�!�,��^ǿ�W�-xT������}���'@Vr���χ�]2�t�z I��ƣ2]8���Du��GY-.�.�ƽ1H7�k	<�5���2���n�8DAqH\����nz|a�θ�v0W�_�w����c�����;�>�����],j�ք����gVy�����[o[�Q��1�z�R}K(���:���d f?p����`�%�~�4c�,�_�Սo���x|��}����z��J�Q�EΣ�e)*k��Y]�>Kc�ﻄ�	]O������ >�.Ka�����=�k��\��&:ʛ����VδD���/_bMĚp��=�a����y������kj���K-���}��Wr�1V'�&G�YXt�ٯ�����R�C|��Y�Y|i�4��y6!�I1�a��h5�$3���M�ȃ��/ڿ��f��J4��i�����$�xC�:d��;�G@ia>��~��<ay�= �& ^��3[�8�ޢ}���~�sj�Л=x��O�GY��`�{�r��K��̱���1�ps��P��)A(�G4n�⌲�_�3��{��3���@ݸ"q}9u��<�3�����2�n??VDk��B\d$aUm����o�0�ߺF���KZ��Jcy��xn������/��8�`u9�,Q*���n�����Z�n��dNa���d�W�r����D�Ď�L�i��}q��;.o�E~ܟq�PH�����%�j"t���e.�Qո,�BA"���؄�:%
��2B����\'�Q�!��x�YW,ܛ��i��Յ��j�Z�{x�M�D������s\`�*vv��u{�v<�ᇨ����Ԋ~��u����pi/n�}���*]���噸�j�6�T��V����U�,�����V+hFb��Y��ܭ%wa�RN�a�j�[;b1c"L�j�<p���S:}��@�&�?d��O��eI3+#Y9�34��{��� �)��W�`�]Q���	�	5L���/�O~�z��;�����O>��}�����po��bn�s/��5܋^���qWk��!�����^����ɍ[�U[V`�ƅ�%ל$	�� �E�"VK��0��Y�G�ax�B�׵U�@�!(��'U�-Wx�۵n����͸Y7Ŏ'@��
��PI�51�� ���b�z���{Q��9Ѡ!�Ե��Z����KL*Z ���j��%��rz����vК� 2��2�vc��r�L�tJ5Մ��ņ/J�97����e]qٰw$��<�,�_����k�|��������SlX�_����g��ݽ!�Y���D8����0a=�"߸�{����=�����j� ;Ǹ|oW:ոg��	J��q�����=(����%S�]�4y���d���qs5Ɣ�Ԑ3�V��Nz	�m��c�aŐ8l��L|@� �~(8�$���_\Ud�R�q����A&�mc�B��XB��k@��� 9;�[d7AɫO�P,}�&
l!�e�`R���Cf���"�栃��e�c���WEWL�@vS����dAr�.�j8�d�M��[f_E�m�X���4	�Ccj�O��؁��?�)1�������|��}%�Qk�}�&�,,I������~�(�ju:i,�r��/�X�qv b�� ޻���ϟg��k�x����sg�8�2�~�_ȑ�t�$/�@�q�8��g@�Kj���0d�Qd�X�<I�P�p z)BI+M @?�KDᖘ��hp���P�g����wA�g~�ȡ��8��z���P8�G9��xi�E�x)�hp�끰j��E�0=�����)��6�	�0�:lf��<K�;2�l�X[��ћ��c�pr\����y=��*˖.��P��%4>.��a�TE�s�����`Q���V��3�����x�27Nd�����܌]V�O�
c([�_��ȕ���W����.���~����Ԝ ��SW*��*d�R��9U�,�$� �+�9�K���̮&?�D���Z���Jp�N�����	V*����DS�t�G:Ɩ��'�t�f�i�9�U��5&�Zl�ט6�{�M� ��Ϩ������7���`������+ �����Pvb���1NqK, .Fm�EtZ���!����B>V�*H2�)p��:栳�Q�k5�|0�'������H���4��E�4���=���1�0��y�]���3�^��g�����֟<!]X���7(G42���E�L��$tq{��&}�arg�<)M�=A*$��U���{��0�e,쏍)���.��a���o�(d[��{�����g����O
,+j�dLuy�qƕBL-���+�3�9�q�;w�4�;k�3"���;�kau6����/M��&>�|��RB-S#gIʐ�̔���?��Z �&C��ڢ1<u:����\��A)X�7�3�;րc�jx��?�s���^��}ѻ� <�g��d�Ҙ��}�����2c8�1j"�d�qcsG�O�;����˞s�Z���^~\���jj�)���@��U��y���������ʋ���W�`�x�-�p#1���P�1�4�E���[[r�-�3������u8�f�	�%�5F�:���߹�;�<-[=�=��fpe�08��8�F˅g��L�8c�
a<����:Ho�41�utm}��鋴��4z���GP?T�A��e�ϗ1�M�t3٬�(����囮�^�.�6����n<L��S�៝��M��EE��d�����,�E�����Ν�b�Ͷ�]P����%��RIm��.�j�|k�ckLݏB��x|/?+Ts
FOk��3�sL��Iɧil��`�yX�Ӳ���J;�rc���g a�7醁\�IC����]�z�]��2I� 1Ć]�t���1����>u���pm�4!�&����E��P�m�C�=ɨF�X��$XG�ƈMm��ƣ�%�&u��3�á��<G��dJ���Vho� �����W`����'I)�~�]+��k��Cf�5�XA 3��Fgg���w����ԅpq���U�dF[�{[� Ԧ0�y9�p �^*����h��P�2�e9\%�R8�R�i��>,�Sha�L7t�8�QY�,�'��n��m������k[������T��_6��>y�;��v��L�-��+b�����
�ZO��[�����ѵR��i�~2��gu��K������H��3��L��ae�z�ϟ=�xjs�9ozʽ�];�NM��$�Z����*O�F�|RAy��kJQJ#�T]�)�S#)xQ��"E�&�Ҥ�q��r���~�`�mn8��=�_ƿ���e��T1��@�=|�Ȼާ��0Í�A�����ٸa/���̾�����/X[oi�0'5$U��2fSX`�-��K��ph�D�P�Mġl��d?�A� �^������kas@MO��-��%��wϻb�M�}��ϒ�O�UF�4��X�P����1�A�Ͽ��5@�� 42]E;��4��Nj��_u�9�ވ�'[i�%����#��?y|��lA����nm����R���/�Y�M�������`a�e��x?���V��+�t�_��M�!bJ3� D�2���}���� �k:(�/���Ng�`�u��*I�,��������w48�p�JH9����Nڈ,���"�]`@�Ai��������$((��~����n6���P,��P�����ta�ޒ�������C�0�`��W�����1 �x���]�:D/��$Eps����f
�I?���ф�?/̚,�1� �A���'�Q�jq�k��M3�]���9��Kxm��@�s��DN-��ײ�ܳ����к�Kn��\{�O�c�����naq^���>���ron��=��}�ܡiv�6h�q��(������'ݜW�@��`����=Y~�uoԛ��獒):�������g�}���&9;��SXg�2lt8h#;,֨�����{���T�ͨ�0�_0B`��=�hX�vB��[3
,���Z7�|C0B#xNh���_��MI�t_������.í��ِ'���M�0����q�i�Y�8�Q]jf6 ��F�}2I��fm�h{����5"���C��'�|��߿/Yg���,��!���>[����^���>v�Ξ�{Ȇ�n�r6^��JP21c_�؛]T���L ^�e=Z�u�r�Z��嘴�^E�����v��ew��*��������dv��n7�J�~���!8歳���t�ga�e��H���J=���݈����Lin!�RH:�ʟ���c�]G�n�%��ft�,}�#�Z�4Y9j���y��&��B:(!P	#l�de�i�^ӶFc85� V�q��BiÐQv����-��
���?��n8&�n��D���<,���E�ܪO�h�n,\0koY|c��ԇ^��{qZ�{8�cgu��|��m�Y��zY�r��g��A�O�,�������V�@�1��a�r�ۄ���t�y7�䉿�r2�q	*L��C�Q��Gn�@�s�#&��?���kz��ج��V�n��8�4(��fe�=*�����p�>N�aGڜ;�]s<݁��=t=�N������B�X�`������h"�/Z���^�W0oL�9Z��=s���O�&y�����-Z�6�٦HR���{�QB<*Y6� ��V���!@ ���A�>���4J�;k���ZT�,��W�U:Xa�w�B������ۚ�r33��%�6��L����C~��ƕ-�°�F<hF��T8��ˍIʺ=XGE�i.{�T���S����QkH�G~0��-(W���{tC XH����{L�������o����u�����&O 	���ü��J>���R�n��/qFN0G�jI�m�}����bG���Hs=��J��ć�ݑ��`���975��6Rt��no*�Զ��s��9h�M����nv`������]�M�� 0�%Z������\x:��-��W(ay��k��^ GG�{x�d-e���i(�l��ʋ�bxK.�]x$�����_u�K M�L.B��L��9��g�)�s��PRs�a���!�b�s�2��[�{����)� <:䄐IGK�ӕ�@�h��y�Y��`�Вhn�L�k{��a�lGD<86��ƕR�v�	�,D�gN���{�t��,�n;tBA#�&��$l��Ҧ�-�3��=6 ��H�%�s:��o�����}7Z�Ղ�Jf��V{��>�&�im0-w�tƵ�Wq�׭�&�g�p��5E��l/���Vܘ1Jw�KKn��c73;��aY�[p3s�tsQ�&�#��	���v��o�e�Tr�zQIh��F���<i�o�7.����K�a�z�:ݍ(���,4i6?%U���TpӼ�o��Kk��� �˄��յ{�5���q�Q���Z����moi/xe������w�O�2{wg���> �c �����d�o��g�{{��4B�5)��W�Y��a	�	�*
����u��dTE�6����e�z�5���/� �0�������F�����Km��;�/n�S�8�^�P��
_��������nK"��2l����"�r��b�$��
�yÙV�J��4iH*]o5[03R/����aJ�>]e�B�d�k�Xk$-��Μ:)3�����z��m�0b,o��I�I����(��	�k�vփ����W,8<\T�M,�X� {�Lxʒ�
���Ӄ|4V��d������ �S4��~�������O���m)�	��M6@����5.�8�.��X���Sd=����x�i%�߻O�D�o�"�n%�n3��s$y�o����[nٻ�P6ۨ9�l.ﭭP����b�8j����w�C���n��{=��]e:<����`C׈�T?��zf�pgΜ#M� ����9@�`m��I��+�h��S+#�.�q;Ճ�FD�-#GJ%�� JS�}�D
�H�F���!��q�0�C�Uw� �^����e��.ͦx�Bo�ĨXQXb"���ǟ>~��ܾ���fH��2ݎ���Ңw�~��[���|�
��{�pt��[{����|}�g2��1!*����V9�8a
��׭B\mSAM���EBw�f���_^�x#�NP��zA���x~tOu����Z~-!�������,>�<�u-&����cχ�#c�£���3��x��jm��ZF]�@�j)Gh��=��в+��������(���x�8��B�����ȹ����s��ܴ�9�M8�(#�E�%�:�Ǘ��jH���i/�ǽ��[��D�����,��؇J7+1�iY?� �<Ǫ����6@s}w�5ե˗�8n].rx4�jd���V��n-�(�)K �v1��4�=��]�	�\�ǔ�A�Q�LY��i�\z��+3�A�,�9lцQM�[#�w���=���V7� ��{�ܿK�e�H�Y�	��t���n�&s������u}@��˅1�m&+s�$ϡу ��p��ZB�D3���z^�7�0����&�d͆�����Rk�ۄ���~�U���y9&�&�闽.�>ײS/(��|�Ynb��:�J�[����l�A�\��\鈑���b�+�9��=��U-2��ճ�gnwk�]����Q�9A��K��~e��EE�_5z�^�Z<U 9kN��4w��L!F��?JQZ�PP	��l� &�t@ڄ�$��V�^�I�K��9�X���<e�_�/_�{-�+�i�:D#�Y�
D��D�D�;�
��b��0�nr&ipu���*�;�7U�j�3s3A`���o��Q��hWP�$����5���N��>��������<� �_~���{&�V�[�}L=��s�u��{��I(�J���6-1��؜  ��IDAT���Y�)'��EA8�p��ɋ�q����&�b�F��=��y���??�UL(M��4(���=�ú�B�s�K��a�V�w�@N�_��_�l<��� �����Ef�.�ӕ��# ��+�GK���䴰� ������}���K���p�g�6u�9�$=+��,��s���gUDbu�86�G�K2>�W����p�ի�X�6��T�����m#����e2!"�̕�|�Ze#����&�`�)���ȃ�.X
��K%�o�jwK��YR�j�ϻ,��r�c�*�Z���ze'�Ҧ�67�`wY��e~��A�RM��5 e:����y>y��}��Oɔ��CN��n�@!�cPGK=J�-)�ڋ8+�%}S�X+X-����MvT��mi��&��+>薛'�>G<J�e7�۔�{�����]p���G�;#���,5�ox�֎�{�����~�{wﻻnv~�����D��|��7D��z���֙�zg�3��Ǚ��ː���p��
�{l9֬]�n�75U7�B�K��� ��������>u�)]���C����j*���'&G
HHD�!v#r���;b�M���`3���5˜r��./5N˭����~f�.�/���C��h-���%[�4����'M�9U��֐Tl|��$q?P�I�H���Q���p���@���c���{����C-�Aܱ�v��J�M��r*4����H�r��' �Lɍ�A�|~^~�;S4��Ħ�*i;��elS2P<BDQ,�����3|���7�`_�K�2�Y_�`��nm�^f��ԗkE:����{����~|���3r>�"� ̵\���h���Z8`��G��2�?C�hm�T^xCt���W�KLi��"kRb�Z��&	;�lqcX45�
_��Ǐ���}�A�u"F��9��@7��6�A��q3��nѻ��?��^%]�	�be���Gd!�'�Z���BWe�cZ��Z�粦R�kmɓ���2	O�]ǽ���oZcu�t��1�����mt�5�	�����3dH����Wr5�:�G�|ђ8�7��Q��Y-9�b�lPa\� �M�2�h���]���9J���D�� Ա"a�@5=j����%n�ɸ_(����	�����R��0wPQ�ZX;�M��TiW��bϤ����{]�8��T������EW�����5���1�'��
^G#�H��$"�S[Y+tsC�B1�8չ�R��E��>\5DUE�D#ž�/�e;7��i<��^�M�Ve�({�$�p��*���x����|�n���76��rB'����h��+��Z���pC�����oP4p\5A�e��s]K�Y�4�T��a-@�����k�?��h])����f�y/�F%�3_tŤY�3I��g���p� W`���g��sGy����b�ިD��Ƽ
��c��N��gS�?��s��?������<{�m�2���nz��"�8�o+��x�1c�O�E��Qp�]���Q8m9�g��������8��J��{���WYf
��7,�F�=w&ԒCؠd�ܾ���BS2� ���t7�\�U���g
��8ϼf�ͪ��1u`���-9!qB6�n��u&��:�FhM��;ky\)�$=��·�D�e�Qb�F,x.�t�0���b@r����V��,1�9K�H"����p�"���Aɳ4�I��9�ZD{��3��$�ތUJ��`PzUs���|Y�,���Ӭ��6�źֳ�*�(�v�Zb�%u����U�_�`)��B�
�Dİ`�I���"�k�@���P
p��樒�IXv�>�R�)BCATւV��:ape%�������Y�KXU�T���f�d
j�lb2Aq� ;��hǦ�&�$�f/0Z��`�C�\:Χ�{����n��z��@����Zi�ĭF٨g�8�މ2��%��8*���	��ӄA+�Do��� �vL���v�1)ǃ�Zj���'R������Eτ����T����Ń1I�G�tɇ@���U�Y7�[N<� �����TH��@�[�U���d��@����t����[�3$6�{O^"B3�5���<�>�u���
�%��׮_%�첿w���>���pc,�e��ղ(\��]��ͻ��I�r ���D%H>_��aI9���D�G���Цl�҆@�o��c��Ϙx%!�}f�y���
�2���Z瑸�uH�[�U7�3Ν� �PO:�72̶��0��"Dk����Z۶w�g�f��SgS�`i,>�*ٲ&3�|L�c��Y�N!������R3\���6>WD��ÝAZ���{ԵK@�78��+l��`��|��Ξ;�߸��j2�2�;�ḋ���;w�|��@�a:\ʅ�*ҵ�����(q��x:��	\�B�5��ψ;fY����L�\�1*���H����?$�����>װ����̀�� d�;� ����^O��$���5J.�B�SV�[2�|����ƫ��>y��	�|#<���;nyiY����<5�Ξ9�8����R��l\r)���C�@2����Sk�d���S9+-��S3Lx
�'�ގ+�L}ejV�U�%�8���X��nôљbM����&Z�鄿�mnm��<t�^�"I�Ac�~t�h�Aa��� <[[g������'����9Zm�&�)R���y�QM�V�8�1�H �B�I��q��;[����<`�L���kb�+�rz�ݾ}��p�/�J+E��D��l��9��X~����K���!OE,���d�P�[�R���1�p���p�Gß�CAP%;K�Y�i�i��f�t���B �i���#.A޳г�R�Y��ʍ���˗^v���_��W/3�9���Y1@gϜs��������虡a�y<bE��&�r�(f��s�H���{̒3o�	?��d�%)�	�2MBۂI�V0{�٘Q �'�m������h�%��T�׿��+�o��o�rf�+�n���	�o�����,��z[2@��۫H��W:���l0BԚ���;pb��յg�\�r�c�h|\��]/��I뚸�A�����d2�H��{<L J 9­�_)X�rW._r'�c�(v��rλqc��3ӓ��	̎0��Y7�?���$��!�xd3�8��x�\<�*0y�=�o��&���!�a\��x�<����^��V�c�O�(.y�a�3�̛���eG��]� 0�^��?[@2��􉠔R�){�f#�J�>���S�O�0�2�w �D�������V����m�LJ:�/,|���CR	���4Z�1m!�E�U�ix�Y~��mi�R}�8(�U�<�P�^%Rfm4,���ߒ! t� ���E,b�K�B���TC�;.��Uou1�R2׽ ��F�	��H���?���]>�PG�]Yd�II����n�ِ��>����DR<D�Xd=@PD��	�	3��>n����gv�PzM����6�2�\8��`�����̻{��Ϲ��&�2A� |���|\~�������8�W�����?�D��x1}�I��8���/�[�X�QIţ�!ޅ�*�Z=e�*�{�9GI�� �n��7����+W�P}��O�4��F���a����,�v�a�Nn�����n��1�� �Y�a�T0�S�����cff�[f��g K1����nC|zp�\�'�p K�
���6��^](�~�Y���;6u>f ��޽{�7�	��x$�>�����1>G��c�c�o�M�<���m�$��i���~�K� �!d
�!�-�6�����m8�4^�Q5Gc�Qs�`�;�{$�&����e�;4?(d���p���¢�I/����>O���]���g��C�B�>sʝ8����?q�k�>Npx`#���l62��X7.��ǵq?�G_#	�q`��J�waub�h�3F�{��I�m��<�����N���&)95.���H8���{�_Eps�ɇ����v�a]�,��Jէ�N�>�n}}���?��{�ͷ��k�����+x�M�ڰ	��NnA�?G�&��t����{�d\�����6��$Xrl�n����^��$i9I:B� ���zZG���L�XO�K
�}�/�_~Ɏ�^H���
f<StXo�'h4H4���:�4�P[i�H�e"��,�H4��-a3�4�U�X�y�d����.z�n�K0qnv�o𛴪8(�[ ���/]d����u�T�kk����������k�¹\_�*��IBg����f��'ZN��z�_ ��#
�4Dw��qR-����b���o�6_�n�J�3�,δ���������Ѣ��?k�"�p�N���w�֑5�"�����m
�`,!I·�f~�>��=Zz�^y�U*f9���[7oz%��^��,�	�Y��=\���-`[.H4�Ki8B~ް�lB�!��]���1��iS�h�~pUp8�Yn��a�M310�� =o��{��?�Y,H��׼�������~�Ήn�r�ze�����������Z��@D�p�v��aً	����N�r:����1�&j���̈́ͅ"��Xz~v�]�������M@��ƀ�/������Pi�=�y��{��)��739���v���c*[d§&��#f�= gha[��OF���n8�ູ�{ŹTiRʄ����+l�������p�f��Ŀ��c�!%���Z.����aȘ��Fܯ��A���<�U��&X���_{�5w��9�
�o��5��i��(�tW3n|g}�(����!�0Q���Z�3s:&��-���2޸ݧYo���o<T����H�`�����l�mB�&��Cmӻ�� ���I�V���(i9m�cwV5���攒������L���L�ފ�Vn�Z��t��l��7��T4��<�Jc�e�L�;]��*����ur�����x�8]i(1��3>������nav�M�&�'է�#�;�αy��DJ��%�pA(��᎛�=/O �(�dL���e���,ֆc^�:�F	�p.���+�����[�F�;9�L+Q�r'�{�����lU�-$�)D�w�4,B��i�I��𢰗k��(?����8*���#f � �MP��t�a��>ȂWռ���\�Ƹ�7��I	�:O��Bb$�ߦy�ۛ[���w�@AK�ܣ�e�XG�����{wٴ/L��Nk��U�4ΰ�� Ĺ϶iƩoB(k{�[I�k�*h��	��t�Fe�G]ϫ��3����6��}ȱ+s�ӜG}��1R�3��ñ�s�N�8�N�<����G1��2�]m���*�}� �m�F?�	[��aor���9��?
�4E;��V�&���B,��4~�	5�}43?�l�p���8����p�4g����4�`�:>��y��B�W���֚Yh��b�8_S	�ߣ�|��M���)��K�.�W��
,��ў��P��w,��B���]o��7N��L٪�:��`��vj�Ub�k���\aE,dvϘ �￰�����4��C����-����XP� ��L���1q��e;�QUn��bݚ���/Ukߍ F0��+��v�Ȕ��a�R�-��R⮂�7��a�N����-��8)�+�J�h��{o�Xg�f�2�h�{58\�_�5��`��37�]�K�Mߢg���w���w��������c�-�+"�p��Ir�~�z�g��)���+��
�%b�=K���y�����R�.��#_y!\Z��k�e��%��PP��NNN���K e��-�� {������>u8{�c��٥������lĵ�l��}��#/h��!�� ,�4f��WH����J�+y�W�h=q��Z�	�t��k>��{y���͝oݣy?2g}�^����'὎�-��i�(�#��+����P���ވ��Z�^b�Pzɔ�ܰ�H6�{ dp��^=x� ?/�n��<�X7��˗�����=.��B]��s�γ���ͯ�r�`&�i (l��uq�h69y8(yj52�/�<׈�����[��Ƀ��`����� ���x�h<��d�Y� �l����jV2�������o�n�����N��.1c���s�{�ݶg�Шm�������>a��`�+���-�hi�
�il�H
R��M�jԖ�u����-�A������*��tqH\|!�Y���&��FBP�B�obһ�^�F)o�[<懝9}�-/=&'����*y���4�k׮q�����݅��X~���{�����}�~����EƵx@haŐ}�|�e�ֿ�Ϳ���԰4�g�S<�;��L�-�|�uC8������w�Ozok|r�]�|��w�ޣ[^xˌ֙��Y�<d��1�e0���s��Y2�mo���p��{�~=���b�_ҕ({H+�4c���e�Z!��J���:��Ԇ;�K�j��b�s���:Ã��&�s��X� (�nq��n_�ɰ���^�+=�f������n����e�܍��R� S�@>��t�n�`c}$���������Z-)�����A���F-���c�!L!J�{K��󡌇���RE#&`�s�l*h� F�^M��U9���D*�GpT"Χ!V��2P�>�v�a��'�fӭcM�VN�.�:L���a]����o�M�㚁R)0��o\sO���b���v@C�/X3Xу�ߨ!�Ⱥ��CX!ˏ�Y��C�W�����,W�u�\��A��, �RH���8���+=_�&���ήL��`��~����{�W_�����.��\p�#��|��Ξ[i���&v_�@�u���Mq������`ʮW�;0��po2%۬����𹾀	����t���k�[��j�mxW�&�~9_ߡP!A�
w�޽��y,(eX\�Z�N$����H����&��j�����!Œ����v�@�Ĳʟ
S�mdZ��{Ix8�O������"5q���P��%��H�euii���3���1tW��;\�I��`#]_ߡ[==}@�	s��F��;(�:�-$s��K��!1,�D�{U�c���L$�O�T�*�2��Ij���f����0{�f�]iim�T�C_���	�'�p#ىߣ�A�=؀E<����$$~w�����!L�C�Ȧh��pC��ڍ�
Z��D�eE�@[ՆB�$خ�C<q_��K/]��CRNam$i<�=�zwWC`�9�
�������{M}6瞬<�0�
�.+�o��f�8����>�C̶��v�w1p��z5�Z��DC�-��nP:�0T\�������.�@�#I����i�k�Z�A]檒�6���l�(���*�?�wi��>/MڌR)�Ƽ����]�� p;�����ǂ|����+a�7�~������bܕ�-�ec^V.���[�[�w#L6]=�Li�S��]HZK'f��o��2�W�\+	X�ܼ�Z����'�p���1J7=��Qk���j���r�;,����-0ɫg�I�Vg�I�X2��SK��PJfت�b�e�Ӳe���M9��MC�@�\r<Pj�=<T�|��_$o��i������0��r�K��C��b�^&S6ⶥ %zZ�?f�_P�nxM��CĠ�#�.�)���biD�qy�Rv=���1fp�U�A�k�K�ڤ|���1�	G\�Q��L�GԪ:s��/u�����V ���b�k��Ş�!	���^{��R�� �zT��(���ӑ/M���8�� �Jً��y
Bg5<�S�<��F����V{��C%�����5�-0Q��m$Y����K+{$��	B�am��8��1 ��ƅ��
���:{��ݐ��Р�_��2*���g�@3B�8������s?��+��3���E�v�|.��uL�_�B|�x�{������-_�pׯ]w��/Tb���.���{��51!䀡5nz;����t��:�g��J�����_�6��2P� ፉ�rN�̤\"�:<�D���Ӕ�7nxu��Q�]*ÝPå���{-��%V�FM�L��6��I^(M��Z�\x�`�]�HY�Pb�0�D�+���s{�>Y!�V��)��@oѰ��6�G��p��2f�)��nH�T�F�$�/�U,��^8A�u���2�.���/����RK'DZ��6k�R��b%��H��J�ė�L��%��d4'ԜP*��8�� `��#�K��%q����R�[�n+�E��YU���_��;���j}x���R��������ۻ�Y�������o���.{�5G�����	���O
���}eSɵ6'��=�!�������Z�7�clXO�~��j�,��8�������e�:H��Zє�0�,�ݨ�MC��(2A�J�L�7Z$��[/�M�4��B�(�]3\�q��٠�ɝ��ɨT�؊�)����o��^�Q=�h蒛���{�-γg�� �^�@h�����m� ZJR k�L�Xk��¶�"s�i�i����lXP�x+����d��,5׽Q��L�.]r�O�!� �=�=�"�J
����[+�U����䗂�6��2�gE!��c?p?8kXc�D��Z;TZU��l��wʻ����2?�*�B�Ą�f(�����f�cM�J,�aާ4����g*�7����|!5H�=�S�٠��$� ��������2��Ȱ��R,�Uj�l�HWO�0d� H����P� �=�X��DЦ�S��`L�����!�Gլ��Qa��8��sB~�z>�$���P�:�Eѽ�h$kL��D�զ#�ZB��]@�P�u{�]bo5%�ji�Eǽ��%ޙ���p{q(%I���@Z�B�'")�t�	����o�T$�B~:>���rP6H��r$U��d����=�e�07��u$���� _ `��8�"�R0�X������~��y�.���3�%�E���l��P�2G�3� �`��ba�-6����ܻ.!�h��yϜ�Q�� �\&�"8+�A�D��j�g�J޼f����|��W�7��
Q���j���>�����<(Z�ˢ�VgmRѕC�y���іW�<;�ؽ�!#�KV�Ŗ��	S���]Κ�]&���A�q��F��l�� �@x�Z�� L�C��'�I�AKmm{�ILDs��ذ�Ų��mH�-���6�䩀ȱذ��B>�<$Q>�ű�;��$4�Q˒�#E��-�%� �o�霐E(	�������/&�j�Y� �?~�;q� +8�˪B�ˎ����9[�/b��þvE�%zP�EB	���eqݴW�_�����X�q��-����`�1�)X.(T�XyX�h���/2�KK�(�pE��*�� >�rO�ch$+,�aYxĭ�W���Q L��l��zNi���l<&l�¿ţ���7�U�o$�pw���C�`�F�i�:�ޠ��r��9
0&r�t������Ub�X+`�![{,I��zr%�����d\�Vkf LeLͱ!M��M��Mv,$���kS&�TO�]�l0Υ$!.=��Mc�u�X�iȑ&(p.^|ɽ��;�v<�p뽕�b���q�px_��8�8(�p�x�w/���;i0J�E��q�pzt�����A��ټ�:�<�^��ɓ��tBx�/"�؍%9	��
����3��;�pc?�Dj�����[*[�Z��>i����=wڽt�%��o�f�I8٤����4�ī��%������:y�+u*��m���&�wx��>d֞�S'O{wsM���F�=<���ۿe�G��ݹs�Y� �ԩ;��������]�g������w_�����@
�ڴB�-�T4\��_�c����}�����,��=솮���m�8/�4g�J�Mà�|$�1�^p������ݝ[wXGN�ݘ�~Ç/p�Q�F�郕�5�)��2.���4ft$��?��%�Ff�1e����5D`��7!�d�S�ix��sZSl����J�ROR>��-�p�1&�{���o9 �A���ASw	�Br��-����g����:���)(ĸheX{��N㱶ė��}f:����#���[a��ԿG%����0)��_H_�?��a�G�LKy�5�.�$��X�ҁ1���[�7��r���߬y�R7V8�����	��a�JP�N�|e�3[��Z__�k�EEd.���Z���OЃ��ͮտ��Q��#���cO�o���}J@ǲW({�[�rV}�z��0[�B�swY^+�7��q�:������g�Z�j	"�\�9�pR�0�u�>짅w!/`�FR�Җ�.2�e�I�^f���b��a$ʬ�C&-[�4^V���'m�z:K)Z�Zk��V���K��k�P	{gL��5�,h�5� ^魭�w�w���%�#��`���So՟&�̒X�"��PP��F�ȣ�$X/d'MSZ�������l1���)M��t%�Y)g�Z���>�Z]�����[�M����yb<�;�����71&����~\��� 
'��@x-,LQq���ys�I��s�Xr᠊"C&�]�L���7����J�����ʒ.1>o�;�� (�^���ϟ�9>[�õC>^A�[�.����Iw��i��&�����-c��W�@`�<�N�\�u
m��g�%�\�h�
r��f����>��1N�O�ҭח�|_ej��U��cB�(�Xh�Za0Uk���]��N��N�9�UJS�]�E�PjV8�`�����PY"Cܘ~8�fʜ�3��ŖC$Vur�L!��N����n.�!�p��B�p�6��b��Jdq��1nn2ڸ��	_�,������#\TPeظ�nbpy��/5₣~����!�ݑD>'�K�sM���#x�@��������,�L�8ho�d45�Yq�nWȚg%=X<����_�����O�;L5�*b"Ur�Tb���2�=�9'����C���(X�� nԽ�(Xbd�m��k������iv<!$:�wS����V}�%�BQe ҉����֛7or�qF���3|^�u�&�k,Jc�끰 � ��b
(���K�ǔ)��B	�lj��3M��H������L�;b( �P�6+.�#�}�1ь3\}���5�.rY�,,��1?�B�����عcYjR��KI�EU��2uq���Mh>�@��{�$ ��� )�����21�t���y�+
1��o��w��,�x�Ɇ��{\�r�xZ$t���G�lp�!���R��6�&������+��{^�z���p�:m�X/{8?��>|�&'��O����{��GﺕU� n4b�)e�Pc��ws[�sn��S�;{�.(�p?ӊ�"-����t���Ҋw�ߪǄ�M�|nܸF�z��Iw��=�;v�p��������ME�7��y��)Z|$G��"`k�����wm�!&&Ƙ�1�UH���Ӽ��E������*0̠�Ւ��C�£:�{뭷x��@�b������>��ł3�p
�J%W�T*���\{��:���j��ȡ.�r��ӱ<2����`��:#Kqq��(��nuhA+��M��Sm5g<����0?Hޯ���"���Z�>BA+M���͋�̽�?���o~�ڽM��O~̙�}���{����S'u�%z��^�w�}7�xF�����W��<�P�k�/l2bNh}#RL
r�VH�*c"�B�+,\DP��!�.�qP����Vknq~�P��K� �>}�[w��y�����1�a��9�ԅkg�;>���c�\��r��N�˗.�v�5�rb�d
u��EL�������/=�&�2]B@���p�B���Vp��� k��~��+T&�ﾻO2���Y*:�_�z��SB#�ܹs�F�x��
�\�ݶ��=��~m�&�J�����}��ǳ�>�l�'���/������b����j*�7r�#��y��E ��Cg�u����S�v�>�ʆv�\0�u�%��G��
���4�2� ��hb�u�6��Y�i�n����4Ie�����"{�Y;���5�*%#�pΞ;â<�4,%���Hr�=z��H��ai�6�^]tL��W��!�a{�7�����,�euN�YqXX$Q>3�5�����P��$��3�?�����x��|����)��|������Ϲ�y�x�u2������-����f�K��pe�����~%5o��ĕ�~��f�{��󠌥%�bḺ?��+�eلJ� ��M#	t�u63
�����7�|#�[-^!�9��>!��D��/zݠlk�E���Y��ɋ|���F.6>g{����qv��8�??�$۪����j����)��\=4�K�F��BW��#ǁ���mA�E�"eC����L��5��/�(��M킰��L�R�*JT��C��I��ސ̢�"��k��D���Y�yn�!M�Y���]��vA��XH���!�6KXAc9��-�,�a���z�*Q]V���F��0��|,ۍ[	��/�� d5�:6�X!������I���������̚��R�e��M����B�'|��v�~���|8�#r�m�(��&�
3� z��*�ibO �FP�	L�@ڽ[�gC���������EZ�����ޛ?�q]�7�����h,�XI�$J�Ko#YV�?��?�<c{&b^��챤�dI$�{c�k�̹���s3��R-���h6���*��{��|�A�I9*�����G�ë���kA�䬶e5bC��'Yzr��dD�`#�X���^�������șG�j��h��S_��m�9�� �`*J9R>��j����!b-�چ�2<!d��(f��{�lC����W]����eu�=jC�%���|=�3��!�I3�A��dy�JYp���BK�S�� �d��zXG�����[�}��׎�}�D���wX�CV�2/�����F�778"�&l(b�^��#�o�6eXl34<,?����k���MC�ԍӔ}�����z ���e����}����:�;�5�se�w�fH�GN�X��mԇ�1���� �,B�kTvh�Y�66w�L/���_�%�0�FKA5�!W�)u�5���_�h��Cf|��G��м�9(T(�"��G7�Lx��%�j���}cM�������	��n���-
.blX���K���s�@��ʽ��Ïi�Q��p�ce�=!	w�04:"ԀA��<�E���GW�G|H��H�|Դ���3d�6?��[V^B��']V�{u��6�9X�e��/�X���[cs*1�Z2�,�<����y0�7�T͌�*ig�\���V9O�����v�h�ܙ����Q-u�Ҩ��P�ʸl�2�6�����e��h�"�:,�<��S	(Z��itA(��o�ܧ�1F�r0���э�f�2�%]S������5���q���Q�H�՟�Tƪm-�f6!�'�s��:�R�L61��8����݆��w����/Ƹsa1,^�J�A����VN�ڟ��,Zе��x+<]���j���TĔ��QId	�L��#��ɶ��.��D&�c3�Z9z�H�8������v�յ�p/Z�����߾O$(~���x�a=�w��������킕�b�<¬+Z�~�1��O>	���s����{�)�H�}~�v�Xʽ����b����!����w~�l����cZ�����D�=YWΨ�W��O3��R�=�] 2��B��-�R��{��,#�1B���@FR�B,(`�)�e�1^SY���T �*��lbr�R�WM�f����,$�ʭ�'��Y�:=�X+�e-���=��#�ds��Ɛ	��ĉc���9Т(���4-�\p��
B�U�ſ~���g��\=����飰�$(!\u � �������v��õ��#��P-Yԭe����h2'���C
>�M�02Ǐ��hZ4�u��b��n���ec���r�F�t�m��x=ܼ}?	B���cQ����gӎ�G#&̌kL-~!e&�|�o��Z��߷Z=XRqM�#VnO��X��-�����.P�"1���Lk�,���>c=���W���u�y����9���"��`$� �<���qgO��,�e<C��	�d�;K$���B �E���k�RT��$�.^|)��BXZ^���\@[�#�4���tT��vWrj�eڲ뵁NXq2��<k4{+�T�ﱹ*j���Ü�B�Aɯ�ޘ ��jo������׶�a�}�2�;%��yfU?*��󠑯'O��&�Ā�@܌�ݻ��z�'�=j�+SF׆Ì�d��1W��6���=�>�
�֚�����/�fV�j��,rNa�� �~���%|��Kt)���ޱ,�����'�w��}�õE�	�m(2XV��bf�9�@;[=������F���Y*(թ;	���wX%2R�� �?V�_�nfV��a���ٳ�ⵞ0 FHc`𵹾�����k��b3�I�7do�9�K	K��d�(\�7����}eN 1||(w���?'��}Kf9�/( ��l�cћ�N��L7>�	��8�g
������PZSh���Ċ�E��9��-X�P5o}kN�U�ެ'��G�&e�`G�5�O�[�6޹7��ɡ�����;uS���%tۢ%)��o�M����ؔ{woqj$@�8���k���C�%�� ,/E��F(o;�5�]]Z� �Ze63�b��#����cЌ�ϖ��P>nj�*g$yѺ9��e��2�;-x��3�8��Mr~�\�,�Z���<�`�(�Ȯ١�.�	XA��Ë^;��]lz`v0!�}$�_���B������)Dp�;�tP�tf^�`W,���X[0�G���X�jk������=ai�nP�P6���J��#M�`�ʔr��h]S=zhM7�AG���H�}	P�=AAC�|��q ��0��1�相�\-�����(�,k��R��I��$�;I`���	�KE�=�!ջ�����cO
b3A� ��W=S�'�R�������B[���lgU��?é��;t��v|9�
P�x����Dh��
�M�㔡D~'Z�^�vŎ�pm`	G�ҽ���,��=Q�A|�e0\/��(�����:�����ޡd���A���󬕍571 �m�0C"� �2�a�Q
j�F�a����c
�P��-�<hf�������)��Ail�����Ef��u)��gm��7�Ȧo��ZB���&r�*t�l6=�U�U�]��
�У�ؐ2�����{�6H<FV�'��N:�,5r���S��P�B{h�ģ�ts�m�g�	�����v�Ɇ犳�I���n��I�Nn>��	�<׺a���<�mk��n�<(N�h�G�����5I�� {0�7[��b.ƱX��{��Gf���9��\;b�͍-��%Xw_dw�i��P����3�:�!k֗�F(,�[�f�ęHM�$.�aG��H�'���'�>�=Х5G�4#T���R��Ѽ�2��Gґ ˉ���'�F3A��cfp�����+�0�F��[�'P�a����U�̂M�\�^�*�o�'�s;N8KM�Ž��|���V�u~�����Vs	b`ZF�e��R��{yY��$�~����q][I��_�l[��+T�Q6��=�6}�!d�hU	Lgo����S��>ȕH�h��C_;�f^�i,p[~�}��������:T��J���PB�}2�����/����-��p�lB���[+aݑ����5�,��B��쀇m[�[i�3<��x�
yZ3�7��z��N���Q{�Z@�3\;�K�C'���Yj�I���76ُ���:�����s�,-~�2Z����-�W�Za>�!j��B�Kw"����S7��>���1�V��'_o�5(p�L�g��൐LV���k堋�x�����a��
�vZT�6Ci��JJ���0���|O��pD]a�8��R6�Nt��\S�V�u*s�d3T�A�7z�9M�̍!�2Ɨ�<�jB�P�����,�XSÖP;��L�����6r����n�b����`u�୊C&�@����:�4f�*�(NT��2��Y#��UHt����m��>c��d���F��k��Y��,�è>Y&m�4<�y�C��@��ņ ���ʚ�5mh�]��6[���5�F�Z�]NtPf58�%�zL+H�D��om��R����ښϓ��&�_O����6��u�����B^���F)�>`c���Y���V����JC���c(��<��}θ�>f����'Z�I� !��<���$N�yp6�%<Chځ��6�m]�#)'d$4ɯ�e�=�V�rJ��6�T�R2�) o����ywm9,���F��1�_K�������J"�'K��~������3��Uz����b�ug�����Y�m<��f��9Ņ�(���͎�р i��"����_Ԅ���^�ؕɼ{�TB6wl���R�w&����
/�@��Bܵ�˲`��k�YY�f"��;F��1¢t��A��<�v����G����Ie$�Ng�w���s��ׇ��H���8:.�ʭ_e��6�Gh�Y
O�@'ݲ{�l1S��tO>u�����
����������vީje\��rM+��d�%����[��_!����!���sW���a�{�Lf��:�M��Ջy�R�0UJ|��싧��?l	���u�.k6S����h6���"�bAl����tH�U`���H�d�`��Ln`Jevk����j�Onxy!�/�Dc��h��P X8�4�C5�&������]�t�;�$���a(2�x��W�{�=��+'+��g���������$7���CU`2�RMXgO�|R���Z�`�Ba��I���+�%�]Ҭ�YȚ��Ь��5O��v����)��������[Z\
�����J	����V�ť�P�f8���{�#0䄦��6+yR�۲vK7BRz��}�]�&*>�Kg�rr�U����
��ܖQ�u�v{a�C'b`�����>!o.�Y��d���Ș�m�$Ԟ�ͭ�^3�.%Kb\}�!��>sB;<�igG�V�P#F�k�j���L�u��N,E:@c�/w�b5�ض.<|f��J�/�4��̕�w����nf;�6\|.�Y����2����w������$ȀiN0^tZ���i�K���4Z	�.d��޽�<�c�2�$�����~k3��q�{�F�Т���n0ϴ4E�BB��������Y��,>��F�2��o�Ν=��t�G`����Տ�[�#g�Q����������x�i�Lf�|�;!�_�[�F�B:K-�aҐ��-�n�t=>w*�&��Ml�L��de=�Aܒ���%k+���vdY�88�v7��<e��asx%�\⒥�W^�~���9�Ј�!��2�B�t`�4�<"����uu����2T��	���$I%+;8N^���ˬ�� ��J�T�a�q��"���$?Ϝ�x���N��lc}�C�����ca~)�1po �@0�PpPIF���'�p�F�nC�{OZO��v�����S���@"ID|�|oG�,�f-�\�U��2���c�ҵ���yj,�' ���B[U���v�׈�
�W^	W^����sX�˗/���
��2���ǎ����r\N����-�s��rs�~����88��"h�D�|W5��МK�S}������p���B�IM������m�!�z��`����IK��.�]�ҋ���\���S$@w�3tb���[c��Үp�-��Vso8���εY�2�Vwlq�3�6�x�W�����G) oDHQ��@B� ��L�S�d�(���_{5|;
(wg1Y#z)��x���G�4��'?�	�կ^~�}燢"��;�	?����:���?#q����O���B<�/s��ڃ���n��S����K=��M�����](�nєkK����]&HsF��H�˦��]^�Ļ𒞨�al��u���3B��l\+���51�.�H70z���Q��0�"��R� ��)g.��[� �e�Ck�������������TVt9ɲ��j*�6W{Q�Xr �U��f��6�(�P��-�+� �o��M�����R�o�r�(p9jX|���ø��B��D�,7��՗%������ny���L3�5��wq�JzI(*;���H�T6X0oe+9����E���P �1�^g	�5�c>|0�I)�E�(�1D9���8;��O��F�%��l�n�=��C����H�:�JrW�/g��6�q̿��0O(�ZdZ�L.���.�ܙJ1v6�M��-�&�э��\*7MNv!/w\_��:~��	�<k�{��;w�ӳKC#;;�ֈ�ɛ�&]8��OB;7u=)�ӏ$�s�T�0�
G�c���C���kk>�AS�UڧΛ����6�H�A�ߏ?�6ꄴ�n�՞f_��|Q�b�`w'<X���fXZ\P�(d�&�а�[ocT�h`1�(���}֖������O��T���]�4���.���9Ѻ�N.�=��"Ňͨ��>:�B�ܢ���-�?\{Ȥ��Ø������aꘄ�~+Z ��3�b] �y��a�5�j��1YU|j$�qj�� l�R	�f4�Cf�Ҍ���1�.�a�n)Z��!x����z�x��s��A9Գx��/���g���ݮ�2�<�� a��T�}Zpx)�V;�@��[|-��I���������&�ʓ�<�oġ5}j-����kM��u��WQ�!i7	b�L�n��2��V�9�ڲܙ��g#Ƈ��{�Z�c�D�F�C�����VI�#��@+���զ`�f`�%�`mn��;�����=��c	p���؅Xh�fN����C�vm�%!n-���Uhj\^vK_���x�瘼QS�j�(uA��V⊗@��o��xe�vI�q>�OÓ'�oa�ָ��T��OLI_?�9zZW,1�� >w����i�������M�*%�:y�&j�-�yaI*��;V�2]G�\d%x�@Y��8	�����@x<]J�=��9�(�n�G���1S.��Q���l�I�����_�}�{���jgB��}ֵn��S)p��U�m�W�����"���󭘚�5b�q�'��
���8�8��.��m�,_��CSD�E�kC�sƽ���mgF�x�)�\4���D�c���o�̨�s�R���9��(u�ĵ�q��!F���Ѻ���M[�)�s�9�=~@����==w8
�okc�n�؀��kk���v����b �g,��(��w3�Rm�3�TC�~��ŰߟL&�E� |��G)�ƚS �:-wpK]���X����ם��_��	�m����3`�s��PʱB���ߤ:=)����/9�ݽǳ��D/5�� ��,����O������D�����?����~�Íʗy�t0������j!�Z,(F�Om�1���nR��[h�F>S*�M:�Ȁs�lB��$/���a¡D�+�.���wj��C*vb��d�@���M��9�'��ypͰ���h�X��&�_�X�q*��`oA�p�*�Y��9Z�O0�y-w�D@���Z<���bj&�	?6 �}0:�p�Ȃߍ�:�eeݐ�ǵ�<����� ��z��ۚ��/��;�T���u��%�[?��:��k��f%

,#�	���P	`��ںJ��s�Α��~��y�z���.0���ψC�?����H$$q~\yC=�Vkw�ҥ���p����ʕ�d]�yB��/~�����I���*N;)7vmYhɘ�_5�M�ǉ�0�����3��n��V�������l�7�#��=�t{y�q��%����	z��C����,{W�A�;��� q*�+3�ڵ�j�,l �z�|jF��Z��ABC�;P���Νe'�� p��Yz�
�N \[C�;����U�kڰ��01AZ�w�&0s�f�j� wY{F�9�c1�_�~al��	}���{���xv`D�
"��7$}���>ۛ$���[�/�B�d��ZB�XK��O5���I׾���� 5r4����R������T(���7I�? ƀ��VOFC��S�˗�'h� f?dj�T��z�+K$������W%�
բ�bv�˶=�W/_	��"
o��?�{�߹�G>� l �T�V����/�i���j���\��{�]݂ ����"��u�䔡�@��*^WeV�)��'$e�z���*�d�y��@B�Q��m!��p�߸��z�M�:��ƍ���z�|�N��N�.P���C`�l\�+��ʱ3 �[s�6w�y"�ͭ�p=Zם�>|���3[/r9_���稔Rx��Ax����~H�v�ԙ���0�8y,>z8Z�5���.4_DO��l& Ԕ�-)����9$�@whnA�?���<z��݈�!".D �=�}���$y8�|�?�U��
�։�2K�Peu�Y`�(��k��v��>�O������8t(���׺`
���=�r�g�c_���U��md�A�{��r�-�'�P|�Z4u��!_��A�eP��2"��@�� �s�B�#z�܍\�"4H;&�̵w�)�}@��E��?�A!b|�ڃ5&�F�*<���
p|�K�	�x���!��`dр9x?��OɊ�C��k����?`O?�8T��W���M���Y$=3�~��/$i1Ø��&1	N��t�<�u�n{�MR�i�X��Ċ�	��g%�|"W���E��{��z��_oB�Y� ��`�D���AԒ8X(� 3�~h����5Z�^?T ���	vMǽ]1��!���⫪Z�M#����s-3	�=��	���':�'�i_|d<6��c��p��Ȯ��V�(����fD+�a��q�ӽS!��w���0��%�x�,b�C�R#la�R(�D�8��)�6(���+Q�['ܐXpu��R�`��P*�_P��@��k4�g�p�K%�#I�vi]�PRR�a�s��?�&bf���8�̩�}:�F��8�H-���ep��*��V�����{�WC�h����[Y#�P܍k/Pd�a�����*�ҳ����Մ�d�wY���Y��ŗM2Y-�բ=T��t\�.�-ǽ�[�/s頯�H2%���ژkv,�F�`DV�������.��Ơ�zqA,([Ff0��z����,���<88���j�NOe���D�>k/�dⰉ��<�LU�zl���|'��  �a��`����`�ӌQ��\��.�:׆kD��?������>�:��*^p�j-�׸����(�G�ύ�8z�����ر�8����̞Q P?�r4x�R|䃴V�=�۴��:�?Coy$� ��)5�ӓ{K�oME�\���#�̷[o/��xPr�.�u1�B��E/�	��3��ߺ�y��7ތ!؉��U��g7>��e�q9zr���S���|��J�,�Pa׸3N�u�J;U)Q6)լ]���Z���ɵ,�M�)-�	�.�<+���V�;4j������� ߜL>>?���t��=��F����q\<�nݰz�a}��M���s������O�{�'��+�@�D����|�����aW���4����S-:��L)��Ą3�h�^���$F1v����M�����.��@�a��}�=��F�	*��`�B&P���saa�w��\�˲�y��!����B��T#Q/�<�e�v�>?�ʕ��+�\Q����YCc�@��]q���{��Iz����{�������׺b9Ȱ�u=qp|��#5 �#�R�F�h�szuO?&xj��|X=�N;��	z���Uܽy+�mKpW	G���,<A�K�;�q�\V&�KJR�V�����Xyҍn�z=y�4��^-�~��l�������U� ?-�	��ú��̷~9�\����)�/z�+iIaY//���Ά^1��qx�v7�6�_1<.^|!�;{��Z��Ml؋����Z���~8�r��?$v � �r0�\;;j��Q�etC_Uv�S�R@�SAvP�e̻:��G���a�K	5$��n�8��l�3v��2'f�2�����q�5���nѽE��ptˁ�k�l���du��戄��GO�]"ɔ�
��h9�N��5;�+��G��B�q*�/�.���(��ܻs��4�S�Ԑvxx0)�,K؅���$�=ݣ�Rh��	u4v.v<��#f�;�zC8K��!y����s���Vz��	a�w��$~����|�bm�M�/v$+����s�������,�$��_ӷ=��v9�G��nM���O�g���T���-��%�h�'�sj�V��(�;�b��,�S����Ù�f��:;�]ܸ��uJ�;rx1��ⅰ�w�����~_Il
^W�<dh�D�
���	��L���QU�D���'R�2�G:uz5\�x���Ç�Du�\���\tm�1���2r �Ȕ#s~��5�ݙ�BÍe��u�v��y�������"�RP{im�T8�Ŀ��B+2�ͤ�<����cas'̡�c}&��-�<����o���#�u�7\�T��!�[�֖*a��wg?[{��9!k�Pp�QA��w��T!� ��N��hi�7A��`�Z9���3�/^8/��L#t������҃j��=���0�b$׻����27:�&��G�R�䜂�������Z��y�x�;��L43��N.(����!e�kiTO�{l�H�oj�n��l�l7)~�X��76�1(�G��B�y8�RKW.s���(Ĉ�K���\��/+>3FK�ڕ��������	X(�Ƙ\����\kj��������n$te�k�1�p�sI��=gqq�b�<��w�H�Ԋ�#x�.��UҜ��u����z�;��|��I�ƛDB�@�j�	Y^`�I˔k�wy�
O�C8�)��q��]���#@}!�����JwB�yH �Ĳb~աw�f'����-��l3���kQS�$�-S�-L~��u�
$\�Wp�%�%^l�wh~��T����Y��^}�n�^no턭(�H2B�a�_T�H�"\�Pg�4�n�;������_�x7��xF��ny"YfM��jB��@{�
���`�>Мo�ο��&�>%K�|t'"�_�Ԏ��w;��'#]8x�kTۉ��acfW� J��(;Դ�����JrZ��ñ%Q�����M���Ưxo���Qs�n[p=���WOұzǻ�<I%0���fVM%�尝Z+�C(.�2lm�3�s�������������&kL�B{us��\n \�oP<�1�֦2���N|hv�k��]�=j�wn�
kk�H��.���z+���^T�%韺�X��_�E+��x/]�;Sm_��+4�)N��0�^Ի�K�S��j,WSQ���)�Vǆ'�{̸0R���� ��։VZ�"�����,3�C����u�z�P��ઉ)�,Sf���c�̅�__���V�2�<�M�<�yDes�:��&J��H�q B��$D�A�B#���&���څ�cr�������x�eWbvL��d]!��x80R��13��U��$�inan �* 1d���fc<~$
0b�KN��$��uk���J�q�ݢ{�6�Q�)����*8,T�	���֜���:
����߾��7�N(�W�����$�E��K`I�]Lq��Zn���I���{�l�Dy<��p:n�.v�^e|�f(�a�2�x��$�� b�W7M��p�6
�%j���R��C3_�v��<���3�y�)��^�����<>s)����%V�mdm��ҵyئ�Ċ���X���@�ʪ*�Y��ܫ��f㽼��o����V����L�32(�v/@� �2�Q�M��p*Iդ�j�Zl���S���퓡��[�D9� �d���>vɄ�$H����O�L4*5�^d�>�R�J��68\��}�k�;�~���paa���42��ÌW��b�����X"��5�q<��Z����K���>	�޸IW~�6V��q�:]�b�:�P7��e��x-�0XO�|�ˉg�(	�/I��^��߾����i�u붱��wA��d��Y/�f\�U3XAD	�ΛPc�m��ϡ��a��^�-�vC��u�5].I%jZ/fE�T�bn$��|�k�~
t�Rbi�W^G%!�&	)�� ��ͯ�ξp6ug��)��1\��5���R��1t/u��Yk�j\0��Z�6Ǯ`�ћ���J�N"��w�p�P4�=a�z�xsq��Z���ͬ�5���dp�ch����%�F���S˧:"qּY�eq:9�x(B(�Z4�Yk��
^*ԕ��z�,n,��&qb�じ+4�5hṰҔ�(|]� pP �q?�B���J�t��N����DH<'A�4'�=��JO�i��4��P��K?�n޾ǘ}gw΍G�%{L��k�dA� $JNnQ�vR�H�19�6�R�P�kXep�*_+��%D8`q+��P��6��%�E,����if|+�.�=��j�7ͮ���7��N����XM��f���sgyV�\�ƥ�{�<��l�lTӓ�f^1��p�ޭ�z����Y��Ҹ{T�GLlvm��p{M����!��h,��m�ʱ�3��p]5��E�G%o0�b��;r+?�����=1�$�fV?oru��y�g���y���a$�N,��h�t�s7ӏ6@��!���\'rk������pa��B�Z�S��䡖�5�%���J�@�0<M��� +�ϙ�,u8
������J�#�( W��s�"B�j�+F�p;M��ށ���Sý��aR�:6ݛ�c��׶��\���`d��-Ȥ֭X��2[��:��ʸ�'�cC�١ۮ�a�q�z����&���G�G��L���D���KvbM��9d���_���S�1�Vۥ��BдGv��s����rG��I���E�)�)�����X�ʫ0ȁ�>*�w�y�}��\($aBj�`��Kcs%	<�Rk	�fa?�F\酹���W"A�Jw3i�O͙_�ssb7�\<w�E`�E�Z7���QP����Q9���([�I�8��Ɗ;'Yeʎ�n��l���,��S��	���-�	�
M+ܗ�,d�L����!�q��a��t��wwG�۵���}�!D���� �FM���=6�?N�r���p�;(j@06��̋��7���,��gbj��K�D �X�(���X. �uL1c�=�ݼ�%�Y�uy�BS^� ��%#�#0����y'O���sǏc��1�i�k�+e�wE�@M����.�ei��!���A��z}C|8��xy+��*��e�&�P�C�"\�]�(��[�/E�����d��7��nF��z�-�w�Ñ���0b�͖Yh``�3�`�n�x�0[|��a���R��SRiV}˚�����[��'�R���Ƞؒ�n>� +|D\d:_���1&��yZ�g=ڵ�b�Um�H��C�XD���ΐ���N����[��mK;�Ⱥ"��9Tq;��:*�ԕ �/���A*k�C!h[�}z=Z��9���'e�+�sǎ=	�^�cB��^_ 		r'���z��Ҕ#~�5@��]�r�����W p�0?
�MN,���*�����̠f�uouR�?E/�뒒M���-��5gs��\�W�7Ο?.\8�z�qO�*� -�a��iU�,�ʑ��C����-BT���ؗ�"�,T�1أ^:2��JM��� ��z:�X3L-��U�W.�$�MH0�n(k��
EV��h}p-�KD�����A"kS�ZÃ�}���%���݊�41hHj����/�7c\�C7���,��w�MO̵[BK^��=.����ܫ98�~��B���5Q�'�TzR:O�,1�c�%���h����ζ9�Ri��Un��K��AL��aqy�.I'�!Ǆn��Q�>����o�l}��'C��B.&c����������nE�����y(dƶ�lmT6[Q�Gw0��I�N�p�4��cϠ2N	2���LPm��9��BהO`������*8�}e(��F�Yd�lX�<OIͷ2���Ɏr|l���θ�D�#^��<T	��T.1�Cw=�]Z� �jOɜx��@	hef1!/����ʖ8Օ�lZ��J0̴Ӎ��^q&0�>a¹�Э�s���	��� & �)�N��:{���+WY)�H+:])�xa[�=���ppfnV�6�e�-������܈�{y�3a����K�6�gh�}ג��*(Q����x��'����g�ܽ ��(Đ?����y�����/�g�w�j�A�<-�:�v����t/�8j
�.��u��]�p1Z�W���Y�.���ID�r�p�,J[h�{G�yUNE��*3�@�-�����|���s�3��
�AI�\|�\T4�a?�ݰv�!C*�ȗAB�� �N����֨���� ���\��
��8\Xl��b��4��gn�ohoK���{b�����I��kM�Y�¡�ƐK��k������#鎤�51x�H�\(,\��uX��h�����������h��*���"u���[r!��˚B՟����eC�-���]��/�O��������õO�q��4����B�ww��ځ@��#,ڌ�ށ��L��_�t�E�/�}�a��>�� Ρ&�a<�'N��rҽnU�R��Iǋ/D���9��}N<'���'��7�8�=���@i}=S�j]~����b�(�j4O�Px@���}"�o�F����^c?2�*㡼 ȃ��-"b�B�о (�y�vx���F���I.h�)�����UF����L%/����"��=�j���e0�tf��@k��ot��hXbv��eqBy��,I ���v��.�o}�������',2J(���)�,���-���&U�m����݄;�������Ȓ+�hYv2ml]QNz�����R<d�5� �5;�Me�*�s��G�OO�N�3́%th�k��-�ڳ�52���Ę���P%m���2\A*�>������s�kd`���j3(Rۜ�]j8�W#Ξ. ��GA���r�E+\��|o1lo<	��1:-m��<�+�I��xl]�QqM�-��;���/^P� "��5�Z����H�L��ʺCq��-ا_D�x#��v|]|r���G�&+w*G�AsAX��Ξ	���?b��zX���9��wl�Q���"+�x���	����$2<�8qsz}PɌY��ug(����?"����L��k��c= X#����b�5��C+����T���{륗.�����#9�{��A���k���݈�-*k��g�:+�q�cGbu(Y7�R9��L�p���1���s��nC7��6qV��VV4�Z+Cj1�s����V���~�1'mp&pP�w�9+��*/*�Oe& � X�7�x-
����g��szSH���I����Yj#���'��� *��+�6WY�*7^���EH��?bʊe��A��f�#����~<3;����G�6�ݵ��>v�� #, �� ?z�[ok�D�[e�*�#�,wAh��>��p&��3F�����S}�x������v��@�ƹb3H��1�#�����%Ν�\y1�x�"I�x j�ix霱�ZҚ� I�l�5^7ݼN�a�ɱ�wn�G }�X:##{o�A��Et��=�a�/Ʋ� ��Z�w �Ϣf�|�N��(�����q��\4EV�vh�@{���p�S��8|t�3��ww���K�dT�����G6���>�fYǇ:��t4JM���8I�Ռ5�X�ܐy�Y��r{;�Rץ�hOr�����W;3�U�.촪�35�TF��	cL%K
��e����&''�a���sN�D����#�ҋ/�2i�����\x���)h��c�H�Q~��;dLy!Z= � YŇ�ܯ�׮�31`;�!i�,�ٺO֘�G�@,�7��=����d�E��Y	4��̎��e0�G�C�PXR<fz=�+��d���^5���W��cG-�h$g���������ћޭ��cѨ���ayq����l�G�H0�Y�����VN���4��\���c��-Fk��r8
Eݧ��Ƚ�(�F[[�8]�j���i�Qvz��Kѵ�-ߧl�hs'��UYϭC'�K�⚊B6� ��u'������8�J�j�!�( ��Y�Q������=d}`���As�X��R��<]V�T�>�����ht���.�-d�u�m�[�%+grm�'�^��Q'圷ZY�Ř�ܯ&��<�Jb|"����y���0�NS]�잕�	G�'Z�3�0���`o;��p���𝷿��W��m�Z�ތ�U�}D����V
�d�*�c�O�īģ��T�d⫓3a���ذ¥ʄ$�(:�"�$GEC��aB��̇tr�4,�0vp�U!�F�3.�x1zs�E�����b4�!~��M��s�ڳr,�R
���Gi��\~9��L��ZƋ|m�����\�T;�聥�9�G�F� xt5P�I�� :�M�EȲ�p��R�>u:|�;�!�6X�(�Y�j�6wT�es[D@Km�ol9���.�~�1Xպ4�����W�E�Ś��W���p7." �Y˯}�k̨#�������l/\<��c�CX<4c��ǦU��RP^��u�MiX��dO�\�yL�v����k�Ul�w�A�w���*t4�Nw*(hH���Et��
q1z�O������.�o�{"��"%!=,T�u��R�cb-Z�QT�3s3�cP?ǽ�{,Dn�	��i�L�W�`�@��Z_DJ��\k.zƏ��?,=,8�n�;c�Z�������#>qc�e��S��%�x�GR�ƍ�X�B)%H3�:�����Tk,� ��Y���d�|w��w�tE���sa)Y�ך����Ģ��W^	7?��>��]G�X
�)}:�x����҉+�@���b�ᠶ���E�����������W_�����<4c㸹��/]b��/�A=���H4;`s�	L����kJ}����iͬ�ޮ֑am��g	�b����韧��'���Q�E�\�P���qd�Q�1`��s�֭���RϽ�����/�����^o���VC�N��S#�E���c�&ǂ��{	����"q�Ѣ;�P���l�dL�N.us�����J0c˥�	�m���p�F�<���R�Ԕ3�O�̅ک�6�FbB�1�uN{閝�jzŨ]8�e>P.�������t9�pnmw/F�8X$`x_8�j�nyZ��/�n�g4]C��/9��I	$� (���X4;��䩹`=C�Lr��& �l%>�ZboĀ��
�S�b��X�,�S�7�Z#3C����bk�[�6������L��:�	�Z�N?�ǅ����/\uGi�L�������x"Ŭ�4p�iK�k훚��	v;Y6)�	v�GՄ-����H�������^m�ڡr�B���K
!�P�H /p�����S����Ԅ�U�&@&�r">Y��~�;a%ƛ`>ʯT���Ld�[�:��]6f�%-:����	 �Z�����M�����vkXb�v	e/@K/^����s۱9��$�Y�ֿ3����C��<;$z1���>�.��D����4mp�+�[������H��"\����d�`	�@'��~�5Ԥ�(�ϔy���*X���zU��
���1�W�`�֑�x�j��v[�_�P�X}�2W��y��$������Q�C��ر1���H���CN��ÇD��>�L�~a�Y��	�kR���^B4ש���r��=��Ӗ�;�r����Ac��:e��E��u6K&^m��������Tr�@�!w�N/�=|js�2*n|������2�;�y- �x�����SR+�5&��n?!����\�t&�8��/�&�GPTc�gaȐ�:��9̧���� ����+���P��s%�G����q{?<;�y� 7@��g�}�c�F6�ɧ�p*P����2aa���CGbjg��7�����ꤓ��I�%�.�>�����V��[���6�x��!����Ry�Z��욇�;㹹�9~����!��{l�g�h`�g� �7�[o�V���:6����x8�˗IG{���Ћ��r��j���޷褦<����4��2ξ�.T�i����6�y��u�	b����vJ5��u���
�}{F;��m<*�dyp��A:x�b���P]Ċ��6���>n�4�G�'���S���o��;����%�Jk��b8��3��A{��q�f�Y���v�L��<�_0�	~�LOYZ$0j�/�A����f���>��5�R�����]�ik�Ii�&s,�؝}�-6���ޝ;{����h�|��YpHX][�R�I�^<���1�Dđ	bSl.�A:�P�׍ՙ<�Y�ҩ�� &�wgަ.d)ن�_6ǃ���R��,�k���7p�yD2��`���!��HRo�P~�$�����֭;T{��ubvQ���[�.�8O�c@����?�6CL���N���䩹�ñ��ܭz�pf2Q��8��5�����z��(s��^��3���Wqm��p3���̛I��
k�>U7�<|��Py��܀�W�2	� ��NFHxe\ko�!�2
��h |vUf�,�����KZ��9y�0ޘ�1�9�`�	b��*���Nf�U>z~���Q꫕�IJ��_�Ah����L15Κ皲���3�=���B�i��]��[�S��ɵJ��i8��>m�����w9YR�x�@�C��m@����m��4��iY���>·�����0���.�����V��ހJ���54P�F�����p�2N����w�Ih�"S�ױ^�C!q�SA�j�;�^�����Be0> 8h�� �c!7�D�!�;����ʹ��u&)K�{g�T�����ˡ�9*��GW�{J�c�ia}��y����O���u!	�@�+���5�� 2ǈy���7����e��:^��A��P�u�ϠmF���M
]�s�jaTHΟ��C�L��.�H�����K�����k��G@�|�BX�V�����ŌR�X���R!�=N�a2���\�h�a��E�L�5�	���f����0�-���#k�>}o���9�~@��~x�ʊJ'OB�3�f�ǥ�5uE/Df��Ƥz����~�u��F�{�E�z���z�7�R}�*S"ÑeXH(����ܽ{�ٿ���+X�6![�=�r��H%�$@������
��ǥ_}�����L� ���"��,?��x�Jdwcj�'�Ѐ?�Z�eP}����Q���'|;���#=���囋�<��h `߯��]��������sSʡJ+a���	AC��M��O��
��W��п.�I6��g*�����>�k�Ǳ�'(Pd�kUY"N�a}�`��4��)m9�ߓ��#���.AT!��aB���^?������ba+$��1�li����+�pBx֭z�cݕ��H�L#׳�����ըb���e��L����S�G��W����}��E}��p=��eX�i"�,����~j��Qh��(Y�ƍF�eF٧�����5l��޹n,5��PȲ��Q�Yʪ�d�>`u�b�ҁ�Z�-$1���t�!pQ����"���a���*g��`�Y���N��v���u�{�[b��*�,$bRE�"[y+�N���}�U���$���?����{�i���a}c��ϗb�4]9H����o�O[�'�m�{�>�F�����Kƈ����:�R�3����IUXn�#º>��ϡ�E
<(��um�M.k���%�Νg��wh�Њ���ao����t�M�%�9�dͼH�k@�b��9zj��5x�	��צ��(�w�F��x�:d0S�M�ݿ��r�xpvF���3��rkݧ���&�nP���g�..�LA�GF�����F�V���%�����
UA�DO-�{$�L�{��9�Yr�G*h���FԳ��@<%w�J�*�N����D ����Ņ� ^9�9R���z"��tm�և�DM���w.�X���!|,��������m��2B���H�˝Ƣ���oxoH��T�듵2L7`�MV��5�O��L��h呥%�g�	�۩ݰN�Nɳi!}��Y��׶P
�'��Je� �ȶ,~3)4�&B��jK�	͇�̜�UTO�l	���A��0�06�X�>y�]����؆'N�CY���=^z⩤i�3�(���&�\zsDc�j|�I����6ý��R5o��d+���Л��D��<@�3���ٟД��i���/�t�u��`�|h��������q�8��>Qg�����n�h��[Jj$��;v�46�0>��j�w�d����ySR�U�gb� �� �{�B&jW@V������r��\Jk�
	XcO��W�v�kVh�-�o�D��H�*�4n+_�{��"R,�z|�E�kLe Ա_2bT62%S�~���@jX����%Ӓ0!k�MO�8H������y������y����B��t]��V�ر�hC\�_
���dM����q@�\��1�1��,�{��>H*�+�DE����]ΰ �T=���n�����1�b�I�#q�s(E�b��D%J�R�9�s7�b=�I���h,�_�:�=yJ���Q�1��z4J2���N=��)$Ua!؛���2���!�	/���p��ҹ��=�0�]06� ߽�Ϲx8X �~9n;t���k��R�Yn㲫�-L�*p�c<��p�xf=�÷n�b�r=��Q��� ӫ����[	�%�hf=.'�S�Ȃ�-�V�A"YC<$ Z sJF�t�@1��l�f]��ś:�ԸA���FM"�௟�$e���Xs���YW�_Z�z2nn�t�������>��^��8R��~��Cu��gr]�r=�*,�2��5$�ru�L|>O�lF��V��{�BPnޭ%��g (>b�" �<�קQ��5�ѹJζ%O���m{�Xz��A	Ɍ������\Y��P�ݷ��Q��?��ܻ����"��";J����?#8��`y�����3����h��\m���A?!�m�N(8(}�B�I:W�6b���r:*��r�^�|=�{3qc�ݿ�ޏnƹ����*��,Kѹ��1$w�j�^��)n�g�sZ{��D�=<O�oh�M�#C��p(��=&`z�A"�,|�s��{u�a�7��?s�f!��P���ϫF�eW3ۘ`�3��-�8j��Q���� �e��Oo��C�e�#G�2��]E8��V!��XV��0k�]��<Oh��wӿwE斄�L2�.]W�n�r*Nv�ͪ�� ��/_���G§�~>�z5��{����gK�W�g#�G9��������������H�ݻ���aHp��YUa���8��"���p�
i���LÈ4�n����'�Zx�yՄ��Q��t���o��p{��e���#�����Y<\��Ү@�Q�I>Xr����\�q��7B����;��3z-���'UT�r�"8V�%�"]�~��1�g���o���(��AV�&�$x�\���Gio���vgket�>��Z�5R� ���ev����.���S'�5.@���v ��f�'R��>��ɵO��h��)�O��_��?]��3�U�!p�J���{J��K���qNmZ��O���Νp��v��&�d�Y>L~X>|8�>s���O�l��#`a�	���I�k��A��<������קݒ4�A#���@�O j2
��^~�e���͛��w�c����Z�8�k��2CB�.*<��BT���\�;��ERnf�-�ӛ�@�
5cpJJ�qB��u�]W��3j��	X�K�4�9Ny���i��	��+'Vy�c�4f�֍
f�$ �E���h=_}�
�%���v4��(��L:S�U������jaz����"�x��TY�L�c0�l4�dԴw�+g-Hϛ��H�� ��z,��u�iS�#G�؆����/�[;��r�k�74��}��-B<+�U���N�I�1�b�	m�c�:	"����]ՠ�d��ݥ��Z��|�cT�.?��c8��[�0��Ñ�}t'��9j��Xr�ES󔈩�#�� ���"++�V�v��Ca� u�>3���+��fw���tZ��������B��#)�a��i���͐Lt��7)8��b������b�M�`��c�c
.�1�	���^CF��@?�CF�v�b�����B� ��P�(O��('*��~��}%��d3zt��-�.��+�Re�QyƿA�!*�v	����u���L,��z��h����VG�?�ZA!�����@�qB�3�D5ځ�ұ"�g���|'��G?��熳� r�!�~\X�x�C� �Sa�^G~��Ƙ���@d)qb����tl��ۅ�I1�E66�w�������y��PH�!~Bf�=( @>�Y��;�c�,'�{��0�@P:HP�Ÿ������7\q��TG�c��,���p��lLȡM� ��b"�Li%�sf�!FG�(���H^M���'���5�$O��u4��7z,�3Y�i��Fo'ۚ�))��L�N�g��m��h�n��}Z?Gt���D�rd����㫟����uyM]\��c��L'8���EG�]�2ՠѭ���m3D�\g*A�>~��=��H��ώ�+,	�?��.�016���T$�~�Q<'׹��r�m��.��}t7\�����9d��c��,+vV�U�7[;���2���7?�]�ǌ�ͅ~7
�!�4���+�0>ꉳ����y>�����Ox ���Po��E��8`c�lv����pD7���xsX>Lbćij�aW�5�t�����Dr#�V����F�T73;(����a|��O�wp��_N��.��G�pA1i�.U������EK|r�L���l��	����
�1�����*d��9��9��{c�.��X��CK�o��6
goX2+:&���+��H��D�S-��g�5rwL�;�=l/�9�i6W��V[��E��C;�XUm�f�nS��{�'X�]�8y'Z/�%A���H��cѼ�܄�ʫ� ��Ȁ�"zkk'x}~0�H�:qh'-�w��r�>]�I���p�ww��h�@�B�u��<|��_�F���`��r��
b
(��?�8ln���'a{�1O#f��<~-���̥�޴�0bF�	���@�<}>�ΜY%������'��Q�3 �����(�����{Bn6��sȲh�:���o������ҳda������
w�ݍ��o���\.�����`�=�Y�!"� �e�^��g7�//+����a$�ȡh�|\
���'Ѳ>�Qs	�N7�����Ïɜ�ӏ>�Β\��w(;y��y`)��D��(:��P������w���S���=~���=���������M:X�K;�6��Νf��L��6��	%�L�+,.��k9�-�m���T���-Psc
��Lɲ��Ͱ���8Oc�2K"�[q�&?�1.��tӣ]��ב�J��P����|,�&�൷�R��ޤ�8�"����&������U�7c�� _���	�|�m��W�	Ζ�DD�F���]Y���٭�2F�R��~�)��{Tث��h���	��8�����0�R�u�������O��_�g���kyH��ή��c���2ᢒ��� C�����ހk�.��/䡐D�BR�0�E|���'0**%��s��2��͆3��~��N�<I�v��z��+��,��Ǖ�����ùZd�*��ow��j���x[���(���1���w���ڬ��<p��R�����c�{��m����e�[� A���+�˷�����	7�q?����%�����x/o������
�y��p�ڍp�[Dj�t�M�ќ�\�;;�	R��Q@	�/���|�������>�B�(��If�ZM=������W)�*�Xq+z~�A�ۥ 6S�X��ˇ�CnF�!�m7Z�ۆY$���^l(��P$���ý�iy@��80��]��Դ㌠%�\�(���o~3z������|r�S�'bݾ͵�NG��Ba�Bm����N�uSH ��ɮ���A�Q"�����(�'b�y���p$6|xɐY�P��Cq���>+�����8zn�3c�.e3���2O\�@�!�HU�%Ћc)^�c]�fs��ހ�����ӌl�:�/ ��������[o1��N���ӧOE.�� ����A:,va�Q67���|=.N��I�\�6�x++�bv��H����҅�N�82"�,lE뼱�ΘD�M�p�!��H� 3�������	j�ݢO���SG� `K�( @���`_]'R�i�LSo�&����@C_��Rx�ͯ�����ժ[��/�E��3҄,T�s��2/\JB��Q�Ae9��e��$&�^~��S�G���d��f��g2	]��?4X8�
�A��ypH
�KG��y����磂B�������Տ?!�c|�5�TV���9�eU#��Z*�ȣ�yB8v�l�JE�x֋��!l�,*���j�܍�)w��m:!�uۓ	��0��7���kDVL�d�Ԑ�����3z��b�� L��������(��.F��ַ���o�6|�{�K�F�P�HJ���K����ٜ�RK�PQ�x�5�E��D�=�PȚd1�"v�VK+�1N����:��p��1:R����ƾgf�7��<X�p=X;@2����c�ޣv���ە&,m��JkZexp��*bȅV�tP��6��62�f.�p����z���}7��GIOC�B�����43�Z $a��I!�H<>z8]9ʺ'��'�������;,j�H��Ŏ�s��Nx�O'��}�K�]讅��.�A���1?�<$JA���x~읷i�PG����/�cǏ�S�V���?)�ׯʸ�j);�:B�W�ِA�Y�Zsԉ��ᕈ�1�^�d�omr/�E�F���q!��bx6L{/~��j���x�5�H��M �U!@�F����Yj6|T�UZ:	?.OG�ۜ`�˳�ɗ2:�������_��_Q�qN|���Ȭ����W._a<���?��d��Q�"�4�he������k*��I�`�^/��NG�6Ҁ��X�)s�\8�����᠍�
����P��:�h���U�9y}�w�b��.��1~�A��6ޫ�\lx'� ����v��m�p���ۓ/!@8��$��ߏ_.]���=�1CJ	,Ÿ���Q�}tq~�Z%����8�DX9~B(��SC�\ox%G��������--��J#.����+�v�Y��vm�uh��5uj ���,(1=��!�s��8x{�+���:��N�Kx1x?�?��?r�I,�S̮����{��Br��32c9���T�0TAk�rU��3�����/*#o��f��z�	W7˛}�=TҒ*��!�0��%��p�a8v�]�4�s���a�wz�c�ax]8?���_��_����V%����}|��^��<0��W�
�|r5ܽs�=��c��T��������b��G�*d��\%YȽ�S�X��X7|.�lu\�0�#4B�E-(% {N�����M�����D��Y�k3�͒��c����OuS=�S$���o|�MN"awX����Q3�I�� p�ma5pt+A�b\�*[Gs%d�N@Y���=�Ѱ��g���}e�蛰�s����	������:�J���F]A�DQě�qԅ�I��0�ӑ���.\�@����pb�d��O~�I�L	�y���%j�v���@�$!�sfJk�#+v�,��Z!�V�������J�ϙLͬ�=ɉ��Hzgu�!
�u������+!P8RLY�}+�$��ԥ�t��/������?�!ҎǺ8#��
����a� �8���F�K��o�_����������ɑ�J�,���M�m�	�1Q"sK>1%���(� 7�g�=p��,m���J(��h���"�t�e�ͳ^�[�2~4�m0< �~v$Op��x.��b�g\�����,[�ϰ>8ȅ	-���LV�/��C���3���,Vl`���P�G�*�-�߷K�!�7~
K&a����foO5�\�Ņ�E7�F8g�UVGi)��,꣋���<���b�2M������$s���6]�o{I��^� i��ު��6�4�+��i�:*/�3�'rK4�H�CXZn�i������Rd�~-��n ��tݶִ��Y�+7KM>��]�UM@R�{��o�7��Y�k�3qУ�R�V���1�� ��={.�x����qK��ݮ�&k�t�����f�R�o��V�[���6ɘX��S"��BxohN5�#y���1�d�w���-�k��6��y���$�)�S{���`���z\F�"ց�.m�:���>�zM=�#��ᣦ�����H$���Wei !~��v����^�$H�i�wDZj)m	�H�ͽ�$�ch"
����/,/��;�}��0=�(ǕOpnCN��+zi`��9*�?P]X�7����@9�]���f���x�ŵj�'�)��$�����6�D�!���>��J�����QZ%�c$o�{�=yG�i�"�:{>�si�s	��'�'1[��N�]����"�C���_�!�)2�4��ϡ�O�
��:��o�ii�N:�.\'O���(���% ��UsP�8���X����:,���m�ֻ5W��6�k� "���KֈQY�>�+��I]H��N�G�k�9.��n�vW����q
$��zag�M�{��C���nm1���v<.S�I��NI,X@���(:��X��M������M"P+S�"�B��Gr���tD;�C�9>�������X|��%�<1%b��.��H+x8� ���$�@�׭c2A.)[}��՘Aɼ�Ѽn�SOZ��#��Y�ŕ�J�twm�V�����A��7o�-OQj����:��P���X�<���yL\�NC5�Ff�Q4h"�8E���S1ܻ�����r,z�	�`�r2���m�Q��τAz������*��Tm�2�E�2���ix���\���>� �f-`] �xݝ�7S)P��q㽻�x�z=m�fi�����t�t�{�;Q]H-���n�����F�T7�ѱ�۸Yݣp xhָ��0<��Y҂`�B!�
��������Q��ϱ�����.L�ܡup�!��};��c&��{N{�y\��s����~n��em9��
�z���y�o�`�[6��^��GѾ���~�����`sq_�'��im\����o���]�z�#Lܽ��냶%��^����%'�Q(!����Q�`2� �C<���ճ40EP�@Km�rs3�6E$�-��~�[���쀟m�+�>���WH <<�G[���b� *��M#��%� �ׯ�_.��a
2�\�|�ڦ�����'l�y������ں����?���w�2u�}:���wɾ�/���ٗ�������M���G��/~�iW���,������kac}�SB�^	��Ϭ]�]'%��,�̅ίɚ��Kf;_�7��Ǒ�����ں(.l�UԶ�T��en�k�̘�J����-�4�k^���=�7>y"�P��8�=;�<�F����A�zR�S>y�����{�g��9����/���z4y�?T���z�����?��Ͽ�ᙲ��Qb,��s�5�ŋ���#G٩�ph�����Ldב��U����\a��>�#�l⧮a�5t��z'����,oޓ=��p�lz�(�2� �V��Rn�$K�]�JG��q-|$��C����G�遼�����r
��?�%�m� |e�"|eK���v��Ox�#��L
�?�U�uA��P�$�([9&��,�r�qV��cgB˃���y��FY��=����y��Ե�\��;4W�g Ɛ�8y����"g���CSry����/X�M�P�(��9g){��G�ίʾ����{_���B�~����W�x�g~�M[��w�d����q��A~�����������>�3ص������<B�VƢP�^7>�hg��/!,)�]7�`I9�Us7��irz�m=���a��
ٟ�"�
j\�'={�0�ss��M������
�ӿ�Q����+�z����?B<��-�C'J�!��ַ�z��1@$Y⁫�C�+����@�Q��X�ډ	�{���|��^3�Z�g�=֯��������j<TN)l.�fx�N˦��0U5��g�}��~�����;���֖����3����������W(�_�/�{��W��.#M)�����&��˳��܅�t3;�f����10ETQ��qT5k&��f%��	��+[x� QS~Vl�BXiAf'Cد<���D��� kzs`��-5g��Rw9�h�2�㱸��o�!Si�)�����^���'x�����>�Yo�DOZ>�<A
	���` x��S���ѣ	x�J�h��C-o���j@�
����g���%�
� �T��R��<�fM2ռ�HJ!{���Ȃ���<T�"��9�%�5�vUm`	��T��O���R*���1��O}��@��+��v��{�/.�yor��B�X&�%�\Y� �`U�P���Gm�즐�~8�k?��3��8�Y0���Ϛ�ξsg?OC:���q�}�U����Wy;i��zh_���]��/�������I��O��'�cf�-���o=��f]3s�k����f�_�{��e&wS��9�퐋����K�����m3)���I]4J�G���[�?�i�C���(�d��M���%���{����r����D��S:���-9��J�C��?��O��%�_�c:��~~��/z��G���0�gx�#s��^�`�    IEND�B`�PK
     ˡ�Zp�"^��  ��  /   images/f159b6d4-7cee-4dce-98d3-76d280a06797.png�PNG

   IHDR   c   �   !��d   gAMA  ���a   	pHYs  t  t�fx  �CIDATx���g�d�u&x^�KW�WuU���@h8H���FK��f4�����]�v��"�?V�)B�!�DIC#J$Eo@x��n�Fh����Y�3ߞ����*6h,VW��g�q߱ׯT*��W�y"�JYG�o��Q~�y��C�Y`���������D���zf{���~S�]	���K�w�������/�����{]��۝����k�����s�0k��%�^�"�~���
/���D��H$������F��b.>�D����ܕk��?7�E�J�Ȏϣ�ڿ���y~-�;�ݎu�p�v,����=G�q���Y�r�$eeZ�!ω{�=2�9$��Dɀ�D�y��dyyY��i�粒�f$_(�H�R�TN$����	=&'�LF���'/��E��(9&���w4���Mijj�t:MN���l����*�P� �TR2z͜~�����b�<��V������k�������Jn�X���W��Α��$��ň�Z�7�%�N�q}�|!ǿ���>^e]����nE��ejj���}���s��s������B^�H�>���ʃ>�Ǘõ�w�޻�.��������NI��������~�-6N�����.�@8g�T��qS��W"�X�� %�R�,nW(�4�}�;�k���󸭭-)�\�X<�s� `H��.�W,�b����3�����s�*n������9�y+es>�In�tvv�o�AN7�	U�*vKp�e���9��WW����t�zx�\���P�����y�����h���oDN
ჷ��K���� �c��E�ʅ���Y"䴸.$8�;L��$���b�H�X���o<|kk�$Ad�/�ex��&�fr�x,�T]9�������y܊ϲ٬Q��h�O�6����ⓘJ<�j��S$D6�R!�67���Z,���ml`�kDp��)��䥗^�?��?�?��?���.#�I\����-kk��~@Ւ��b�#lO�"��� �,UĔ�Lo�򁜄E�*9�w��N�D���.���m>ħ�+[Cn���f�G�1k,U�d�\4cE�^64C�{yyM�ᙷ<o����#;���U�n`��f2���N�W�E^�������2�X��M�,q��!vz+���h���o|�*D�����~�����h�,u�"��"Q�l�AGH� �օ��z��ll��F�d�CH�;B�
x��H���,V9�SE�j����C.���3<�[G.�x2�v�q�*��@:;i� �s\!/4�N�D"�8��yF���=�\�	�E�J�T2!����M%+����VW6evfE��W%W��Q�я~D���?�S���O��ڐ�T\�ꥵ-)���آz�I��u�⡡qY�_��!<�O��g�MC�E,t�7��!=�[Dܱb���OTcIp�x�S���2H���
9�g�r����=���B�f�=$f�jGy���|�߼�h�j�����*�LƤ��[N�<.����=���z�ե�U�~��|��5��J<��#��� ��Ԅ"�uեE��n�f%F��̩����w�~;bܑo�2::F��T��EB��� R�F�B������}�a��_U���
u���Z�>�3�;�l-D�%p��2Y�l�b�����Խ��S��ޞ�����ݝ2���ڽ�_�;�#T� ��[�g�j�T��[ꥭ�Q���G��ӧ�W�8&x�Ԑutv(��7�Ϸ�d"5:��C����3e�-����ǺŮ�lG�߱�a��9������Z���ƦE�����z�婧>.]Q*SD�U��ʺB���i�e���LZ�i�;���ߣz@TN���bNv����ӧ�]0pL�쫱.�;�b�C�ߎxF�G�J�_� �������T�Z��/#R��vRT=�H������ꕉ�HgG�AdѨ(^$�U�����t�_~If��B���*��F��MM�r��)��:u�2��ѡ�P��;&/�Y���ıc����b�ma]X�=t��e��H|�"־>,��I���������޿�?��S���W%�	,���.Z��vuu��t����]��x�4��ϖ�Nilh����(�I	o�Y}���qj�#|�Z[��a��I��8�È�}�.����<�N������e�����vM?��)Y<x�m�1,}��R�l��?"�Ql�7��%�
���X���pAA}�K@]���лţ~��n�X�}������:1�TKt�Pf[諭�sE�d�~A&'����64R�v�E$<�9���Դ,,,�8��A�|�,+���Q��)ɫ�H�7�b��t��5��+���߅���n���kh�h�B�-�[E�:���|�5<˱�|pE:������z����L��W(������Ii	��M�����r29� kz@sk���xV/�Uh;.������� 	k7vC�݋�����Skf�wۉ�!qw�Aj󫠮����M0x.��d\%�;���|�s�S_��̪�H\�U�e�3��O�E�Qb�|QJ���R+��*ɠ�o��tw����Ac?J��D���؏��r�c��B���n�Z��sx�>v7Bڍ�~٢zwy��<�LR�j��h��o(��?��988��3\�����_�?�Oy6��T?/�A�es��?���My��M K)���D�t��7dyeURuIFg�>��]�쯋��w�F������Ң�NU�[��휿H�j�W�g�/Ʀ�㈪}����3��[+�J�J�:wی���5P��R�5<����/�L.\x�
�D.�!쁰7`�1D�ҹ����&���>�ο�F���4	��m�k��Fnwd��9�ƨWAH&���tFL��L
_�m�c�]��3p��O)�Qc����3�1�f�Ƃ����f��+�sT��I���Ϝ qU	حjv�H��M��.�0Q��Ԟ?5Em�)�.U�����o�T��&H�B:�%�@�I���FDMۥ�+6��k3͵w7���_���۹ο�z�@[~�k��X�{��q�٭��f�v�v��k��eRn��%��ٳһg�lm�+Jmן%������J�
m��w&ߐ�1�x\1s9"�|�&7A	,躐�<���Ҭ��?�/�~��~Bsư�>�fq?��Ǟ&�({w�����m��^YY�|.�f�(q������P�� �t^�g��؍���%�	ٻ�O�[��x+5W�e;�Qj�)����"^��:��_�Uvr��8�Q+R� w[�@j��N���=0
XyEv�^e��6��cH>\`~�\ED�O�!>~f4�0璈����|6�J���޺@e`S	B�t�������d��]��`��>Iikn���&��o��xO8Ư蝶47ʑ#���EJE�2:2N���Q��}/*���+��+ʒV�����۵�O�ꍇD�6��D\H��R����oN�����[��@�rvv�栍w[�),1ypnP�X�(�|�1I�E~��I3���){I}*��}�	)(:��O/�:(g#���f`Ҩaٍ}g��w{['cNݽ��ذgqimn���:�l���Ꚕ��ҭ(pJo����K11k_ȗ��� `rrF��}�ԓ��tZ����"S�3a5�g�<��J�dł����$��_��u6�fS"U�r�C5�b��+\Ш���������5�[�����g���QĜ˼e,*��?�O�#^���"~Bc}��@�����eɉ1��"��¤���x��A���99~�:�K�x���0�X�����v�3\O��W�IE&_@�
%8)����7o�M&����ih����aY[_Q�g�z��
}QgqD6��m��dv�+nQ��!/��0[ED.Xiћg�׬P)��˗X�?=5C��UL��,5��:q�}pvEU[E~��˺�e2�	���,Ծ�_������dkc���$��^"�o�d^��j��R�H�U5��7oɆ">䀚�[�t�%X\X�)��>����!�~�{������YY][��ʵw��O���R�U::�elYAS���O)�[��J]ϗ0��ࢿ.�	'W\tپ`'	����k��a�~Y޼��K������L��߁�=Q5-��۩�=%U5,-���]��m��h��}V�YYZZ��JС{�`u��e����v�z޲�X�˞����PUt��=������a%b\��7�ʵ����/�=�n[26>%E%DR	�4!_�ݸqS���MH8&�bFR�z9p`@�m��4���
g#�GG��MK,RP�ʩ�r�ޓ�f��9���*��R�j%b�{ԏ],5A<k#�r	W��
�șPvјQ"����׊�*?��ׅC��a�@�h��Z�^�>��C���S��׶TM��k�]T�l��PQ�(!��;�����y�<�=�!���Όȝ�iU�1X����Q>����%�PQ6���4�/�i��My����_|�-}����07#�ܚ�m��ֽRQ�蓏HcSua"�Q;�`�Ҭ;��5��fc!x�V��C��jT�@nF����EV%V��u٬4B��+G��(�璩��c�#4���bA��b��2=6���/����ի���S`� �YV��V4�D|�uPMs�sO�� ��'��L.(ưR�Q�Tb|�_gR�%�� R&�1]l��Jr��y��	�54,q��R.K�-�J���?�U�E�>��B.��]�,��e8�bl�p/�ȄB���)��iJ��]��M��|�RĔ�Rʂ2����AF�`�ʅ
k�"zouҹ�W�v�I2Q/'N����=oh��#SjW'dtxH��; G��əYu�r233GIŚēu��	Jn���������Ӆ�EW���E4b�3$b�x��O>x�<��3
#��^'7�;/3���%���;�T6�
�+;/70�6��R�^a�h{��&�b�@�B��~����PG���k&���9rᵩ�4[j�����kY�UCs��))�W�C�$��#]�T�b24xS8�����#O~�Yy��{���|GRɔ�z�FeLm������x1+F�Wﰳ�]z{�e[=�I5��i����/��k?�//� �6˱cGU�i%*�98 ^A=�"*��TQ���r���هN�g��bW����S}(�q%�8R`���^�,���⤑*�s�у��t���DM���de����*�Ï�4\����	%N\ҙ��)���54'%����&9}(Imŭ�;R,�髫KJ��\أ���iT�F�Y4L���G�k�z�g�ޣh�GCA!k���MJN��<+MM-��_~�PlbbB�^��VD��{zdH֗��Q�sgoh���b���� ���V��<D�چ����gm$A�kr+j��KV\T�xkk��r^2� ���)�A"Ϭ�-۠_ UHmt:�t`j��E�����e���\Ad~� Y�����&����C���Qu	���r�7�K��j�c�:�U��Holl�����tuw����s*��tu�ra���޽�;���p;�.ss���/Yo�(��Q9{� K�� �ntw%+�+6�0Fc��Q�P!�#�A`K�˵)�j<)��\h��;��Y��b�����!ڢ����r���W]6��g���'P�����ܲ��G��< AD�H�=vXפ�y<_��ߺlppH:��J��W�N�k�S �֩>[\XVΟ����l����F�;nilh�Cj7"����"r�=�eoW��*6��Kuv"Rm�.��C��Ui1ר�'�8�� W��h�/�E[��wz+��EW�QI�Sݔmͮ��۝�$˳�g����Bzфվrz��ٳGN��O�>\���u�=|G.�~^�ʘ�ۇ��,/-SC��[XX���SSS��;��Э���d�6ַ��W��R����( CD�\�!=tN�⯮,�b������K]L��)AC߳i�r|�b7!�5\e�+
�ᄰ5�Z�떈mU�.�9*��ך9ua
�!{6\m���Y�b�.jҨ�����/�ۀ�%#]�r���$�T���)�:D`�߿@��}��lfT��H��$��MH�d�FLܡ�R4<4)S���Ee��@A��m�lg�[���,��Gi���U�Y�XZR�Q���|�&]S�m�agH=�z��A+.��Y5S�����C%��JX9�l��j��!\Ū�H�!�z�.tP1�R�r�i&�]�",�?���gONLʬ����m%F�����OA�;H�}�����. D���!��)�:ˢ�%j�t�g�)2���y^�$�"���n�BL��#�1���~E��'+oKwKL��RMm�����F�,��"V��a��,�#�	�:d�J���
�(��6�ǹC� 4RY��*�w���{`
�}�8ӫ�[�]R����[[Վ0Ң����T�������{�R�������*ձ���%@�ɒ�K��"��"6��/@V/$Ա��;���������������+!|i��ȓ�~Db^L�gl�ު����
�%U�$�#a�b��&�"��8ڰyŖP���q�*�N8M��Yj�E<_���[0�g��	ٗ)A*!�G)���X�a��ԩ�rD9��ɂ,�n���<+�O;.'��TTZ'.^d1�W"��J�2|D п�΂h��hw !VA�!|��ػ�_>�OP,������:5���S'�+Ǥ�E��ָ���&IĈ��q�mԂGĄxB�q�E���*�R�j�.�]p��(.ZV�El@qgћ����n�[5�\�`��&w��F�N����.�����M������@�ɹE�q�ܺyC��%����r����O(zj�6� *�s��Q������������pkk���I΁������Q��Rr��)58	iid�����G�oz���y6� �ѳWW�T�$B��Z#|�k��Sņ�%����]��]�w�U=���Q��8�s
�W�zc�&Y�Z�Ń��n^��[�����M��!�X+)�Jɬ"�VP�gO���C=��44�ɸq�����O�/4���.c�344��yE).>��8lqaA�_�.I�N��y�����-ɗ�a��j��"B���
��9E�������vAmV�e7��Q)�+��3���*�q�0Hm�BmR�Dg�$~ةj�kV�I���Øg�PS/03;-����JrB��$���+�4����dO���:�&DjI�$N�$�pw��m]c����� t��oPL�eEu.[�K�ޕ��Ey�'��]^\�EEP_��Wƥ�-&O~䄘���u�v7�ݰH��ደ�7Bq7\k%���h#���Ɔ����5Յw�p�c��T�β�����RDX`|S�T���9[�������.�Ν����[�͘W�Mפ]?�$et���l3�D���##c�_C��h�Hfe������WqT}?66JC���e�}��}r��Ay뭷dzz�|Hqt_�T
������>���`��.S�����ā���0+6���D��A��L���%�p:ir�lj�"bT��^,,��+��#.΋��G�Ύ�y��F+6�Qb�,ρ����>0p@�L��{��U���~���������nS�m��ՙ�V�Sϖ
���Ҫ��}0+$��B,/�ʝ�a���Q�<Ǜ��N�����P̉2*?�[��D�N�[�����W�&�L�:99���"���H,b��mڀ��'W���ICt�C�Go��tCr�@�N���Bj<Z��qy��i؇M��(�#|����v%L�x�Qb��-PG���Y_[���.8,+�MpN��@���ֺ|���`z�$
�o*�v�@���ƻh���\?8y������ȫj��L��0H��@r�[����
���ڶ�\�̭/�;���d� Y}]�l9GB΁S�A�A'�P2��7�Y� ��08��� ��[�� t.�n|��#,{H��8����FQux��Wnn��uq.s=<D�	5I��(u�V��kf`thxL�9#��nʂB�e]��׮���� �b�T�$LIUc����	���P�A}PIr*!^$�j��~FBΜ9#��],��79���¼�˿��ݼ��uiV_c{-��3��Y"�i��B cV,a����
�Cs�>l�	8�n�D�=pom{�	`&�˿�xB��8�=H�PTf�sJ*��n�I.���\J��,ڐ�QV�Oq`��Ȩ�#"�S˲�<J��4(�(�o�c&E�$�e"��/����f�a�Ǉ��GM~�9g�@��9z��<��c��+?3��,��ܾu�`���|����\�5a����oC���]�r�+��@g�-B�Xԕ��Q�h#�	2mW���<�5�����ؚ�-^@4.o�J)r�c��f��
]�l��G13�3S�y�	���18%˛��l����T:ڛ��JE�%��Y-�[	�"[(0'��OtB��/ ���*��El҂����U}�p�O����ǟ!�Kd��WTU�B�m2l�pq��XHa�B���:�`��Loqq�ʙ�B��Vk_�r
�p�6�A�Z_ål��36�I�	ח��Wi*=��D*ַ�7�����Js+�|�d|f^}�%����>(�ȓD`Ͽ�܀�����X����7�r����\x�~\$~�z{$���E��6�����'��(}�g���ʕ+T@Y%Ճ�ɬ,���<9z�	7^����p�U����`x�����]�Z[��^��ҥ���rL��sׂ�6ݩƙ�L 9�.�L��!>�,���K����LLNHoY�Q��&��o�^2ncs�}[=s��Fu�{����N��[R���6 �-�ꦟ9s��IZ����YYR_	�18xG���P߮���ի���ۖ��aIDӲ��-�R<|�0��~�dSaK��掶߰�]j
���R!EP�,,���j��Xl,4
>Q�:�gh�}�1��8��� ����o�(�Q�\-����4���ss��_ӷ�V㝓���=@I�Q)8P�*kֶ{5�كI #�շCdtl��	���!�F�ԡ�hi�ek;�E���U�Q?c�*���K�K��U�h�5���GO��bJ�?Π��!L�>j>s�ZO�y�)@F�f�`��r=>Â�P`�S֪9�"(��̚����{�w�� CM���z(0�ڐr��o����V�Z���$�u�y��a7z���Ԟ����A���5�eEQ�j��:�|tȂa�6}<0�`1�������_�� ���|pE��^���#���J�&98pP���_N��/�}�\�tՔqیB"��(��k	R�~-A��v�X��P"Ը;�������Ƌ�
5�xH��3=u&M[�^W�Iu�D�@���! �ū�O,�@�fDte��:G�_�VD5/#���.���7��������I�4���4��L��`�~qe]n�fjem�)�UU�&NOO1�����:n�������?"�����*W�{Uuf��r��Wdƽ��q\[�z\��gw,UD܌ƃ]�SՀ�\�T$a��ʕ�@�xJ{�H%�W�h@TP����*�(#�h��!W�P��B�%%X%�T�f:#��]���,�j#�I��~�o��!��!�3���Q�\�Wt-Ӫ5┢b��Y�� KL"I�|"4�}��?�(��`|	����Wo�g�%�хq��i0t�a�+$,Ŭ��T�[X�!G�J��9	)�~~��8}Iٻw/Q*Wj�1�>W�RC�Eߣ�mm8߭-�3�w�/b�l�p�ip�%]џtF㭼,��f�mB�~��AES?�a���
�6�3�4�������BO�`~~��p̅�@E� t$*��Ŭ·)����;�Ҳ��^���q�q�����R��n���!s_���j��9u�[g��ǁ�����9z�iX�l����L����bL�y���F~�AuN�@]Uҧ߰��&�A�orfUՙ:�Ϩ�E=A$:�*����)I+؁)�������N��7Y2��*�݂���Or���o��6o�3��u��VwZn��a~���WH�ڐvv;nf,]���4Fe���m��&��X���֣��G�d}m���|R�鱫jg7s���zݫ�>7���4�ʪj��>y\U5�����Y���)��I��<��k��R�����ԝd<e�2��T���&"��HC/�Q���A
��ˌ;�U��w/��K0������E��o��dmyX"*%�&s�C%�^j���x��F����&G�Ug����p�ٙ.481���� �� �_8�*�ф�ج��Z��PBl��=�R�o����dJU�!��z�tY�U�� g��>�ő!�����nkkb#�V>���s&t�*�dD��viU7�(�~�ŵ�eb��+��ʇfF�W�Kߞ&)d�%�Y`�'�!��uȜT�:qN�@@@;�#�T��zV!|�w�����o��r�V������\>�I��Gf�46��sf	R�mט��3�l����!�ykp�6è�
��h�Na�޽��`l^{G��u�u��-,��s玸�aT�(No���}�L%����I�UC��K�� �H↡?���3�r~sN�y��X n�QCb���Z�1U  p�c��ֆ�` %,ԍDō;o�F�O��b%rg&0�6V�Wd%(�$��;��Ih��4� M�ClQE"n�Pj�u�3+
���<�eYȆ�d �x�� ��Ih���B剉q�Р�QC���;�_�q�Ȭ��+g��ƍ���Յ��P::� 9hP9��֘<���,j��ʀ�E'����8����F߯�Xk&9�c�4e��avs�g�..f�;��nײ+z0yxal�63�(�Ί���qbK��11�&(6��=rP� �(�-GTMh�9��ݧϗ��@��:�X�22:)��yi�u2R�yS5@�uq�ݼAw޴)F���xq�gGG�]�=]���U��45�R��,ͭ��W��"qU�%P�����d��㖲�+��`'��Ԑ��~'h���rx���%|v���&��4b�p-�s�H�[���*��"�����#�Q<y�ɲ�����Ԝ����x~6����� ;F����[Z\㳬(�c�*9Ugcc[���6��ZL܆#]*��Rw�� E�p�>%��̧$�����W�b����!���ī>�����
!�B�(*�!	����x��o�g�qL�vFa�{{{ކSB���uP �pw����q�{e>ߩ/[�bZ���[YV�pD�Q"��s/�������ׇ�c�j��tE�l�3�索O�#��,���dX>��(�����}��
��)E74����c�R��ޠͳ�0�j�&��lE�a���Ϡ'q�Ы�`�<ҤFw;Մ5i�|x~�ze�k>�E��.��I��Mpn;$J�d�U��x�墉>�q��C"������l >�����^!&ź+��Aţ�-DT�_����Q�(��U�Dd��(���4FP}yyI^x���̕min��^���P�T0��z�X0�MYU��#�ˁ;�-�� �|�[d��p,:0��� aq-|�Lt0���cw~GSqpQ��ʅ��C?DJ�kk�r��u�^/�p�`�?~L�eKM���P��s��@���p��aJ#+v!�y.���Ux�{��A������cJ��{���ES��'m�1�*^��e����p!&\�@@Vx���p�� ���w��Ź��8��JP�u�m%`T!	���`���Z���a�B�! J�#�<VZ>����˲��j^m�����=�{�w�wY�t����ߙ� E�XK�B`U[�~�3�2�M3�ARX&�������o\�~S~���rH	���b�:z}=�*Us��Ȳ-,��RD�3ak3uX@,0�@l�م6`�A@[�15�H��:�P�w��[�Z��;W]�����
���bw@u�(rٖQq���,�D��F���O�X��
}%���-�BI5ACJ��>ۚfr�x���"ێi��ٴq����֢��~x���#����~���W�[b�_{g��Ϯ�����<���ĩ1�(Ԉ[|���u�^&�V�'X�$:�s��Aa��9rGn%⹒OW2��8�f&�6��`~&j�h�x�>0��B�\��7�D��ͭMy��Y�R�\���$���
	��ЬнG�`�k�����j�O�<&���-�/�Qe�D6[��=�	�p�x�79?�&\�%��MeUW
��ծ��p�܂���)M����q��l�Nf��f�;ZClwWR�g�s/ݓz�K�HH��R87*aJ�����\��-� )��O�E6棗�L`�����>��lg�2��!Q��t6O�hh��O|�c���ܹuS�GJ���;~Bϙ���Q��I>��TC9N�z�-j���2�^VO���Cc� WkkQ���7�U�7'�qy��{�-PCSs�x.��|�~v^�S7�@�N{{{�i>�q��� H��)�V�E���Q71�S�{���[��@%�F��52?�(�Rު�����3�ۯv���x�B�4���'��8���h�����u��ұ#	��r��!����߿&�cS98�������uG	(�'E�I[sJN���	�y{h2!������ˮU].��p�EXP�h�\��El��O�@@��ф�a�YF��)��S^&�*�?� Cc����߮�x��jF�_�w��������7~�Y�`j�#���O� �2>1�L���-cW�����y�=�Y���A����Ĭ�ίW��`��33�2;��o���:t���o_�\�rY��'��=�:�]��#�.��*!j�](3/�Td<]�3��W�n���Z\��E[����Cmi��p����
�g��L	�	4
��F���#W��k8	E���De;cmӍ�����elM@cc='��6Kb!!���W�KK�����#c��8±Eԙh
ɣ|��FzL}
x����Dn��@GO���fg�lpJ�M�ć8K��IjU�[@��8��:�k�G�x-8�-Rs�6Ad�v�溙&����@"� Lh���&ekS�t�j���(���?��������|���0M>�-o\X�&��Ƿs��Ψ�����ܨq�Ѝ�����}Q,g<��s�C���?~Yu��v�,=���0/�{����j��-j.ݱX�M-�T�AE���$�rgMj�r�ЋCM����d�)N���@�n;^�r��T?0���)�b��ų�J�M{ZN}��\���%Sa/FK�W�4�U)�Ц�p�����4;|)1�����8�o<��How�<��9u��e}3mn�FH�E܂�s�����U�8(�=զ]wvG����6Cꍨ���#��p�^2����4d��܇�=�(��RtgtR6���[��������?��dT"ꙏ����e�cὙ�)�L5%��3�+f�Z���/#��b1TY�ڊ?�/�r{��eivDV�c�&�1~h>�@͕�y<�$$���quJ�Sv�N�t����M@Kq;�T�o�iMe%���Ɛ�ٴ+jk�]r,b����Mt��U���!���|���w�}�����G������/�Ԯ�2��4ᔨ�*���G"�����>���M�ƛ[���~���������9�*�Rc�B�+*��2���!싫k�2H�j��B��J5|���Dw� ��vCb�y��5��#µ�%.>VK@#���6���G��V V�H�6}��~����wRryTɬ�)�J�P��V?�mH�"1נ^�x���b�n��$�(>��t�����ʨA�4�PU3�3��o�30l9s����$��9iiT:���p��v��Ty�i/f[ ���*6xh��j���ֆNvۏ�p�X��3w�jMR��5��6^��U	��q�R���/��d�`���#B@Y}���(�^Gg]dU���dP]��G�Y�ҫX�<�_�)�
s�Y�E������7o��`R��3��}��n��<zR�T*Rͭ,Z�m�2�?�8#���<�-6yS���`�yx�ª��9�Ȱs��5Dj���-�������@�M�	
��K&��
z����ަ��C�eQ݁�%�L��8~\��'�e����Pk�D��s-����A�}}c��dfv��"n�-���Mm, �7��\�;�^J��cG:�v�OΘ
�1C�0E}����<��E��$�y��B���ww���:��`�
*;�*����%���r��vT�U\r ������U��S��o~��څ�Tem3�
Ȏ���yǽ�i��z���z�8��]K<zs0��ƍA���T�ʾ�f��#G���I(��(���}�OZZ:��Γ+�bث��@O�Ũ���x�V��PV���zvg��fA�4Tђ��ڿka���6�^{��x��N���J��wN�hl�����Ӆӈ|8�iݞm{c�Y��O��
�����0�O;	��]c#��I��3_4��"	�@(���W�_�"{���� lm1M7�ٶ�w�VT�qEe��i߾��O?�1��)��57�h�Vw��F���s���z��i:\����d'��C�*b��@ѹ��)�Y�gǴ��Uy��7���sv�E�E����B�Ͼ��AI@1B��M}0 ,���	n�<�-�Kv�:��3���"������W���3/+iI�E��W'�s��;p���#D�|]������;|��"�O}�j����R*X\lQgm��-x�4�ı���U�8������9�)�B��8����d<!&Xh�,�c��QE�PO`�����T�)�����nn�4�a��Z�������4J@�\j?9���W�0ވח�L��|!xa��˯*N~�]��\��n�=Iԥ�����ɣ����F%S�Ք�T�,�*�U��G��1�>�)��l+4w:�7�f�XS�����"=g�f�9�Ĝ����C')Y��;&��;�����m4�+��Ԡc����M	��c���g>�q�T���֥>�i��0cS��Ǔ�pJ����
��Q5��sҝ+���q�j�FU��%Mk,gJ�(�x5��
� n���G���P��x�:Zdi��4�6�����Ƕ�;0}�=� c2q]���W�`�LQ㌧��1?�h:�$"W���m�8��v�J����c�P�+&���7
礃�nc��HZx��a�����f�K�}�R��'��7�ę{e;_T4���nmm������!�nޑ�����͍TQ���ޠ^*͠Gu>QK�JŤ���ATBL�\�3U!����C;\yL�� �QL��#�u�z�kfW��u�������g�?#��6	��2a�a��=}���Ԍ5��u���2��N����1ͫ�A<��0c�3p���L�0��Q&��]йb��`�<{.C�A�!�˗/��ȄL�-��{�<����Rb��;MTU�BA��<� )F�MT���,g��N��s����y"��O}�
�țo�Egejb���K�H~3#^.-����lٶdX �YB�\��%�|(�W5���*A8"�Ǻ�>q���S�
Bb�]*�%�Ǿ;,:�r�L3~E��F����q%7r<N���B��Kft��=|�8��8���5�&&��z.[���E����C;�T��.y���adS�l����cTG82:BqSQ�l�P�ԩ�G��>�rU��FN�K�&@<J>��b<���-��^Y�膖>�RF��-�3�b[��]%͍���f<)�!߲T[��1��DԼk���p	��
r|�Ob���V2%�8�59^��d�׎{a�a�c���(Ů$3��H&l-�O�V7�N�݂>���=i�^�y��7�����Ё�����g�9�W3��:�U�l�þF��9fa;�3%1z{�6"�q���
c�kҩp���zR����Mzz1�Nff�̞B^����"g �a���v���2�p�$#�j�����i�@,a�&�ɗ�;j����Ī���]d��ڭ$[\3���"��`���gz)��IU\!�������l�/|��>E�T������a(ĳ������Bŀ�f% ���W�=���+r����omd����M-��/�ٳ�K[�I2�����o�ҩ�����R���9ʜq��T���g�SQ(X��n�{�8������+��9(PM��lzYBy�.|}*���D�<V*f�x��W�8>"b�g���pz��n*�����kq���-��f{����U�]������^H�"C���@���_R&�<�Ly�N�3���J��=@z�Nb Z	�y���LM���c�G'F�PH(�>s��N�f��s�%�S���%������2�tK�ǧ���1��"�Þ�n+RK��9�3��ɺӕ0b�x��R���ƂErs3>*+Eq;Dbsx�����Յ�+E�V=��@+���;��D�Q��Fj#��PHE%�6�jцˑ�����F�	�7G�W]�y��7eQ�Q�f^����B���e�l��&�gTJvؾOF��̄�<�{�X챴4bs�F� �hiA�����]ܑ[F8x�v�lOoU
��}�����F�U�Tdg�&����[7�{�p������ȑ�� ��z\��=�����g� I�#�Tô3؈2�1����z%hB9iYvM�D���b|uJ�r�ʽJ��n3�M����Y���: L @|���Lx+�FvK���e$�7苍<�R`@O������U�~�2XE޹|S%cV��[^y�*��J~�qEX+jK7djr��ޕ!_�'�\�C�C��ḩ'����+�т�c4t\���'h���CԱ�uD��2ev�<�~
���%���nK�Xb����5^A2\k��wGAē%�ŹEim�\u���A��d��E�ؘa����Ũ3=���:�M�a���Ҳܸ����)	�6�R �T��H;���-�Si���{�p�3sܕ-��BueL��=��,�F�
�]�m�n��ɓ'�O�Z奩�E���oY�,KcS#CAXKP��P�O�"�D\R*���3S.����^��G�)'7q���M���N֭��X�5e�Q�cP�����{��@��B`�����e�pai��E	����Gz:�L|Ս[����ۭ*�l��Qq���K)Fo�(S��b�M,bڌ7��]�1�}��f��ꡭ�?��R���St�gƜ��]W5�:Z3�ɤ_1ZU���� F�_�عX���e.��g���SJU2�4�-�v�j8}.��cq�ͺ��{�_6vCz	��VW��ڵ�����n�d�7�]�8i���Tj�|�j6ςqFû� �̷3ٲ�����%�A�r��aiji������{��K?�|EV�h�����U_IU7�����G������cJ~����P�2��c`���Ҭ���{WoI]�^�:�ϴ�=���ԧ?/�#��S����9s�� Y��C#�r��}r��C�Ak�^EiSXP�k�P�����t����&8�~�P:*!A��mdR0��[�l��d�:;�Ix��a���M(��#��(h�7�m���ae6ޖ{�QB*"(��ڌK���i4я���F����sܻnaiM���SO�=n�a��:���������cI��x��O2����(�����W�O�饗�Pu�$��{X�z�K�^�e����Ϫ�7e3�ڀ���'��3���%+�~�YY�oUn߾%����=z\���!\��=�fUU�h�i�w��d����@5�ړ�q�"�OD��DE����e+�I�!��tvGA��";�����CYԶ�F|nfFF��oBXW��sT��ɕ�cc#�cb�_�.�"	7U�$��>��{P^=�� �?�W��L�L��3��`X�	4`@��hf��[`��A'�w�B�[��nU{���
DHoT�9pˉ��u�X�)fymU�h�����J��uN5 �v~��e<�	L Ԅ��k����ϭ0|�ٶ/������b�f�>������4B�t�|�~�l��Ҙ�냛�Pu�`t��^�����D&� D�i$��"v"��H1�U��� ^L@dem��{@ʴ�4C�yTs�s2;;�ET���伷߽��c�N����Ȉ�.�$���ta�߹�v/-+ʝY��MlM�Ӛ����o�)�f\���J"c+���J���b�d�#l�G�>H�20��(�^Sg������섅�Mb\e#���%�7n1�73�:�5RK���'��[L%vtw�k��v9yv۵w��D)��^���������1���Bᩢ���W�Fs��?{U�\���Q�on�?~������P0����¥�Q	�/}�� ��T��_��>x������� �_�Bo|ey��g����2�c"[%"���O���G�r`���ԆZ
�R�r��+�f/�����l�k���<�+�X\$O��F�f2Q��ivMA�rj��+1�� .��4Jz��+��K��h��z��_	��0n����0����=�p%)p#�W.�1�N�D#�v	6�ȼ"� ����#!�����0�eBQD���Ί?�6S��Y۹d��!��+k�.jj��Rbi���!�,\`�@̞��ĸ��H�!��&X�ݹ3$�	����k ���<�˄�^i��M��aN�F�Cp���!T�6"�j�t�2���-1L�;�I4@!�)5}�ESdύ�I��.�D�^ڊ]$&\Dj���j�<�X�T���J�JΓ2��a�}��{�=�G/Rf�cO�DlN�]!5n
���,��,S�&�Ԫh�$ �Aɳ�,J�Ƙډ���5�Fv�4�� ���)x@Ͱ����U��-��&�e=��ҧj
_B�%aG�> �x�#����t"l3n�y8,B4����ƹD������N����f5;7�MB��\�;��&�f*�S�e���lK���w [Qiim��Ʃ��� L��v��Ԙ���ϊI�����?�����1��9�ԉBi<��S'9��\t-�{ɔ/=tV�zJ��9����~%�*%�͉<S7����]�̜t?̽[��8\o�����-���F!�2���?}�.����hk����>���ƭPn.3e�S���#� f��&�&��n~���E��7�c��2�����B؟�iJ�/~񋔚�^{�ja议=�����#�h����ʢ���țj�/]z�j���O�&!�?�+L���=r�����>�7�����	!��m��c���f�OAa����4>����>��?�O������!����R;��Q��N�¡�a�N7, Q)&~`�=�ru��� ��g���C��_�[�kTE���Ql�OybB/���R�g�����(UQ5�x����[[[қY�JŌ>������-3����,����$����9�\���,���O�M����nAN�<�}����ɽ�ޫ>��L �"��NK��#�zN�{�ul��Hn7��QV���{�]>+���G堺 ǎb\������{��TR&'��^fU�Oq�����2��bP���A8 W�^�$ �����G�;��xb�Dd�PƳ�h���!�Dc1"�J��+C%����~J�{�ܼ��l*\�����#��f9t�B��������GsK�؜<�������a����H�^���(U������{A	��&S����F������hR?aQzz:"�d7՗��k�0T��ө��Vx~B�:Gbp��JA<�M�?���P �����/��T]$���<��CT�##���]�����19qꀪ�Vi��&V�juU�˺6EEO�*Ec��S;���[�ף�-�T3��P�ة�
Qo�,���8<<���+O�bw�8���ș��rRԄ����c����c6��+$���PR��No���5�e�	�Ѳ[ ����xT�I��O�dF%tie��7?7#��핼�)i%l[K�ܼ~��[P/��*A�T��@�ޕ�m���~e$5��,-̨�,)4V��j�e�j��޸�:3z�>߼}S��K��6�� �z�y�Ԩ��J*�n=|h�<��Yy�7�#�u$��:Fk �7>n�R8}&L�d����Un���-�c �:/����)1q����8W���;
	7%�j�X}�cY	����k�n��u�g?��I�p�*�}r�@���_g�����J�s
�R�V8����:�G�dk�7r'L_f̓�I����[��+����m�v���*2w�{zd`_�t��S��='mm��������*�Ӵ��zX�S$`�@y�D�2-�#$����G�J^��kcjS|>@m���Ŭ,./�(���Ʋ��\]y��;t�{܂�\�� 3y,)��lMD�{����Joo1*�4m4�@��̭)I|��32;�&���o�|������%�7?>:��aIf�i�"J�Y��?��tw���G�B~���S�꽪.���L�V.8�{X%�K��0�[$�w�~9|�L��u�Q|�~X�{�HK��+#���چ�����0��Tk�(�m*"}�L�ɕ��jni�=D���i�L�͓r�����C�@�΀Ѱ��>�<���a�TY��5�W��@*~rb�g{��䱬F~��Cі�`�f�)��܌Ik��8�ݝ*��$����� ���E."�z�N!h�����5i�o�s�*A�'���J$��jm�R`Р^���/ǐ:��9d�lcW�<��ۣvU��pȰ��C���}��������cO}̌g�U3�����%��1�2�T��*���߾��4�
4�sC1���b�"PUP.r�HE�L�t�&�!�oz��ZD�+� W���������ŘYȍ��P9`#���5��
�C+�#�Tf
�:��~vn�����ъ,����_RuSgƚ�7�7�E5��_h�Ιwo1�����z\}����!�k ��i%V"�&q�|�����cx'��B�ZF,j��Em��oQ���e��U%�p�οv^

maS�<�Çss�0C�Rg������Tc����������~m5�j?ǝ��劭��V��& �~���aj�ȘZ.3_	��-��!&n�n�B� �]LL����A}�5u��L�N3h�I���?R�@E�3
C��sj��-��ܨ�=%�w)!k�M��اP�(����*��ݪJ��P{096M� �ުhmcu���H@����=��d�F1�F%��w� �����.[����g�tN϶`1Qiz��a&�N?���k�_�f0)<^Z</�j�==}fh}�b� ��;�%����$�:ۙ4�0j�6���}�j�����վ�;2#J[�*��Ӫ���uYY�c�MgW���uI���zէ_��?����u���������S�|��W�)�ۚ$�(iU>����.��lϚ�v�0�����T[ {W)aY�d��e}i�)��zR��^�*�j�����E��-��hRa�~%^Y��u��"��<u�>��SG{�B5! y��1u���Vo�3i���p3�4Ȍ��^�Z�� L7S�M���T��-��>@��R�СԵХ�j�W�"���Oɧ?�YUQ���/���m�7�Ӷl$ 7�Q�q_��r�a�Ƙt�����"��}�IHLSc�l�1�*�U�=�X"٨���'N(��}�~��?~�����@U���[@����*���AY_^g��z6�)j��9��zJ��+Ǯk�{z����V�~gB~����n�E��m�=�Nc
���3t�/�ȿ��o+ 8��̞ Qvb��H��O�X�M)]���?�fe��J\lѐC毩��CH���Ӏwao���2�882����m�zPS;���TK�m�4p3���y6t4Il�A�����WoS�ns~FR-���'�U�hV��,�O��}��&������%3� ��%} d��l��O6�A��|�J�6UUл��	9��	t�0����_�=~\豳3
FԐe��C�L&����4H頾��6�Pp;�f�T����'���
�F&�:ųs�L	 x���*�ҐM�jw�o`��Ʀ1��@ܜ��CA6�7��Q�F�%��tl��@Y�~�}�"x�#�#��R|��s�� �����·B\ַTElU�a����{�_%P�us�C)��,�[������\GҨ���x�KW��bJ8l������W�U����l*����!ڗ��1��ް0�`��	n��z&�5cq��A���?}�4�K�qLu���(A"4��z�c��Θjz�Ӛ�3�	����Oˏ��%�/ b`mm��wq�sGf�����%z�9�b�� �b�>�[�p�ϟ�۷��FrS鷥z1+滱�+�*�;�ٶ��7�K�L� 0�����<%�-�ŤvuN(������6ߎ�F���(m��9,T����x�K,�i�5E�׶��m��:�L�Y��������3� ��Ls�[:,ŁM�۲W���3������=��cDx��J���fy������]����x&7L��X���Ht`���@���yZ<�:���O�:Ty��;3.~īو� �D��{o��n1�FF�t�!)&��J�H:�03�]�������,����
�C����[���.Ĉ���V���4�qyA�"6�
G쎔�AU���Ѕ"=p񀪛#G���Ҳ^�U��)�z���]�~c��ŋ6��������]��U�[�g?��yJ��l_'�EAz I܏����A��Eͦ�'Og����kT(i�7M5y��u*���#���M��QC�@3��LcmSb(iֲMˢ �-@�]7�ŋo(���\��>C�_����7oޔa��oM��c9~ ��#����uӚ6.����I��1��s;!�A�  &`$����}N��d}�3�a�+�����d�u&����W��5)��4�k�mE�DF�-�ǵI�FTM#!�b���2E��'Sgi�qt�����%��?����� øi�qj�7��3%�)5�̪�#,�����������گ|�+����5��x��'�9���7�>v��g��)y������6�8wC�ڎeu:�uCUj��(ۡP3�i@�A2ٴ��0���z\����G"O@�mUMZa�#��Ɩ�)n�ei���`�!��0�D�� �k�CD�x�r9B��c�R�LM�ˍ�eb|Z�,%fr��P7`���d$W�^�B" �@DQ���@�-����-1�F��3gv�s~��OR%�z��(��'<e��1N��������&UF�V�ls�5��)��c��9�vHcm?9�^������l�����������߫Zq8�\�6��.�8��L�3-jB�F4���D̀2����d�^����'&��D?A��B��U*��D,��:�n�����0�Q��~�?p�[o���������P��)�կ�b.�NUÙ3�8�u@!߻�^�˗���D>��eF-��`�����o~�a����	K}���{z��S�:�3<2�D[�0hA��c���!��1f�244$n*C�l��g���})EY'6�D��A��U؂V����<�i�O	l%a��C0j����R3��,�tnRxyd`/8��V�E5�&���W�A���)ߡ�~�һ�v��.]e;�E�\sk��s���W���[�+P���(e�[�d]��Jhj?�uY\����g|�'�p���������w�b3Ҥ-�-l����>mA��$)�J}`t.}�S�!�~�Yֲ�����U7���k���Ԑ�/���J`28x��j����ɬp։/u
H�F�H�2�f��u������鵕�%���/�?�<�����ӹ۫j-�*�}����1�7�0˖�L�>2�8TmҨXD ���M�>��Ӻ`CD�2eq!�5$���w��.V�����L�(�ؠ���ׯ_U0�H&�&�ϰ����2T������r�S�8P�5�WlD�L���ަ�E��A�z7�յ�NC C]T��{�r1���D.�C��/r�F������[%p|b\.���������'�(.Ξ=����8����rP8�8'�$�=�����u�)BXX1�@.�XŇ�6@�1��d(l9�w��B�"J�MT*���#Go�E���+�Ј{Ul3$rzf���pV�+�̳R#H'&Fɱ�����
PB"��J�+����@m���bH�Zd�ץK�H8����Ʉ#t�8�XfB	93�2���ƌ����YR�� `*� ��[X���k��~�8r�(5	@�[;�/�v[��� ������G]�z-$��2@�����-o�)�K!�>6�H�kC n �cp^w�ș�N,�Ç���/캮��}��u΍�h�n���!&ILey$�dISS.�?���*�k�/χ�<U#�RyJaF,���(�D�C�D""�h���	��{�z��Ϲ�5��Fv��Xhux��{��q��HWo\//_c8��/>�$
����e��F�~]m<L&wM�"OF��d4��3�	��s ��'��%��-^~�enHd���I��#����5��=V�u@=�>�|�L ]<CkS�2�����jrj�#h�&A8t6�(�����A��'�O^.s�32�i�,���ߝ�����,�ό@x�]L~b� 7Ɍ.����e����=Z^��y�<��q`���}�O��ݏ�UiI�UF�^����J*u�Qg�nv6>��t8p��o��J�c4� ��5#�EU�;q�/ ��p��6"6�>�)CE�҂���O���H��q�p�h
�qK���w��JO
���+ʫ���>����L��'A���f����1���@ce�y��$�Yn�^/��4�=�4L�>�	}��8�A2����3�e`
�5Dy��ٓ��-H��. 0q��9y�ט�Zi'sx׮_����sC��Rx�mφ��4���p���۷�~[�~���ڽ�x*�(8�]��@��|I�#mv�/���{@�8�ﶶV�!6�ic&��9.�p��}��p�3�Il����k��h�]��$�J��O�;j����-�R/��Q[U�0�![�h���Mꢙ2X�(C��3jO+t���?95��Aqi�G�����zz�ʏ�#����L��~`��,y&��' (8>��T-��}�����i2�d�&�{������*&�0�\�P��o`��15q �0AEֶu�'j_�}! ��f�<yd�<��c)J�$7V�޽y�{�Ο=��<u]@��'�����<>��J|�%�is\�S2nim�^���UͲq�v&P����u��.��7�+c��E�	A��#�w��Vy��3<��CJ�_��CWO�iC)_�R|A��Ԍ�@�Ԣ��ͰTD����fa��{�wog3	C�#.kjy�yN�����F\�2��P$Mq� 	��P3TSW%�c��F�[]}���7�cQ�6��ueC_АN��EzA��|�! �ߪ��#���p66`Mf�FCA4�l�W_y�Q3ao�Q�}q�G�L� p��ь䏀7�f���vq1[�}�Gŧ���Bl���͆YE➱ٖ��4����X��S8��@���^^���(�rh�ĉ��pE{��LI����[$9���-z�%eE+�3M�ؕq�.����>��ZG%�e�	�;'\�p<�����h����
{��\�)���g���n�5�:ه�s�LN�3s�ﻩ79ǹ���m�ϑ��!���"�N�~�1�D[8U^�a��IW�cɢ���	N��b��|�+rs�r�d�L4'���ӄ�N�O3�jh�Q+��:��촃�$���+t�I��J11֗���JK��jE�g׮=DE���;{� �n�fdȅ����q!Pc�`#���yv�<�y!m�M�D��``niFZ�W���}�fBL!��o��D��~�,�2�0|�B�Sd�/��7Tr������v��FeZl@L�]�Ο!� E`��ج������z�O�:��H�f������Q`���:�
�#u8@:lۺ�"�㓓zt��3@�����e|P�nn�S�	�_0�������4��H�Z[�4����v��3� ^D���C���wJks��Yii�������.��~\F�M�-=-!�Y�dǾP8�?%	��?��4��&�hx�;8
�k�tڰ<��n*��M���Lss3oD�(�#�������$�d��'�xJ�I�����^>���{��Ǧ�p�b,�G�D<\+�j$vC}�ܾ3*C�Ä��ׯ��a�S����{� �Wt���j%2a���>y��ރ�Ů����%�����\8yX*}Bv>�W�@�Έ=+3t
������2���9� sr��]������ޫ��"7 U7Ac����� �)���=�[�vo�BO�#!髮�#h���N�_�&|���c�1�j{?8x����ըe��%�d�&�i�e��'� �M����֓Ŵ)J�/�r��̈�+_�(�9�&8�i�OH
�jd����{I��d��k�9�'�E[$�ʒ��'ȩ3\��U��+|ѧqt8�R=z���j��b�q��}"	�
8vlf5-h� �AY!�a�� 3%0qȻvh>���̀�}��f��l�����B=�c\3�)hV���,��i� ��{f�0�c�ވ������O?%�5�mhhH��FS�^��;�rnb�h��e�]�*EA��7�ߖW�I:\��2M<����ҕ20<!�Kf�ЧP�"�WСJ�J%6c�?.��	OD�y�!���-�?m��FG�m�*�����Qsz���i�>8x�T���r�#%)4eH� #�'J�*���L%]!-�Zʁ�a[����>È<6h�S_]*��ܼ5���Am�P�T���s �?Ķ<������<.�T._���~Qs�@>'Ee�pNM�аB��9����c��z3�{�	�  -~FQ����ſ�_D�8����;^6l$�y�~�A�4�TO�C"	�\�6PjB�HK��ũ
r�p�v��R��Lro��3�>. �Z��Fa�sA�GK�\rچ�u�k��K����x���;���٪�s�<���������4�;�R���/M�r�H,����u�V@NC��u�
�n�)�7�_���	�g�j�^a����<`V��׾�e>S ��ÿ"`/�,e���r��G�m�?0?Lx'Ⱥ@`=paf��lP�߳g��pJh���o~�mjO�4��m�6��4mij�A�h��0��i�����f�T���5KhTֳy��]%��)�Ӄ�G���/F��X@�0�'���Dq�נ����0�xМ�_����u��w]
 �9�H]w�M��8�_��-��������,(Xꛢ��nM'�`nA�x&���{�����n�	�ds.t��f�ehz�9&:(� �����	�HfN��>׋��yT8�u�Vy�'Y�A��g?�� �� ���.r#�Z�0���^{"v��{�2�<sg��*T$��8YYc⬊Ě�˔.� ���}�p�}r,8R�{��4�7�Hm��#,�Rߪ�!+Mq���4Q6lY®߾}�4�l%r0�+rG�B:C�g���c���'�Z��*�כ.���f���2���8Q�e�2y��ȩ��M���,	V{�p����ň�g���d��0��	(<%~�M�Y��\\@��D*p��eM��p��U���c�ѓ�\�^�����7���8�o��V�2ǣ ��ט�H:�f��!AȦ=w�	BӢT1k1ԭ#;f�����>��0W&<�Yp�ԫ��,�$���=i���]�����$�X9r�d�+t��4�e�H�->At�.R�b����_u��h�ԯqNDb�w��[\��Zkv��,J��r�)G>�?mj�p��ʰ�u�W����_�cص��(
�5��K׸{��)�E��-\v�	�#�<�\ 2�)o=
oЗC��F�
�Q�131&C��	����2x�_���Y���8eY�� ȟH�+s�����
�YX�/oV�9��{�	4���	�T��$C:#�j�K5�wF��L�L3�ĉ��)����}�:��ȝ�}���8K�Aγ�B���C�DFI�L����|�%��L�H��l�t!K� ����Ō+�� ��+��䇧eaf\�*�k�Z)�(��gNH�T D�;۞j������<�C-Jܢ�M���g�W�����/�?--͚O�'���� ��U�$r/���� ��b]����;5)C#oq�Z�c��m��e��r�ՄO�ga��03 A�mXOc�q�I�eJ�\���ś�1�<��dܰe�� m<m�L�W�;ijL�kg�Ͽ�C����5�j�&�Ϝ�����(o�=��Ф�v��ro������(���ifx�0�*ڠ$:���x�C �D��k��&M�|��j���g;��2딎���?�5�:tjCxx�xͼ@N�8�^3�pJ���燊/�!��Y}C�f��
�$2��@Ӽ�<)#Ccd��+VG��4���,�3B3�i�c}7�9(n��c�y�L���y��s0��ī��E�7�$6?QdY�EYfƊ4W0�lJ]&�� >��<����bZ >E��DO�����5A4bD��B6� ;�2�w�l������1����O I*k��~E��G�4���"p��	'���~�n��;7;-Wz�P^��P4B��SY�Pc>�`޴ ��y3�F¨�4�#+8�E�k\ZX�/�Ƴ��2�nkj�چj�
��M�NEY	����Ѝ��v6��� e�)H�A;G��廃�C�۶藍!�ҥ��d���r���5�uKM�M�f�(����#��,�\�
i��@P�#5b��U�̧?���Y��Ґ��������e��$S9�P��Pg��|���Vl�D�B���Uc�|��h��x`p�<G��d���׾"k֭���7����!p}]��餥���Q'��pR�1���+ngfv�į@�H��b9��~B`��E5C���ֻB2.��s/s��rәrs�A��T� �Ͼ�b����u�{wo������Ț���>+ǎ� `@@��(�qZIA8����1(�,|E�r�_�����,�wj%�L8p�>J�4%��6G�>�P:�W����c~�Z]�]r��]2P#2D(��Wd*Y(��"[��S��4�p'V%	m��SE�`� ]�,����q�Ӵ�Yx�y�d:DP"O<�$s7H���{հ��g�gV;<t���\.�@���/j:�^�y�\���(��V:��N�'ԟ4"�s>@܂���e��i6�n�C���h̝>s��������)�Gy�C������@�B� �7��OB#�Bb8�Iё�u ���ݭ���	&{pxe�U�9O[#�8��+�	͔�;A��͍ֳ�?66,Օ���֪ы~�r��L+��s����񾈇�`�	e_��L�ݜ2���a���6��a��V0��1SL&K�Ѫ��0����t�t��M[���ӼF�_AG�r�E0ڦ�G��IʴECNr�W�i���{�MuD4��֓���ƕ��|#&p�����9W��'�'"���S~���i�����}phL~��7�f � e6��3�_�L����Y"1 ���::G���=Fm� |���<	pK�Ս��e0=��-+-�xq	]ԙe�2�1-劓�;�����9#e����Uu��s/HK[��IE;{ĔP�����wFX��$���K��'<8h��i0L���<�m�N��$l@�mo�(!��@a?�L�c���{��?)~7G��B�\)8G��o�w\�K�efn������>�Y���Eq�dsح�.���Fї��u��![^\���d��E���=�{�R8�hU���Ǥ)���?|G{�T����-�H{�N�8�zO�A�C���sa�Ӻ�Ġ!t��0�<�3p�s�&g�1p#;v� ������
�S�oxavT'm�r4x�I�/��M_���$J���]��9tXT"{�<JS�D�Ƚ�a�~)�}w�9���T�OD����^��rY��@��SO3k����U���Z�$���E���4�rK1a��aX�'/e1p�&|��!V ٣�G�I����h44�Ǽ���P'�*|O�� �	Ȃ^Rx�	����T���'��$+;b�svI`�~�
�T6	�����O����Cnξ�x�Q�����U5�w�^�|��a#:��4��u�2y߸k�N
��ٹF��߾G-n�?�ן��SrR��� �L38�ضCΟ�(�����\��]�\�EK�S��g�f��%���G�pw��-#}�%Q(2p��ϔ�a��QdR~@N�ß^='/�K�2��7�T �i$c����GofU�Y�Z.^:�9�1́���	�.]te��O�0��>� mm��5J.���.2r�nWw�����(J��:+��u�UtrZ�_q	�L�a����ӷ֫�Q	gd�ܸq��Q(������i�n��$DV ��JF��Vy�7�3:��EM�*��`F<��í�|�*����z��3C��VL��6�҄�%t�DnrB+)�� D�;J航p��)�w�YP�$=ji���QO=�I6��@2�N������#l��;����0u�E)7�����I%�o�!r�r/��Z����B���I�LZ�Zk�WvKsG�.�.y���x=��%��7�\ȡ>��9�Q�-��w�ʣ��M�z�A~�W/�_��kh�'��i�u;v����lݴI��{Ɖ�གྷ,)q�������l��	������F����L%�b0v6�����u�L���^����H��0=۷o��8|���0����d�s�}I����d��+�����f���6N�0p~��cc8����_���1���-���J]���L�Y]۽V���b>����|���0�	,<`�����@��5)�*˙ۀM�8c�0���}�ߵKΞ;G�~ 44��c�=*���y���j&��p��s�ۻ"c�Mf� a�@��`-�ȅ���g#� ��ʢ��B�����NSYv8<( 	E�mp�O��^�rQC�M�H?�x���źc�D��8q��QC�*�%��=vT�n��#_�r��҄����9��kNA�PZjd�^�f�����x�/^��Z�b&g������$ӓr��e���Y:���vǠ�p��q~,&S��ְ��?"m ݘ!N%�	c�e�.�6�%��M�J5�P,$�=s́{�����*Z���u·�ǜ���a�"��[�͹m�,#>�\���Äx�7Aʫ��)-��!X	���(T�,��b������d�5VQ�`���X�ij��GYe=�6���u��r���]��qP(�t���Hli~��Z�f��:�V��J5	+fug��f�KL!�Yo�Qe��dʙ�����R*�5xo��pW��ٴ�{n��&�q���Ȕ�H��@6�aV��rtC�+�6��'C��w��x)�(�1���PC$.�c��'H�L#��4ìr�����x3&^�uD� ,��S)#pKa�b�V�g�t��	
��$���w��]��v"X��I:�`!-c|΄+�r�h6�x���3�D�?�y8�����D��k��a�����L�\�_!N�+��vc6���
��`������F�S�,P~�#�J���H
u$&HQ���b������u�Օ1��fM�`F7sݕ�7`��B��#M ��$l�,��9}�Z��
,Ykڬ��8,�Ü�Q�e)"L7(N�]�E�\d����A	��|�*�L��j�%����?C�XU��긯��X���;2�w�4���&錇���G�MF����yS�����fQ���� N�p1�8$9�.X��a��oj����&�q-1�+c��JD>���BV�`���
$����ZJ��Q\bg���4]��۹`{~T��$*��N�'�g?��{	�3���`7p�>��+�aŠ:?Z��6_��5'_��7\|�9�g�5��n�/~��TF^v}�G?$�@	��Ⱥ!��i�Y�&�I��Z�< N����7���sj��H������A^����~�V@7�N#��Y���#��0U<Qb2׾����;7ZRz;��&|U���$�����W��u���r�!��߽�Tw�ϻ�-O��˂}�1�O8����m���R�%}���,ՎQƾ�(Ñ�{�GQ����	EO��a�eTD���y�� �P!2��Ƨ���ی>0��DK3� ���q���/&��kh�cN�ȅ�`��ed�N�r�31�yF_$j�л�RCc��.�?]���Ϩ.
C��f&��nAf(��#�����<�h��B�)$-��^���|EA����5p�� @���8K΋^ͶA�V(��Ɓ�+�|a��G���L9���g��xF�L[��w�>���#��w�~Gp��A  ���<���Y
N�<N����#B��������3��2گ!)���<�p=׋ݹc?�'N��#G�R��#d��5U����,���9��=# 6��D���Q��� �. ��K�/f��������q&̇�Ŵ�n�u]���2���Сc�'D �vAw�rnI._��&e��h�{G˚3I�p�%E��?wv�K__/f�葃d�A�v�:>\�9YҘ#	�BnNC�yj��!bC� G��-���Z�5Lm&��j��3`��L������d.�<�R�t�!ԅy�;�o�aM����"I�O=I|�jq1��:�Ml&!?m4��F2\X#��h�\��#�:b�I`�;;Z�aݕ������Y�Zv�y�T�o��ݷ�`8��#��s��΂�����UZR$۷m�E�����i����S'�0zq���4�ȴ�J�n�鲢*
�<r��}���s�Ik����CŔ�D��]:jl��~F	�����ٹ�a�Gg>"��'�M��kzr��`:TfU����(@�F�3Ӆh������ψŕ�r�%��l����'�?"[�ۥD��'7h"�ʞ��g ��-&Nc��Z�Y?u^����&Q�_a�1G��S'Nh�|Ym�u��׭�|�2�i	fQ�,�z��l� U�t���Mu��$�RB�P� ׀�<}&(�4Ԕir���u��^OnE�HB]ȭ��T�X]f��K�$�!��<4?h97m���&�����l��X�� �?6E~���}���Rz*:�[��Y�,W�i�]]ۍ:ϒL5C��Uu�e�F�C���{�F>h��dI�����}�_�R���o+("1D"�$&�T��~���̬��W�Sʌn���d��D�E��HV'�x����$1`B@a�/H�֯]#@Ц�x��[�aR0H#�����gdljF<�g�8� � KQN<������*n{�"f4�����S,�&|�B�{<6�W
���
*=��C�庐�S�����b�AEY��9��m�]��T�ū��|�4��P�K��F��1["�u��9�����Egx��/�%�3v$�AzZ�	`إ!/�)�P�dA/�YD>��ڴV5r�B2&��I�)�	�((3��7Q7P�� "�f���SY��/Q\���X�����I��:�e���]��UP�!�C�������z�ۈ����CC��K'I����9t���]�ɬ�R�Ͷ�49��:<#���&�x�1��(�빻B���pJ3E�QS��>c ��Q�>���4��IZ��;{�vqp�'�� �:�Y�-�I2"�	��'`9^��0��j �63���|V�����\��dsÚ�j�YN��7<��X�źq�2|64��{�Q �JN,��sD�B	ۿ�uv�ˋ�='��la��P�����?`��C���G�˵�A��R�9��'�БS�ؾ��k��6���EΨ-��@!	�O�ߧM<
u ��cI"��w�� Mͫ�p�:m 3�thv�g�(�݈]�~jZ��Y\����EU,Ћhz�Z�'ʢ���&5���F����rs�����Q�
 �˦�}VM���<%��K�g�wB��m�����9s� �尶(��O�Y��4ʗ��5A�XY�L�Jv��If5󫽗� (2��X$iY�Rag��V��2�4SLm�k�O�I�sJ�����T��u��+�P!�5E��f��VW��%�Ikt���~�s��n�<�������(ǎ����N"u%w9`4[5/B�x\���Z�؀��"c!�N.4Ğ�51s �/J�'=�����/}�}���ac�RC�-�7IͿ�����w9w�E����T�)*�UU�2�l�D.�$B�!�K������K/�$����ka1�J̲O����X��LK����{r��myd�*-OOf5R��x�����B���.��8Z.�$�f�%i�c�bd:�A�Vo��˾�ۤ������x�D��'��P���I��*�|Ry�Ʌ� �X��C�z�	)�wm,2X����S^|�y�ڧ�is-,z�AX
8��kȗ�ᖕ �o��c5��X�T�P��	&�P�"#%Y���!k<�ʲ*R=lذ��s��5}j$������F� �B:�m���84v�7_��B�?qM��I@�����J������TQG�Jмbl.�4��)'�5�)Kk��a8�itsS�ɤ8?R?�5��[�Imu�^��(	�m��<�9���[Ni�"��������P��)��xA����:���3)�Jk�*�N=��jQ�jWiL_K���3xg@Z�Z�[�lټE�N��M/�fP�~�Hx.Ԋ�HL��������N��711A�:�O;״�d����B��Kp�ص eA	����P���,e�\����{���OS���$%�j+��1�"���(taP�!�&p�U�<�h	 �9u�,-�G
v2Y������,
�h��c
��E $�'4r�D3u��>����5�N��d`t�%v2r��AP��}��4NNL�%Nu���F�T���뿕�=��/�C�������O����֟�;���O��?�)����� �̩���@&���I�	��l��^�c[���1m)!����Jo�HS�6��1���f;�HL���ߡڀ�*�6C��ٲ��d��UVɌ�1ZZq"�)��3S{�c[��M?f�*�&���E#��t��{\�  s��$�Lj��̡�75�L[�X`'o�+������Ӓq���HQ�׼e.K�tx�&�U,Z�M�4� �	>�XߣI}�ר4��׍s��*��]��+�|�R�\h�$���5X��9P����!�T �#]�N����NTD$SJ��Ҍ�����}��cj/1ʵ��>ᄞ�<�ǎ'����{dh��na=e	㡅�"G�rr�j�l��t����two��Ҩ�$F��K�dE�M�.c��;��ʊ:��7�}�d�*�q��� a�߹(>��V�S��- K��ڗ�����y�lh�}�[}7���~G^z���,H�]gO	������C�o��wu��{���]m1��{�]��뿔��v��5̘Y�ӕ��;�$��nVH�߹K�X8�2�6�����V��h]7d�p� 6�G�c��F�z�&#����J�$�r3����㿵�ȗ�m�U����8[IZO쒼w����	��1�:6:,?���Z9�H�9BUg����J� k�>���YJ�srC��f��I9������31>��'�!D�zA����,T��pA&�����C���oꢖH�+_�������;�~sD�����AihX�^BS]L!���&�d�����(ܾs�6��$d��H�*#=�vɹ����������v���x��>��44j�RI�4hPu�2EI���R_�%N����n�kO��*�_ WWZV�'��8"u�у��٤N���V�E�>#(�rB&�Yo�{G7Fw;ƌ1��6�˯����� �&�T��##��{�)��D��B,��߼��n�����l���O�an�m۶���?ee�׿����*J��q��4Of�i���(UJ��<��Q��5¸��G�����H <Y
�t�{s3�+z�������зDf0_M��i�ȔZwN��B�Q p�K7�}C�#*��z͎�o�.u����9G�
H�������7�^���K�j�p,L����2#�[�b����Cz���݁{d�a�,_`���}����@%�
=�ϩ��A��O��|��_�)4(����.����)���?����Kj�n�2ŢLOM]��T`�k4V�P	�r��G�;eef���M@͉����E��-��d,^�7o�o}�[��ɩ�l싃,i
���S��QZ^�9J�)8�jԎX�
�K�g��p_���ѓP��4]}o��ah���I�Fu�w��� ~�f�&����o�4��p�%����;�zS��64�5a���R�,� qê6ijI�W����Bx�2�XDs��/�K�s�dK�͕������gn9����y[�\M���8#&6)���cQQ�Dl��<O(�:Q��5�K]cK��8Z%Z5�B�L;����-6������&�
����ϸx�&^;eߣ�����=�=��oC�CtD��~F�A�!�B�Ĕ�:��aP���~�~�&�iǇ[ �I��૩�����{YN3����J���Q٢)���!���j��6��Dk�$�LYi�qV8����nLM�;�+]z�*�w�}���)^����䷿�����󷢇�TV$hh�\Q��ֺ�������yd��s�c\���0��e�,���d���.��<�9�=uumd5?KkVr��P_}x�}?���
in�����^�~��R�;_����'����ߥa{�_YF߽a#�.t�����+,�G�M>�	��b����~�L�;�R4�Y�t�[�(f�>KSs+�M�m��_���+���=������b����vٿ�e���;�3�)��X�('=���z]��a�o����Sy�^!��<�:�CݰeA������������?�Y�W'#�-���xy����/4Gź{Ke����Xk�����;�(��~��*)=�M�Ү�;��E    IEND�B`�PK
     ˡ�Z��n GV GV /   images/5a738b76-89aa-4728-b8e5-f09c859dbb14.png�PNG

   IHDR  �  "   �?��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ��IDATx���|w���������j�dɲ,˽�v�$!q��;:� �H.wGr$��B�����s)$�@(C��;.�w˖l�����&�Ųg������gƊ�7kiFZ�|������LB                 d�]                 � �                ��@�                ��                rw                @N �                �	�                9��;                 'p                ��                ��@�                ��                rw                @N �                �	�                9��;                 'pϲ�Sgj�vړ�&���{�����4��oxL���E               ��s9l��n�ץ|�C�M���>'����"�Dc�h`$�a��	!�����"�^՗jz�PUE>�#���B��������7���aI.ۺ����_{���w($               `���/�kz�@5e���nE�/���8�?2�=8����ݎޑ��j�$��&�Mf�-5�j�-֜䲱�/��a�~v�����2��֖=�z�[;���               �Dg4�6��sj�S���ӊT�e_����0�����}ښ���h���T'���	2:�7V��tf��55;y�oWv��\Z�\��P$�W�Ն7�j����               �(�|��Ơ�5�k�2x�Y}=F��Y�E�q��7?ftvqg�6�qD��w+�A�� �~��:��Jo[P��"�r��a��Ը�]���~��~��ں�               �#ľ��\�ϩ���rٲ݅�/�,H��:u���"z~{{*�k�	�;��P���;���u�*��DU[V��i�fm;أ�lث�li�X8&                [�������u�P{�g���<�Cg/�I���~��~���T�j�y܏���]��A+�+e��gɟ0{ZQj|��yzr�A���]j뢫;               2'��҅�R����ݚL
}.]rrcjl�߭G^ح��R,��/���c?mN��&���&;�ۡ�'���e�S�!<��.m��%                ]j�
t��3���5rح�����Ƒ�=��.���}G��A��X-��R���E�J�4����+S�xB�_�ܦM{;               ���4_�9�IgͯI5��j�~�>~�<��Yz��z�]��ϊY���-�++�|B�+9U/�qD��|��t�               8^�]vv�޶`j��P�ש�٬w-��������{�'4�pO2:���y:if��-kjɌ2�j�A���f��               +�ݪ�V��{Ϙ%���*�w��w-Ѕ�g�'^�;:4UM���鲷�$��x�ϲZ,:{AM�����E�oث��~8               ��ȟ^w��z�?�h�}��W�����oT�����)p�_W�.\���A�c��v�,�����ˏ����               �����Gϙ�j���Y�\�Ee��u��g�P|
u��rw�Ӯ�ϛ�s�	�oNm������Γ[��s���              ��9}N�>q�x���q;m��s���\�{�%��T0��M��|�RUӵ�N�M;g��7U$O��               �.�æ��>G�h�1��D߾�,}���䦃��D��b�.Y٨��1Gv�E0���R�w�Y�����Ү#              ��3=X��w/Wu	ͨ��s;tӥK���L_{|��&�Ip�8�q�"�1�ZH�B�K������3;��_lU<�               ��U�uㅋ�vڄ�9gq�+���|A�#��&u��<���_���!��N�}�LU�鮇6h,<y�              �d�Xt�;��ғ�̘Q�׷>v�>���ڸ�S�ͤ�Ϫ.���[�@�KȬSfW��W�����9u�
               ���a�?\�Xg̭2�����?x����+�ū4�Lʀ��͕�ǵK�r0�A�ԗ꟯<]7��s�t@               �<�>��x��TSjd��f��_�D����ׯk��t�3�M�'/Y"��"dW���?_a�ܟ��{              ���(߭/~�Օ�e�H<�Y�<����M�'��&U���%u��ꅲZr?�>4I��;24���{b1�`4�*֙�[{��j���[��-�|��Z���k�y�������v��|�C���)��ߞՖ��              ��e4@��GNUE��\���50����	�ĎF��X<�O$�c�x_"a�U"^�t�J���mV[�Ӯ"��Y��9+�
�~�˪w��z٭V}��W'|�}�܍o�u�/P.f���Q�92���;��p�H�w]{����ښ����v���@��꒼y��y�ֽ����<E��g�              LPF���.?Me�e.:�=j���=0���ѱ_������GN��w?:��?3��:���s��`ae�י[�ݤs���f��?|I9�>)��XT�kϟ�S���]�c{����	=��}׌����Z���so�ۍ��|��*<��U���k���s�Ż�iӝ8Y7~�)�<�'               L%}�ç�T�}$M�~�g���������������|��&�{k�u�:{�՞��|���N�Q^Phɑ �;�h4��ߤ�j��O�S��,V.4-��7��ڲ����_������k��w�'��0N��k+��5O+��rز�U2:��'���<��G              ��W�s�:YU�y�~)�'��m�ݻ;�w`���Z�ӕ��кjU4���[C��?��$�w[Su��r�ש,�py��"1���-��&t�}nm�>yq�����z{�'�?�v(r׃�k��o�<_5���?8�wͫ/~oe�����w�V��{���1               w96����-+���	�_z�ȓG�F�.]�ڏW���\�=��͇/����2zi�5�]���ԙ��գ/��D3a�E>}��S'M�lo���v�����r���qw^��HrqY�uW:7��ܚ��낅�l���߫;޿R��)���              @�1��7^�Hsj�������v�����|���wk�֏_���������O�-��������;_}�|��s��k"���|�C����*�R�-��;^?��mW�~P�[]�oimM|zcՏn]�P������L���J�n�t�n���H      &0z�x�	y�q��	���.krݦ�H���O}�1+����vKBV�  8nƵ�p���蛿n�K�B�aU8&�Ƭ���,�u��"�Ԕ�      �M>k�Κ?-+���m�u�?��?�z��!M0w\s�S�ł�o>�����;Kggg���q?���^w�o���_ń��؛�_�⼌ﻳ4����w�r��VMp���;��������+=�zZK�{�.{FϚ��z����      �ƪ�
�	�b*�Ǖ���Hȗ\7�5{3] 0nF�}4j�pĢ!c�����V����&��     �-+�+���ge|��xB/�hߴ�;|�;��&�֏_�Br�r�=�����냅��ܿ�i���[��~��	k"�p��٬�f�gt��x\vtlڹ��_����jy����o����8�6�Ȣ��zK��`���ơ>���!      �>�5�wLW\~gL���#� �4ޜ}$�R�b���F,�[���7����B�      H���<}�%�p�q�?:8�򮎫?}�E��$s�G/�Akk��u?��)�+/��82v�+���Sk���{fB̨8��g��g4et�:G��Кۯ�������%�%���#7��Ss{�ϙ�����o� ��O�k`L      SY�=�2OTE��J=��2&�� ��+�|�1���Q�z�6��sԦ��z,.      ��鰩�=��se.f�ƴn�����׭��I{�筿�U7}���Λ^��9�%�L���a�թ3�_O�T��0�|�C7�Y�
Dg�˻��ٴ�{�WoXۣ)����u��xlac����L�����k����<�xb<     `�cm�7�
cxbrڸ6 �_�'Te����f�=���sԪ��'���]<"     pܮ8�EӃ�_��h����W�z���q׵�lomMT�}���V�q�2����ok�ƽ]z�`nG�'L���ՋTV��ȾFB�ĺ����_p�����[�-yҔ�y��Us����C��Jt��3��3o     `��Z��'�
�Wzc*t�  N�͒Py���1*����wa��Q�B1��      ����fŌ��o���/�?���׼w������_t�}�����U�)-�8ҽO�բ�/]�������V�������9U�WG�p���G�q�ի�i
{�9���~�w,���㴧���eok�;:t�sP      ��E	���ɋhzAT.뤝U ���'�PI�D�7qרU���7��aw     �?����/Z��EV<�Я7|���w���ۮ\��#_����/Ϭ
ҽ��"�.;�E�x|�rU��}.}��y�����#�nm[jt0Rn�|�]�{9�΅5�+�:�:���nM�`\����m�     �Detj7����EU��i�Z  ِz��K�E%!���t`ȡ�a:�     ��+�1W%��'��|�>t��Bʗ�]����jFñm�LK��V�T��lnӖ���E9p��y*�:Ӿ���z{_��?����~�g?��?��x�����O�޴N�<�H$O�G_�-     ����WCA89�r��� @.�*�*o45�	���ƀS#F��     `j�=�H�-�K�~��Q��}��rŚ�
����C��>0#�5z������ܗ�b��^�HW��+E��wO+���t漴?��M{��v�u6ߑ<0�?�k.~*q�#�N�]�|uI^Z�1�=0�
�	      �٬R�7�Ƃ�ʽ���׭�n������~v�M��^O~�� ��y5�����n�XF����y��Z�͋��pԪ}�v��w��     ��բ�]�(zN���p◯��ȧ?zѿ
ԃ�k�J-���'�>}N�)��WMi�.Z1C?xz�rM�܍i�?~�ܴ�g{[oϮ��-��n�K�z�ƛ����3L�T�O_[}�ˮ��6[_y�U     �<G\�
ê/��iͽP�Vw�\�x<�3�n9���p8�a�[,D� '��G"��cccM�����rddD�P�5����j	����mخ�}.�	     `�8Y���
Һ�p4�'_;x��csͻ�9��~����%����Θ�'7P���rI��ߵ�^��i��ގ��W�zg�y����u�%�w?�γW=�������%uz|�^�<�'     �\R슩�V]^$դ!ی�yyy���W�ϧ��2?�g�;��� �{l6[j���?�D"tJ�Ac98����Tg�l2~���ES�g̪��N�t(�\&     `��8�U�Һ�h<�������+�|S8f��>�eǯw,�Q6#]�����Y���G_Q.�ɀ��i��jN�>����zx�>���0.�]�z�힇���%���<��rUט��#oo�?|�Y     d�q�&/���Z�e�u����B��#� ��d L Ƭ!>�/5����>�������7G��z/rǵ�=�E�T����"q��     `�y�iM*���V߸�����+�|F��VK��{<�����<��4]�y��Z=��.�;�;��s2�~�I��d�����/|b��|����r�#��W4|ޚ�)���jnm�6��     @v$T�iAј���N����U\T$�ߟ��n�� L>�;�^UU��X,S����z{��ӣ��0>�I^GB�JB�����t     �GQ�[.oH�>~����7]v��q���G
���9�}_]Y�'�0r�F�۾��rE��=N�֞:3m�㉄�m9𩻮�d�pBn�j����w�>�zU��atq���O	      ����/
�ȕ� �ѡ=�����D%�ũn�  LU��Ţ@ 5���Sݾ��ݭ�.���f�ûӖм����°vt     �ĻO�)�Ö����t��qι�	���]t�{�c�z�u��rQ괖jͨة]�}�9p_��A�^g��?���3�\��.�]�oo�=2�:P���skK4��D��u	      ��Q-(	)��L���p���Le��*M�=�.� ��.���_�h��W$QWW��vv�ȑ#�F�i����3#�����~��	     L8�<�޵tz��w��6�m?�VK�ȝ�n�z�:����[:��t�7&~�M���F��[�[�:�����/��8[0M�Uћ����A�gs �mM�>.=���;     H�GL�KC��{���n�A�'GQQQ*�  ��xH���"5b�:;�q�HF��n[\KJ�4� �M=.�r     `"��9�Խ=O���_w�5�S0�'/�����~�����g���)�+UU��C�Cʶ�
��9�Z�����$^|���~xL0�]׭�����.\���t܌]�T���|�     �ٜF'�@HM��,J_V�՚
�WUV�:�j �<��~�#n�ݻ�t���T���s�8�:�|T3G#z�˭�PZz     ��i���e������CO�z���L�vp��꒡���<��V�E�h��ߤl˩��%'7���s�ۿ���Y��^��������JM��g��5���<��      �bUB́��BrX�l���Ju���s�r  ���PYYYYj�B!�wt�P[��ҶϠ'�s�iπC�t��t     ���5*���R��k0�y0�ZH�����}���n�,�}3͔�Y\���j�G#ʦ����RS���´��tp����j�������\v�Ϙ3�U�'^�H(�S�    �ɯ����2� �h�^W���< ��p�\���M���~8xP�JKWw��HCADվ�6v��ƀ㭏     ��է�n"��K��n��F�����ߚ�ȯnX<�l�ٵ]��6�F���[ٔ3��g��x�dyew���iu��\���������]��댹���K�     p��ք�B���"��|>��֦:�ӭ ��RXX���1��Qm�i���3}?.[B'���.?�;=���     䎙�~5&G:���s�-�_�U!�v�=7�}�Q�u��a��tpO��:cNUZj���c�W��!#��=���ʁ���
<f�>oIw     pܪ�ZZ2*���`{iI����U\\,  �ی������L+G�h���4}?AOL�N��^���8��;     ��jH=�&v�PȈ�?z���=��w,�}�ٵ��<�H��Q��D��Ԗ�TK{��#1�=2�>!c�N����ue�6����"Ք��@���    ���&��$��s'��X,*+-UCC����t:  �c�ZUYQ�]��ڹs����L݇͒Ђ�1��E�L�[}a��     +�բ��Ԑz���uw��E[��Y�w�C�_R�9̮}��i��u�����;�^�QȨ[�Xݺ�W��X[��3��i�c�?�m     ��(q�trpT���i5�`{Ey�f̘���< �����X%+V���v�RO��7��ΘΙ6�W�]��g�o��;     ȼ%�A�{���	E���.2�hJ}R�O�_���ڧ�T�?٤��#����=-j(3�n4W[��Ǆ��r��[�e�7�]��9��    �_dUBs���w���577+??_  `�Iݓ���رC�����6��/)S�7��z4%�     2봖�4�~e���_�v�^!�v��?���ݥ�S3�E�nͭ+զ��ʆ��W6W�n��^w�Ν�W^������?y���k���\f֝,PuI�ں�     ��8�:58��˼��~�_���TTT$  0�!��+��ѡ;wjddĴ�ިΫ�sn���:     0Eج�Tf�l�hL����⾫����?z���K̮}jK���/k�^3�Hh�ၿ�f�ZK����W�>�q�p     L�/���Q9��tm��|�5k��e��@  r��bQEE����<�7v�R86���ת�Qm�uhc�K	��     ���i���8L����[��K^��`��U����=NS;��#�}��p�Z��3̿9������/���UG�oG?�q�M�*�$y�����     �o%4�(�yEF�����6�U���jhh��j��  `�0���֪��2r߿��҉K�%V�;��;<��     �ϲ��	+����U_�amO�COn>�)8�̺U�y�,��pϰ2-����� N��������u_��=]syrϒ�3�.�^*�æp$&      ���*��s����>{�ly<  �7�á��ͪ����m����kJݠ'�s������l     H��i��}�{(�ُ��!�u|U
~���f���2ߔ:����KL�i��;�?%䄃�C�,����5]��*�ڼ�[     `j+v�tz���������2{�JJ̿f  &����X�\Ԏ;�DN��/�^��U�Z�����
     S���PC�������Z�	����-��*>S;�ϫ+�z���b�k�~����׼w��⍅��50�����-G�&O�     Lm��:�lD6�	��MKud���
  ����!j�֭���8�zV���lTgL/w�u��     �i���Ե3�	����3v����2�;�̚sk��z���-�7O�<:�_B�h]�*z��x�����̺-5�;     `��kqɘN�Z���ռ�sUTĵ  0~N�S�.T{{��nۦp8|�5��9^{\��*     �	KGC���w]s�z!gt�ޞ\�p/�w�"�S{�2)k���<xM킟z�{$�-!�t��(�05��\�Mg     �"��Ȓ�1�,<��]� �Y***T\\lZ7����|�a��ݫѨ���     ��3�:`z�C]/9�k.~�̧�G��^��u��M��{Cy��5v�|�ڵ{��2*�}�x�6�Մ���R�s������1    ���nM��QUz�'T��vk��*
�1  L]��ͽ��-��=��P�bWL�֯y51�     �zґ���<(�}��{���&3k�'��_�vP����{}:��C[��s���,��3����f֭/��k�Ļ�     ���&��bD�����4w�<9�6�   ����j��q�N����ۍ��a�zC��    ��z�*�w�Zs,U<�!�t��>�\�p/P�e-�>=h�_���'BNj���P^x��5��Ћ;	�    0�����FR]L���bь�566
   �|>�V�X��;vh߾}'T�mK��a�;�U�M      㑎��{�t�^�vH�9�C�{���ƽ1�L��%Y�W�Z/���X��m!'�FO.L�W�|    ����S�v�3~�5�^�.X����_|  S��j���f�~m޲E�h��k����o;�j!�     �ݴ�|�k���*��^{��S�Z�x�f�,-���)9����#k���gj�����;�����##�6�fy�+     0y�9�:�jD>��ۋ-\�P.�K   �PQQ�������>�:vkB�*���G���v�     L0�4d-��"/9�k`��"�0���>���@�2%+W�y.���v���r���^�lJ�6��<(���     �>{Bo;�p��i��2{v�{*  @6��|Z�b�^ݸQ]]]�]�jI���=��U!w     pґ��<#䬁����´���"yM�������Ccto�a�����Ӟ�)�7�Q�2�WV�E�DB     `�p��:�rDy�n7�F���  �
�á�K�h�Νڽg�qױZ�S�G��ݫ�sJ    ��'X�1�^,���J�Y��m��r3k�3)+w���)����;���=8�US�_cV=��"�ۡ�Ѱ     ����uvը
��n7�cK/V   @��X,jjj���Ֆ�[�8�&>6KB�ʇ���^��;     �ӊ�ݦ�����^�vH�Y�c����̬��3?���d�W��az͑Pl����G�{���B���;     ��Ӛ�Y�#�nw�\Z�t����  �ˌ�f<�^y�UE���a�JgT���C^u���     ��<���ݞ�P����:�kx�ʤ��������~!�E"�n�k�Nӫ    �LKu!�Q�����F�}�%r���B  �.%%%:i�2mx�%������a< X5������
     ��۬�������Bnk�1f4f4K:��NV�y�;�+�.!�E�	ӟ�1��"     �yƥ����*uǎk��߯�K����:  �X
�r�
��a�FFF���1Ϊ���ͫ�!w     �?|.�L�8����㻈��i]�*z�+n�ʹ�~Z��FV��!fKX�BNK(nz��ag�M     &��%c�ɋ׶eeeZ�p��V�\  `b�z�Z�|�^X�^����U#�ת�Q��ͫh���     `�r:��X��㻀��EL�;���攕��#���G����z̮�s�    ����֬�8�� �d�r�R!��/�������ө��m�W�      Ғ׍��CB�E�Fw)�Y�2ݐ:;w�CɉDB;��v
9-�v�]�I�    �	�6/�E%cǵ-�v  0�8�N��l�	�ܫ�Q-)ӋG�     ��!�����
�L�g��\V��ۦ�hBѢK�
9-;����&�    `b�;cZQ6z\�������y�� �I��/?�$��a�������̂�zǬzc����     `��X�OY&d�	9/��ͬ��c���J�=3�k&k�6�{�$�zT�Y���욑sl    0Ѹl	�^1*�u����Z0~�/�  d����ҥK�~����侴,���MGG3;u4     �-1s3�)6�
���v�f֋D3�\CV�ј�'��/��f�)w�%     �>F,}epT��������X, �  &=�áeK������踷�*�S�#z�ͧ�(��     0U���g,�6K���\���h���������i)r��j�]3�O�     �3�8�*ot��j�E�Z	h ����r�e���/(
�{{�=���G��C^�<     �T�����n#�>x�vSo���a�?'+����ob�%q��T�iv�������     H�i���������j��Ų۳r)   k��AF'�֯W$��%�����-     0����z�_b�Y�BNkmMX��ͦv<e6������#㿑��8�r!�9l��F�?�     �����V��&�����\����RK  ��(???5���_T"1��R�&X�cv��      S��u;��尙V�e����	>^a�ԙZs`d�3��,���K���BN��8�̮�74&     �ی�+�F崍/�e��Ra.����  `j+**�ܹs��k���+JG��P�F"�6�     �є���cZ=��H�i6K�4�k�d�!uV���K�������L�O$4���3     ��Z!�{c���b��B\~�_   ����448�={��{[�-����z�ͣ��    0���L��^w�u��U��BN�l+̮�?�G�GM�Y�uLrZ�ߛgf���1��㟊     dN�;�y�����بʊ
  �̚5K���:r�踷��j	����%     0ut����Ҽ�BN�Mz�Yr�9!'�sͮy�oD����{W�����V�:D�zB��Խ�o(�:Mm	��;,     ���քN	�ʪ�=�^YY���z  ���?�^X�^���x�}Į�M     `jHG��fM�.�9���nv͎�)p7�nI��"�i5K�ߍֻ�k�z퐐s���f����     �gAQH���������ܹse����<  ��a�۵x�"=�쳊D"���x�pEpL?=���    05t���v�˵T�Y��R�kf�)uV��=C��mV�������9'�k��5���    �\U⎩�?����Z�p�lV�   �y<͛7O�����%��ΘZ�!m�u	     L~����Z�9��{VQY��Ys`$������;QY���ВASk�;/��TU����{:�     r�ՒЊ�QY4��U��٩�   �˂ee���վ}�ƽ�ܢ����	     Ln{�����V��&�����M勴�XCW�Mn&���n���8a�~�"!�|��_�u�����=2      �{��U���̚�UUU	   �nVS����ԛ�a�H+����6��     L^G�GRݷ���jx��h��$WrJi��<�kN������l����'��x�sW��3��?�q�M�::�����i3     ��	8c��k����nn   ��j�j�z�g��o��wLM����9     &�D�ͦ�sk��S\��_�sNU����{�f�!u����'K(��a�ԇ�d-�#rYr��B�()�\bv͝�{O�o�s     �~K�B�����n���ϛ�Z  `�<nw�a�M��6�m���Ю���     ��v���p�(�rʧ�y���4�cv]��ɴ�ܣ����:sO���C"��S����Cl�.    ��R�Q��6������   �_UU��vv���}\�9�	-(������     9d�]r��5gV��o���i_��BN�{=�X-Sk��� 2-kw���ݦ�[j�[Z��ӂ����|?|������5%�?�%y�     ��a�$��$4�m~��O   N\������Q(4��d���w�;dެ�      �l�o~Sa�æ
��3��˄��P^x��5��V��'o6MV��R��8-������O
YWQ���f�4N�m{     r��@X>{��?�f�j������E  `�r:���Ң�_ye\��Ɩ���gm޷�     &�ޡ�u��8�Ժ�kD�='����S�
ͮ�y��G���7�9�p4.��jj��҂���{ֵ�[gov�-2����     ��#�f��:�655���
   �	��������qmW�iz^D{��     ��K���p�Q^���o<|��\���U%�����X�7�(�p7���vjic�Ժ��*[�����+/�)d�}���/+1}>�Y:Y     ���hL�q�/���Wmm�   `���fuvu)_����!�v(���;     �ы;�h�I���4��E�O'W����5am�^��u��C��ޯl�j����GL�;lV���O��.dMS��o�Qw�.�     �BgLu��O͙3G��    ��r���Q۶m�vƬ<3"��Ow     &��{�*��aGעc��>x��_y��7����U��;��f�5R�	eC���l;���3Of��\�Pv�w?:�+W_xPȸ��{�YՁ"��v��C}     �aAQH㹬SSS���/   �O]m�>�����S�[֮��tq    `�����#Z�Taj�B��Z]�wOru��sj��IG�g_oW�d=�~�oD��z�<��,��e�����&W�2�����t����CY{     ��bWL��b���N�C3  ��k�=[�=��㸯����hk/]�    ��~����wâ���Z�~ ���CBF}��Gn��̮;�j��)p7�fK��w���w������7��KȘ[�}�Җ��`:j���&     �����=��TӬYr:	K  dBaa����t�m|�VZ�T�P�.�     L6Ͼ~X�h\N��Ժ%����Zr�2!��Ԕܘ���ooO+ْw�+�U�'����
�NkMy���w	�\U�5������{���P�     @���c��F���}>_*`  �̙9s���+Ǭ;ք�
�z��%     0�]�_�Ѯ�Z̿g�xF��Z����ׯ�2���������t���k�mH��΁Qmx�C'�,7��ɳ+�k��ѕ�W^���v��2����od�/��8f�     i4'��7Ϛ�t<  �?��ri���ڵk׸���k[�S���     �l�xi_ZGI�����*!�Z�~ oYc����=8��ugSN�?ٰ/-w�æ�?H�N����<P����5�c�~��    ��+p�U�;���EEE*++   2�~�t<xP�б?�htq�Q��~�     ���Ү�:�7���kz핳*��������/���VŁ��*޴\�1�0r�ٔ3wcʃ��Q�xL�=�����o?��[/_}��6��Oण����     d_�?�c��itmojj   ��n����A۶m�v́�v8gv]     &�x"�'^ާ�5����Ms���_r�TH�۾���+�+�LG�����>e[�܍��c���#g�������[������k{�Oܬ�Y~Z��?�����     ���U�9��7:��~   {j�MӾ}�422r����qMK���?���F      �߰W�9�IN���ڳk�J�����r��� �ESM��v�w��^oWG�_CJ��	�~�����&y�濬��1�6�lr�Y0U��~Z����H:~�v�զ��     �7�0,���?FC�   �]V�UӧO�֭[ǵݜ@X���v�:     �z�B����$ga��TU��yf�vWie!��tD�!�lc����}��w��x�À�H��L0>��AY"!$��rZI�����U�uuO�TW�U�V������SM����ݳ�����y���ޏ7���)�������憛��+�i(��?���F���7��,Z��
��%����}xӅ�1>_z�ة����>��?z��@ƺ1�W���;�����Uk�a!�B!�B�:V���>�����!����B!��<�6n�޽{�J����17p,ٜ�#B!�B!��V6�u�m��4���]��r���o�s�c{��r�!|��o���]�ڬ���$�?�V���V����ۆp(@X ^}֖�&����x�[R7���?{�i�w7������!�B!�BV�-�YDTS��;v�B!�����[��SOz܎�,�B!�BHr��<~��!\�{cS��Xo�ቅ�����G�����O�Z$�<��_~�$Z����N�����+.<�)�k��v��������WN���Ǯ��+/?c�����'���9!�B!�B�ǎތ���}}��!�Bi6oތ��?�LF��nKW���"�7�͍B!�B!+�W�.ݵ�)-����O~�����ǿ��={Lu�������4�5�80�{�=�V���_��Sxݹ[mҧ6u�/<e��w����y��}I���S/9cӏ:�����/���!�B!�BV������!}����A!�BZMӰu�<��ҏQۺ�xj�i�)!�B!�BV�bN�^qFsZ�E�k������w�/����Ajb��[�:s����OZ�K�=�V�%�s)�t�^���On�k��y`d!�}l���={yw��#�ݲ�=4� ���8���B!�BH+pro6�U��靝�!�Bi=�����a��c;{2xj:��ŝB!�Bi7����q����My~����gm�6��7���\yH ���?���]�/h�k<��8z~�DK�-�v�Sx�ٛ1�k�k��st{&wۯ�×�H���n�8sS��-#��|�ʯ�>B!�B!��<�b⤞���Vh�B!��&�Hc��8|Dއ��8�l�ݗ	!�B!��r�\���~�wi�J���a���m��r����o�D����͟�|�Ʒ4�5���A�Ѳ�d&W����7���׹��u���~�����=�'V���뻞>}��P3_G��i��~B!�B!��;s��r�횪b� �B!�˖-[�-N��2�N!�B!��)_���x�Y�1��Rꡞ���]n�?�p����'@<�䗾��ל������;�}���x��,Z���[���~���m8}�@S_�glz�5߼������u�:H��M#/����i����Z߹{/�o�?,�B!�B�Zek�|{����A!�BZ���~���bffF�1�:��W�Z�!�B!��^,���¿?�?�yM}��C]�W���a�s�zͧ?��A�|��?��Ugn~��67�>��ƿ��I�"-p7L���|�W"R��Z/ߵ�������_w�K���I����u��~�I#m��n�k�N�+?�s!�B!��V!��X�)��e�fB!���gs����G�>?��X��P���EB!�B!���m��+�܄�w�6�u��;�o8�O#�~����o�7�
��_t�8s㛚��nq��l"�V�����s��O�_qZ�_��#'E��w����Co?��y�����-?]��Y�����=�d&B!�B!��VS����t������韏'�B!`���x�q�!�����B!�B!��?|�!|��F,�5�u�:����;�ڵ������s س�T���ދN]w�r��=���9�VeU(P_��i\|�zl�m�k��28��>�^���~��o��0����>|��G�[��ȏx�={�B!�Bi�t�}Æ �B!��P(���Q>rD�1~�B7�� F!�B!�����T���(>��g5��:�!�?^��:���W�?��+��Q�?��f���M'���;O۴nx9^o.�-R�2�"������õ�{"��g�7�D�����C_��������Xc�sϗc�2v��wm�l9nq`qxr���# �B!�BH�QM�������@!�BV�������9�_�B!�B!����y��Ņ��k�k�4�={��<6��C�|�=��k��_{ӻ.ݵ��=�e�t���a|&�VfU�-���u�X�
9sY^/֔ן�������k{n�e���7��ϯ��������z��5u��'�uiyÜB!�B!�gCG��g߇����@!�BV�5\4E:��~��.�wB!�B!��1M�o�� ����@��x?�����w<���������:���1վ�?��36�)�6����-���9�Vg��-�w�^��u��޸l�y�6u���M��ػ���Ц�����g�l��y;���#Z��JZ\x��$!��V��YLwT��vɏ;�*4�D<\�p�,zw�)D��;#�J~��B�z~/��Rƨ�H���J���
���T~�0̧��q"k"�3A!��6t���_B!���P�p�}��I?fCg��DE�B!�Bi_f|������D��^�z�7^����n}��ǒ��7x�a�)����{ֶ_]����|��������Up�>�Ė�l]��q��u�����������ؾ�o�����m�_\��w�����z;����O�|���@!�ԋL�pzwDAGȺ#���j ��)4E�f�����0��>��f����T�@)\���+ӥ��Y瓕W�R}�4����gߕ��fB����
�k��f,>G8����P!��B�Aՠ����o��5dMYCA*��uV@>mb6�ͤudx3B!��P�W5�;�.TU���(!�B��c��u��Q��@L�DJ!�BH;�)
zb
b!a� +� �Z�f� +�X��eW��g@-�^�뭔����gК3ET-q�j�P��3U~�0����P�-�l~�[�2Yʳ���n(Hdd�ߚU�5�2���x"!���<��8�t�c�ϯٽl���߃/>m�٧oJ���9����=��6��|wө��/8uݙ���]�H�s��7�Ar��VU�����Z?��s9:c�{���[Gw�������ѭ����g���Ǳ����ι;7u�#�,������} �B����J_\�`\A_�j&:4QE�j�Fz�L
�\�T� �(�%�_����f�5���tyV
����Z��i,/����� �(Ў����k-KJq�t�W��mk��\����f��������3��o.>W؄2��H!,�E�0�H!�15$ti]�t
�H���A7����B!��P�@D�3�
�:��B!�����G4E:��~̆��Bi)�2��}q�!a�k��������/�Ӻer.�_z.�l��2��`)���7"Y|��Oh)f����A0]��y+5z�&
6�U�ee�#f�T�0�P�P�e9���"gj�ME&��TNE"�gML%ML&�	B�Z盿|�n�%�/�|��b������F�֏^���|⪷܈U�;�|9v���/:u�]}�Qˌu������9�V��h��?q�}��;^V���r����37�fvg��o���}'����\�V{��݋���?���3#��g����~�TF�V�B�M11��o
�"@WHGT�A320s��z:��aŐz��������Ei�ƪ�����=��1.�܎�Uӂ9ט�C��ޝ�v�q�}�q���o����X~�o��m�jB�U�E�D�����2f9�'�7���A!��V6tȷ7����B!��^���q��A��;�<2!�BH3��������S�1�X1EG9(��z�t�t
��%_1��Z*���j���*K�*�n����|y(�k�p�$
��sn�Y�y=��L*Yy�Y슏���ͣ-?p�,d��,ܽ1��B�
�`���-op.�ê7���7H!��v��o݇��/-ݗ�S7��o���;&a��y�[���=�������go~�X_Gd�����1����&Ve����g����>x�9+��=���/K�s{�~��w:>��O��O�����7�~���:���!u�? R&������&�A!�=�*��c5���3�bj!33���I"�J��SjQ\RX�P��uk�D��t���qI(�;�����\y�q\>�8���w� �`��8�;+� �^5���t2��2�(?�
Z��b��n�X�_�B�!��0�u�I�Ь��d��E�Bi;�u�ܭ��	!�BV5���cVa����r~!�BV7a�q��x'���3d��a�*�JCϦ�XX(��+P�-Y��;7g�
1���
���Y����qŜ`M�B,ۚ�o�Q�U�o���\�l�2o�5:�uX�`���c&"=D���ݢu-V§�׌�i��M�ӑ�=H!�+�i_���1�ױ"��b���]����O�����˛�-̇>s������9g���c+z���b����j��}��o���:�!�]/Νf<��柏�=2�oG&�?�>�Sh>z��F;��r�H�[G{zW����о������B�������jAp�	�Ur����$���ֺ�Y����%��P��s��֪�ν[���<��׸�h�b�c��`�m�)\��c�\�����¼�h%r7���������x��Z%�kC�D�+�H�j8��ł��������!!��DTQ����tw#��B!��^���
͜�e�����p'�B����`c���.�/b n��s:�T*U8OɪPf�����~"�c�2,�W(
��=��.�
�ʔb��nEYw}v-�r�ߝk�ݢ���ߙ�q(��!���=@4G$ڑ�MFN� i�0��pl������ҢL̥��ޅ�/��;^��������_v�=�ؾ�><�����+�`����8{պ�����ypg̺ Za�Y,_��ꀻ�o{�
������a5���uh8��>���S~�����N���o?��������M'G��{7�t��i�ևC+��2F�b�o�}?�z�0!���a'��� �CYD���M!��G:���Q��T�V�-�^��6g��j^6��f�lmw	���cѱ�\ðO�)��X4v���Ea��̱m�j�c�$06���`��^2�!��5_��p,�bߌ��\��B!�1�!{���vB!��Տ�i�����c�c9�_�V#!�B���l��R1ҥ` j�S�6��&��X���Ղ�f�E~�t)�WI�_��/��c�oh�w���Ex�����7t�Wy�h�o(����YR������[�i`g��X<�XgW�>m�0�a"�60�a��BV�����_��杗r�+�XGx������_v�3{�L�<=�������>޹�˱m���h_��N�v�?x�Pkv�������_��W#m�:]��� 	��قV�+V^�s�t�ħ�9�������{hb6}�����?~�l#_��|w�P\������8�}ڦ������]Xװ�t����o�BH�a�O[��Fv}V��������\!Įd�TzYPR-����z��]78�kp;v���u��v�)H��-��Ƞ�3��5�p�{߅��c�@�mξ�ލEa�~O%aZ�������X�@�3R��p'�`<�bߴ���	!��F0�I�k�!�B��gp` X�=N�BY+��	as03G��B&�D*�(�s���R칠�X~�!<J��ʰ||� �X���ߚ,n��hͯKt����c	��*�B�w(�&�f�����Jw��7�#뀡ő4#8��p`���9^�B�r��I|�_�§�y	"��������s]oo~{G��������g_�I�6����'�z�Í|���!r�X�-����_��y�����x$�Z�],���V���"�n]���w(�[%�^�jO_��sy��r�4�����dO̦����s��Sɔ�h��)9�X�B���O�緎X����n�Vԑp8<�ARUm[wG�̮h����躑�x�@W�e>�!�
�]�����{_ !���%���>��N]�,¹$��y$�I@W��C��E��b/m�av�M���ã��)<�hw����cѱ�\-�Xx�Sn�E+T�S�9�@�h���O�����^��Җ�Zߍ9(��P~m0d :/�����S���a6�:?�J!��#�a%5����B!���	��E��5���-��B!�Fƺ5l�Q07Сd��)��g�Ng�.�@BAjџ�t�*/Q�3���R,�P:�� ��k��\?�ЎlIV-�a��X�w�0;$�C7�P7��w�M��k�s�C��;�F:�DS�̘84k@7�BH����?��_���Hk�W�{���vr~hmW���s��ɹ�љD�d:�H:�}.��'̜q"m�Љ��#_��ԟ~��C�Hh$�P6�5e �����l���uD�\p+c�ۭ��DZ�Ъi����ՠ���<��To�hZ+8���o��Ck;Wt��?�(�����}�A���} ���tGU�P1�Y��L�3�@ƀ�U�Q�-
��.8��.��k��#��l�{����kα̱�|��;��	�;�A�,�h�J P��9�81?��OCˏG��CQ�����H��X��ϰɁB��/o�r�V�ݺ~$�B!�����B!�rr�C1Gmc7B!k��'�����) �@ra.�CM�P�
�6O�d�W��~�X���h!�'z���A���q;����z����Z�� �wi߰�M���Kw�N&a&߰'|�1*�:eFp<�s�:����͖BZ�����t������Z�����ߺO�����o����oi�̮����}���-�Jq���>��G������
��d�:>y�����@!����Ul�+�ٻ��������T��U��H$�`��PNAJp\d�m^����~c�9���8�X�6'��WCCа{#��}-c/+ж(J	��ǆ# �����'���0�]0�]��E�xa�-�B�n�$3� �B!큥m���c||\�1��B!-��ʾ�?�>�!�̒����L��;;[����
��ʰD��L9V#|D��לh�7�5�9�?4%<*/��y�h���Q~�W��7\�����x0?71�Y*ǚ΅px����\�ޝ�B����)�ٗ�ħ��b�wEAV���<��}ý��n;Ж�ӗ~�O.�_qB*/<V��d��ƣ�&@!��Xa�S�4�F���H-X�LAM��0{rQD*��W�݂�vAJ2Ю
�-dB�ݽ�d���E�ns�&h��~,+X5#�$��6_��yA��jl?�1�N��\�C4�=��2B��z�'�<;i��\{\�B!�����p'�Bi+�0	�Ũ�B!�D)�>�!j$���A:��:��P�av���(��vg����Z�e���ߜ�Xt�7�܂��n/�z�A|C�p��7���B��r,s�%�p�j{�f9!����Ӹ�ڟ�Sx���?��E����n���V[�-nyp&�R���}):ca�����<>�ջp(�'�R�bb[�қ���Zfr�Ш��)�.����X,^`�
���U�vQ�]-Vy�#N�"P5"��*J'lk�Y��'@�0�;S�V5o�1������d�)�\=�w{K{�p��O����3�����x��R���d�7��򶅄Bڗ��\Hɺ����!�Bi��@�G��B!+�h���*�#���X�����0��.5��b1�B,�2,������9�2�N�	����փ���k���m��G��7t�c�ܯ����P'���xvR����	!�ɱ����_`��_��NY>�<��?~߾�9�mp����cxߵ?���~!��!�¯�>�O�x�YB	��U!f�c~z�n@�ѐ��P� �_��)H�lo�8�'P5F�*|��[Zp��ƕ_���Ae�����).��5gؽ�xI���ī� !�ZĪz+_�E�r������}���`L`(?���DGg�xf���Qx�BB!m�l�������B!��=��]�/TU"��i&R:uB!���U��!��@R0Rs����:�!����߿C�����w�=��z<D���eB(uY[Zw�����*��[a��cY~��Z-��Ҿ�`���aw�oXC)Vi���͟?����9!��r��ځC!<9�C*BY�X����+w�^��w�� �g6��_�p��ڑ��[<1��_{;>��sq�� ������;��o}�pH!D��!l�3Ы$���F*��VhUА(QjQh��{�=�)��%VY4C�*�����$���Ħ��űR��l�9kns���a#L<�Z�2�sf����̥y����岗�jia�Z���֜B�0�.���[6���:��ޠ�ԡ���XP:�oN�S�Y��BY�����ވ\Qoo/!�BH{��*:::��� ������ɶ�	!��eeK�{��P
Jf��@F�2�")�ó�OT�%Q�%p���7t�#Z��+|��;ז\��R�X��+�2�:#�U%Y���X���p,(�rY��+t���~���"��^�U�oX*�͏Ǻ���>��.Le#xvJ��&�	!k�0q��?��L�CW��X�EI�������_��T�ʚP�����7��=goƟ����C�`��$����o^!�o6�j8u�D��Bva�D
ꔊ�b(=��"�@��0����#<5��=P��x��/�
�b]fw�P��zU�]�IKU�AEH]�KM���y�LM���e�tQ��ۃ�n�w�9���iz�a��5�\3Zj�K�T�}�|�X�:�o��)���F]��v��}Hk�8��c9d�cBYt�h�ܹ=�� �B!�GoOO��{�wB!�^,q�@�}UKC/x��;</�w�H��;��C�����_�ݹf?.�����[���K�*�����EEY�	;uW�;b�",ۼ�,{�+� �;�P�+�j�w(��b���+�y�s��ǻ��B�{?���U��x�4!d-��Gb�|�m�c��>��a�e~��{�ٜ\i�jeM�M�>�O�������o���B�DSLl�^�J��	d3Yh�V�]+�H�XLf����#N���P\p��u�r�(�s�y�u��5{�])����|�u׹��ŧ�Ƭ�">G�n.-���Ax����ι��{�~I��U	Y�q=A�~P���ǂ�{�897�?��P~���^�H���1ު�BHk�ѥ����!�Bi?���G�H��5A!�y4E����!�g'��d�N��@���9�٥�C�^���z��^/����v���/>��_��/�U�<��}-e��|F�c��8�.�z�a�k���B���/��E>a�k��l�o'G��CR���!<5�C�y��Ҏ���U����T��?�Z�>!�15��gnz �<sk�5p���м������N��_~
�!�Z2R��B����� �����0N���e�ca���mZ��*p)��l���R2A�z�,*�C�Ő�G�� P�C�g-�����B����&?9.�����#�k�9��!�5�6�7����5W��e�|�
�/>�,b-�ŮF�1x�=� !��c���N�Ø�-�/�����
�`�\O�@gk!���/"��`]?1�N!�Ҟt����!IB!d-b�b�:��]f��	d
�Xb���=B�A|��5�[�z�c�B,�",_ѧ0��R,�1��Eٵ�ؽ=��Zʱ����{e��7�n�	]�l~a��z<CO�P�7��m������I��Bx츎���;!�����'�������`�0�\�{��õ�<����)�^sw��n��?4�x��􊳱k� �k�
!��1ءb׈��P
����$0a5��д�a�*��)L9ũ �� A��*{ �z�,49��kp�+��z�}���5�q�׼��������qNuнJԪ8�<_|w��ͪ���U%j���P�[��|������k�42ip�
�/�Ǝ��H�rΥ������ul��XON���D�B�J�%p�F��k�0!�BH����l����	!��Z�ܫ���bC{bz��eR��/��������n�bE^��G���>�Ǹ�3��W{��u�|C[Hݻ��x�9���P�	z�y{�e߯xP9��/N��Aw���
��л�Oq��������+4%���ݠ�0�xu�Wh5�?~���&�����{>�3���O��]v
B* e9<�����C�	�5�d��ľ�������ڀ���K0���γ��q�S�ˆB�*��;���6ųP3Ә���:c�]`�U`w�KRA��T^�v�|Yh�X�Mh���"��x��J��s��c����W�U� 8^���V�9���A�KbW�\Y|*	Q�/�9��*�+��� �h+=�Q�hd4��%\U�6�D�������9��\�50��QL!dy�
ɽ�ttPC!�BiW"�4U�n�]FT��e�ӄB�.*v�J�&�L$�Ni�R,U����=DE�����
������%�rNX�e�+��j�����Bqٕ3�.w\9W9_�&>�6�����
�� Ǖk���⋉}B�\E���:K��J��B�~�w����X˰ܼ���Fb���x��^!!�m�du|��O�����j.۽ĝt���o�|߸�idrk�}`M�-�����g��헝��\�Ѱ�ĉ�$�������_��"�����C!�ܫ#n�bnjX�_D$�"R�%�^�ك�"��C���dE*�P;��$C�KBՒ�T����}�k�^t���׸�c���s�GD+� �����|I4�r�
��E�ҾB���_�D����{U��?�^�`U�pe�D"�s���\٩���u\5�52�\�/΅�رt��1!������w'�B!m���utvbnnN�1�!��5B!k��
�2�����R,)U[,Ŋ�U��l����7��s+����v��l>�T!�(��]�%���z��Kߓ�� �Nm�X����q����U����p���R,Q��'t��Ω�����%zy���d%���Ӱ�B]#�0"}8��c9dX�NY�<1����{�ғ��������%����<| _��1��Ma-���%��w�/��8n�ճ��ғ���@���ff!��|7��ܚ�!dmb������vf��sЭ[jZ��H*��f�%�^�HU!N���Łw��Q�&
�/���Seؽx�x��<�s�sn�n������Տ3�.��jw�,q��z�+ /ދD��^�w���w�<6cQd�	��d��^�Uզ�Us��<��Y���6��Ąى��I�BH#�1M.�g��B!�����$�n}Pr*B!���ҧ��!]�,�'af�&5V)V4Z� 5M�˯K&�^O9V��Q���5T̋����?(�Ek��Z����)�p1VsB�2�X~Y�X�`՜�V�%��
�aw/�P�����	��2t��GCW� �n<vB����	!��{�9���=�Kw�ǻ^����������y����'�ܑiܫ�Idp��?��޽o�d'^w�VtD�֏i|6���z߿�y�2LB��*�U0�. 1}zRG:�n�+lX��$��JcUN�r���<Ghw�{�ճ��778ϩ^�>��w#��n؛j=�9_ٞP��fV�S9�
�{�Tr�����K��xe��o����F����RM�.BVb�"�1\1�5<�t�ON���D�BH�X��^����	!�Bښx<���0��!��V����rK���40�!���B�$�B%��������p{ �j�sNT�%������j����2�~��>�������潎k�y��by����/(S���\
��۳��X�oX�u��)(�N7u���j� �'��͑��4'��"����!���a���M�򒓱m�5�����;�?�o��4��Ybm%�`��?��G�՟=��>�x�v��V֧>n��s��#�3��u��Z�1���~��榧�N�A����T�]��D��F5�WRj��f�|D)���6.��T�0�S����v��Z��=W�f��������߽,��.f�"R�߽�~�l�]J�4��5��]���C�K��QY��t�B��˿ot��[#!�BY��@c'�Bڄ���������G&�.����q�7��^�P����;��}=CQ�]^�	�׶�����m.��r��)��+}��W�5�`�h�~�����=C�B,�&.�*yx��XA��A�n���;�e�0&��_;�;ABV'V��և�㶇���x��;q�����n�YHeq˃���ñ�H5��0��M��_>��|g�4\�_|�z������H��'�rxp�qBH;V��ׅ�)�@f�2�4�I)u񶁚V)Jل(-�H4�.'J	��a�B����E*g(�)L��J㒈�?W�&�w�����YrN��݃��e�dB��q���h�t��D,	���Ʌ�����+��%
��r�����>}#8�w��:2�B�&����b �B!�K<��^\��@!d���Wîa]��&��(H�E/0s	��q��F�ܫ�C�2,A����h��ʗ`y���(ƪ���y���y!�8Y_0����݂���{�Y��d��
C��z��B7�0�_�V��8g�	:j�NЄ�Չ�W�}�+l��37��݊���)^z��4~p����#���@�a�]�B�
�[�`w��ސ�6b���U�)�l���p?� �~�(��BښH����6w���9��BɤVhi�B9%Jl��Tv����Cx�;o��T�t��m��I�W�L�c�9�9��ZƵ�:��F!#f��ڝǵ�+*��{�л��%��HUja���D,�<o�ۛnw[��Z�EA���5=��(.� �7c�����̦i:B�&�ʷnZ%�B!�K$��^�wB!�E1�k$���Y��H&�	IMC$���P����B�OP�K�K���b=�X�>�!��(f_�p{=~bа{#B�~�bP�Pf/xt�op���b�*��:6�������wQ	�K�]�͕��=|Ɔ.��A<3��v'��>�&��/?{_��)��s��׵ʩ;��/��|�?z��ٵ�D������Kᦻ����8.>m=���:k�0b���B�?{�<s�<}i��	!�K,��v���EHN���#�ZlY��
�va����.ѼPk���ցN1�~�ڃꮡv�M��&H��굼�n�ZE�Z�%�n�OȒ�d����㠂�нz�v��W����ұ|нV���X�]E+]tl'f&5�񲘁��$"���0��[�B)�T�B�Њ]B!���!�:?�R_ ���h��3�4l�B�'
��t���bq�",��k�ӳ�]���-����b-��⠻��Y�b��
��6*��H�,H�=h�=�_�<�u,�����B����y�~�X�A���v/o�*�������tF�6��v�Ơ���(9�� ��!d��������G[�{*��1�����v�a��������80�{�)~���	�u2>��w����C*vo�[��{� N�4�xde~�V���}xt�	<��	<wd�p!E!�J<��uj!Ԟ�<c�(�,X�O8�nZp��۽B��!w[��j��&Q�]u����X�Z�*[��B�[��*H��Ya�Z��+���c	 �N�=侜��hι&'\Ʌ��,�ycQ��WF�q���.b�,GkC��z	ZU��v�%�^�怹��ѵ�v蘂�s:!��]��ܕ��	!�Bڟp8��(�	!�� �b⌱0�u���G*�F:]y�g��������9���"��j��ay{�~>��S���m܌@����M�e��A�B�|3��Z��Aw�?(�����r,g��t_Zw����g��j��
�-;q#��7��ƑL�=�C��]%��0ٜ���:R�,6uᬓ��{s1��R�w+���)<���x?�%���b��y����f�����y��F{�}]_a�~�c}�0|#H���Z��sx��la�>�qxr���tET�t��e�'�YB�Z(�HIp���{�۽�)�US��.Fم(�XdW=Z��T��TK�]r��]�w,s\�+.���J�p{�d���������A�P|���f�Es�8�^)f�D,�he~{#�Sв�9T�5�R�{���oC�Gнj\�l�&���g�:.�2��P?8�`|�awBYk�49�"0�D!�BV���Ȇ�bZQoqQ�!��e�j��G&�F**x�V���;��A��@ޡ_)� ��ӳ�����z��Av� {-�ߜ�8�Zй���IhY�����?��fz�A�B��{�r,Q�������s�a--�n�a���ŽU"�m�x�`�R�������BZ�'�����P8�a�X/N�oV^���Zy���Ɣ7Y��'f�8<1��[��<���N#��'��M���\
��쑃�y�w�;���8z:��?<t���G���R���h�,�Kf
�LV�\*�م4fL��Ǧ�1!��%,Q���al�/6�O����HYd*�QU��8e��ك
U"TU��.<�ϭ��	O� ��ze��W��"�>�Z-c�qa�� �=�V��pCZ��E�r�G.��+X���_<�tY3������U�w��X�����97{˻g�]$^��*E���g�]6��K.�Cї���B���P��4��B�Z@�u3�wB!������"�������U��BȊ`��箏`sləcГ:ҙP�g����ޡ�Xk!V�R,a��Q����^[1��g�,�o�����m��V<^T��b�]���kz.�x_�����;�ޘr,�gh���6��ݱVtX���:�n=�������8>�?הӏ	!d%��K���=V1��0�ׁ��z:"�툢+F<Z�PwD��Lgr��F��`>��L"S���&��Mb|&Y�������o}���!�����A~ƘVhZ��Cv!�d�x�@�d��L�P�W��k*TI��]D)�0�� UZ�Zs�������mέm�w^�V���F@��{��%p��=�ͪ)����Jv/���W�w7��&b�ir�γ�W�M����SsЌi\���ً����Bڙ����6OB!���X�}�w��ƀ;!���eǠ�����Ez>�D���b�@�X��w([���.��]K��a��yR>����oݯK����	�{�؋�U��^�Ң���z�9�{�������������
»y����B/O�o�o�+�9�?ق,�]�EEY%�*�����@�9���+���zh���(��so�"�;��x�h6��-�aB� ����㳅���HBiY,Q��~��1$���
���
U�*�2�^��`�\�\�,����
�����(���9�X��{��[���B,r���y	\vAH0/z.�����լ����K��W!`���M�}�F�@[����0;��^ӧ"�?Z�-�d�S�"���BU�4U����B!kK��VP�x�H!��la�@Zb���'��v�?��;t�E�`M�v��t��+Ū�+x�=Hx���{��8)7�5�&��s~�2jG������J����)Ò���A<C�sd�����s��dU������b�*�0X�]f=P9�c��8�����c1(��xx"��r �B��BZ�����I����r�!�(%���{	UKk�bT�%�;ŨF��D)�F	R5ڋ�c��TS��-��p_\��d�[!�����ye)�M�����B���p��"��9�V�W4�L�*	J� ���aq���
�;[ݭ�u[®\o�C���<=N�B�U��G	t"�B!���w�LB!AY׭�Q��)�MO�C�T�%��[���!�B�Qx�+����<���X��s����K'+������^>���c|���as�kz>��'�?��ceʰ�ޠ�M�kI��^k�
���2����X
�W��;A��>�X΂�z��@~��>��?f� N6r8k}7�C�暴c�:!��F;!��'�7�pc��,f'�C�P�)����@�� Uoc�S�*�-1Gu�+�[
���T�[�����%H��~Ⓦ UK���@�St	N"��)z�͋ϭ�V�v�"����y�g{�Z"1Kz�[~�w���~���
Y�Zjog��+���K{�hUo�]Z�ͅ���HO�V=��ū���H�^��Z�$/�4�	!�B�A��4u�il�BZ�Ψ��֫�3�0;=LhHi��x�=J��Qޡ�oh��˱ľa3J�*���{��Z�Uw�����e�+��LY��9N��k������f�Esr�aP�Х$�����c-�_((�ҍ0��4��~�����6�	���&�Y���B�wB!+Ʈ�N�M#3}���(�
)QȽѡ�ʦ�@{EÂH�rIբT��
V�-j�)D��Pu��+�6��$�rZE��KdQʿ6��$��� K�xQ0�3��<�	�;���,���}��Jf,�� ތ��E�kȽ ^�x��~�m��wWUs�������!3{q��rԮ!dU!۸�ɓB!��N7�C�z�B���O�I!9yƔ��J��Y�;���EX���7���C�2ޡA�E�Y2k��A��~��<���9)���C�-ê�c���0뼴�`�e�J�dʰDs�����ߧϾ��XA���EX�aw�b,{�=h���gX����Uw���FD��+zT��G�b��濏���BY)p'�����T�t=Н=���Y�&�����ea�qJV�Z�J"�(��#R	D���vQ3�E�P{�w�qq��x�%@9%/�IF|�<%���3���&�M�*=����K�x�s+E��H#�;C�N��X(f	ּ�+���w���л�^!8�����"�3�^KSC�s�x^bv
�	�a8�{O���d�BZM2��0�N!��&zݧ1�N!�Fƺ5�7�#�p�DɩP�ۋD"�eXn>b�@����+PS{�R�꠻ES����.ǁ
��u?�P6�n���3��F��~�[_�=XQ���Y����Uޠ���A�t��g��Xr��`A� a��V���-��K��Ɖ����pź.�Cxp\���BHp'��t4����������Q(S*ҋ�v��v{Ƚ$>9(/A�O���D*qۂ]���WTn���U�
ԮP<p�&��Ϛ����4",=L�Y�Z	x��s����b���ʊ^�w����,vy�.������Dw7˹oD��y,v�U���W5��45�v݅c����<�����ԇ�� ~u��B�f7!��*��9��!�BY��0K�$�Bd����ׇ�>\��I9��?�
�{b�|���K���:�����9����W��Ƌǵ�k�m/U:
pn�*dh�W����~�l��z����}+�r����cA�}��cy���=�V�*��t�~�g���+�
��B�@�m��p�)vcB��wB!McK��s����Cv!�D�jZ���+�)�`{��5,D�%1�[���d���E3�����`,j�M"��Kp�
��E!E�Z�����J��Ur�v��T�O��	Ż�S���b��Jl�
���i��6J�jdؽR�2<����%�Z�rXU��R[C#�e��zy!�L@���e�
:6��Ssx�X�BZ���h?���	!�BH����i'�"ÎA/��!7s��,��?\�`���U���;~��/��}��ڽB����縟+��y����}�{z�~�wн��ޡLA��?�r��.7*�^�7�˫�=�.��Z���tw��3��xU��h�������	!��À;!������1y�z���>{�(ғE�)j�-8)Q��!Hɶ���U� ��(U�*Ũ�}��$
���-�p/��s��*��� ���,��x�9���V����7��ڊ��U)B��Ĭ�k�V!�6����pwWT^!�+W
X>�U��/��K�r�V��P(T�&�bC~��B��]������
��2 S�i0�N!��&z�g0�N!ąΨ�K6(�L�ca~��P�۳�څ�v�b�Z�����^�%�!z��[�K2��^j/?s��������~^XU����eY2���<:��,�f`�PQ|��`>aб�_������VwY��t��V~�3��;����#ؤ�p��>L���&�Y�΄B*a��BHC��p�:��1�����h4Z�dC�v�I&�.��C�Ά��H����dw��6��Ū�|\�/ι�P�S�Av?A�/�.+5>�n��~��H���D���J?/w�M,���.�|��c}�����`,�7�s�$�.+X��J⑟��r/W�-�.hk(�[ZdCg��!^Y����.�V��c31<=��B�JbH�]�|E!�B�pיG!��`�@gd��>}*��B4��{�ڝ��A<Ċ5E�������;<;<�z��V���;����<(7_�-��`������]��ׇd'`�<O� ��tԋ=��\鑐��ʌ�����C�>~aɇ�)Ʋ���	�;ׄ�"�Pv/̇�J&�����u�	!�T��;!���Q����&���T����m�@�W�H������r�}�i�l��}��XtA�p{�gԘ�{a_<�
�{�M�(�,'<y�N�b�L������g�������[X�o��d�Y�\�������)rn�V����A�u����/`���e��)`�ޥ�*A����](^-�4l�sص����~�~)jW����������wB!�����o�@�>��BH{	naT����r[{4�*�
z�g��vg���7��ٽ��ܘb,�F�K���t�]�#V���U̕G.�kb�I&�����Z�e<?ْ,�c-ޡ[����U���w�7X���.w��pWUk_�_�����rн��|����
��tq-D��B��	!��/���Lt��#�0�D*�H$�f�im�	�ˉS���8�liث������W��!��av7�?�4�^k�}����$h��� 'A~���k�BU�yq�J�r
W�9W�'�^��p��w668E,���]��hxw�ݗ����{�!w{��+�^��Vwun����_���G�&��N!�v�� �	!�B�F@�L7V��F!��l���,����L�-��J�d�����|C�B,�b,wqJ�dC�>~bc}�ʵ�^��kʲ���V�������0|��skg��;tΕ~�}B,O9V#
���� �a��ݯ˴a��	Z�'|h�_��0B=���x�~!!��Qp'�"ͩ�!��I`~��)Gۂ�0�Ӹ\�r�P��
B�b��0U�(T���B�W��O���{�O�
�7ShZK"V#~��� B� ��P������A���fq�K�r�J{��{i_o�]�� ��\���{i�5��U���л]�
��-���8:^�m�3}��p&�kh�:!�T�K���ks!�B����}��N!kMQp�z�p���G��,���X��/t�e<C��h���m�b�P.�^z���b�b�+����y���%Z,��׎c�ʲd6b0x ^�#,�U��nw����"�z�����z����*��z=C�b,��
�!w���.�"�0=y��^�m��~ܵ?��W!d���;!�O,a��M�kS���@bJC8^�B���v7�JV��;C��R��`Ws�P��],JY42��/��E�T�|�������yy��]�r�H��Ĥ��~%:y����	�~�Z��	Z�߃k�C��}Ѐ�ۚ��%���W��+��.�� -�^��-�[rv
��q\����QܾHf�\BH3�%/	ҙ!�BH��	x�g��:!��֠'���M
"s��^H#��J���J�Dޠl��������ڽ}Cg���ؖ(�jH����{�^�E�<�V�W�Z�[�%�Z~�_�c��;\���	������?εJP�����R�%*�r��aw�B,/�01;�}���߄�ᎃ*�S�	!��a��B��NK�ڠ�3u��$��@�x����R2��^b�(��lmwګ��m�BTu���M���Jc�x<؎j��[p�MA�4Bj�����f|����e����z���{#Rq��x1�n�<��X<�tN-���w���p�lg0�D�JQʴ	V�	W^awQ��K�*�4d-S=�"^ѫ ڿ�>��Y6BH#��;�M��B!m���n��=i�wBiw��p�`ɉ���	]��˔b����fw��v�v��>{o�V���!����j;.IΉ�ۋFy]+�����ѥY+Q�����]|��kP9�^�U�K�K�z��=Cw����S�U�ݟ����^lu�'������t{OdA!�=a��BH�{5�;�Cf� �)YK���7&�nkd(�P�x�J��	����)�@�ŉ�����
Q�"���P�h�h�g5H�NПaPA��f��i��l�T���:�,�Ɔ�~��Z�+籼xe���X�r���~��2�Uy��\���a�D�q�a<���o�0�N!� �˽�gp'�Bi{��`!���@g�"!��-g�aG|s�Ǒ����9�w�G���J��C�2���$ˢV?ѾV�Ń&{�K�ιz����w���֊�؈_g�!�Fd�[�U�O�<��8X9V����q�й.�	�<Cw�P�˫���@{����#ؑߟ�m��~�u �����[Bi'p'�R� Lu�c��Q�'�BS8$L�����.X{�&:��^"�P����nXO��|^qЀ`{�k���r��k>V[��Z�,���(QJ��j�=�%������/�Q,jW��]��ڣZ�
"\��5�	W^��"�J,bم+�`��p
���Sˍc��^L����}:�4�	!�fd7�����!�Bi?��t��u^BH�)�x����1$��Ȅ�D�
�/�`)~�a0�P��"��X�+Z��Z�ܝ�J)V+z}����K��khdAV�ʱd�K&��5WU�UK�=�W(�s[��	��CgA�o9�O1V-���f�������	\����QܾH�0$����wBYÄU��-��Ǳ07W�*n#(�B�����[\�م��]��R�	��V�y�~���fo���V�Z�ZF���<��8%�J����!��_���aq�+f��n���ܗD��vww��?��'^�-2�v_�$X9���|&�@$�<^?A�s=n?,���!�%����=#�!�BH{��]�Ò�BZ��.��0fB�֑����54���>>�"nk�mm��-��S+^�UK�}%K�����F�Y�s=��Fd5�����y��� ���2��2Aw���Wh˄�E>ae�U���Fc���z���G�/�=*��q��0��1�N!��	!d�Q���
"s���J#�����b��@Z\�%��u;A�G������	��	V���@��
�W�_��_���;̾��+!,�F1KD�d��d����{��{Q�Z
��ķ;�ޥE����	�{�ޅ���@�@��VÂ{.�i����>\�	�6o�]G#8:��B�� ��T:̀;!�BH�J���wBY��:��y�OEn�n�~�X2�v��v7�P����u�g�Zi\�+�1�.p�d�K�X��:�٭DA�j,�*=u=��Z��^kK^a����+�����X��a1���8��B&.޾O����BBY�0�N!k����7���x��b�bh�'��lnw�j��o#轷Q��9�^�p��
���'o!j9���
E��(`-_c���ts{���_�h����m
{{��K�j|�=�he�t��e@�+E,?�JZ�r��C�!w�}�4��8��4];�၉�0�!�o���L&���!�BiO��{A`��BV/g�aG|s�Ǒ���D����vY�P����n��o��b,���Zq�R�:���h��Z)Q���Y��ˍ���3�n���+%j��Q�dz���qgq��m�_�5]⿪��E_�=���.}Ӟ�N���b7q;v��E��$J	�  ���3�w�ޙ;��|���w@B0x�����x�}��p�
����u���w�=�KU�e����Aw�kKs�`��3WO���靻� `�@�  � ���S۴�x�����^�B�B�h P�	�+ũB�+0�����ٝ�!bQ���i�Vq�&q�a}|�Z�EL~N�Ǐ��%N�	��BV�<c�Ƕ�͏)����ʦ��Y�]&`���>�J�lo/��uZ�����*��]"^9���=�Ӥg����G����  @E���kx     ���Ɔ��Zw  &
�}�B��P��W���]l�;>a�P7�^�x�A����]��^�{�}G�#����;J�Ϊ�w^ܹi�sTH�$�FA��r��y6˱��^�{��.�����W����0�f1�q�����ame��4����ct��_ߪ��g|� ����;  �0=P�'��h}�.mV��QQ��"�B�
����xT��@�	�A��e(H�P~1�}<H|�܍;6���sl�Թ���-jP^���63�|�:���Z7��=_o�(b��v����c�'`��������V1�t��:�TA�����umu��7�ӣ�;�կft  ?�u����     #M�Z5or-	  `p�
9z�b��n�Qm�J[�"�۷��;�l/��}C��!�S���
ǈd��y�}Pb�9q�%u��?�-l�e�>�
���U�.�

���B��eeX]ϰ3Y�������+@�n��mA��n�KtB��w�Y���:j,�_�;D˥����&�w  @FA�  F�''��pw)An\(��%�L�
�z��^�]ּ o[��l�-��t)1���ڶ�U�*��$�eߛM�I����{�#L�OK�
%��;��K�_	�{�js��U���A���UAw1�n;��R� �J��pU]���%��ţ4G'�׷Z�2��  i­�;�w�<��.��    `��6��7
   �,����D��Y�Zڢ�bg�g�;�B�wh^�lW��lhO��ݽ�=�Οݿ����@�(b��a�?��ų�U��c�r,��s�����>�J�B�����V�(�6���|C�,x�ۛ������S�i����M�$�  s �  #�g&�4��V+�=K	��)�(ſ�jW�=bT�(�p�	Rq�)�jW6�+�)�Ͼ��c��)ہvS�b��I�L� b%�=�	����ΕD+C��x"V?�8�}��]lfh��;�����y��{��agG������}�R���R�f[�����p%��=o��N����si�t�~9��� {��;��9:X
�!�    0�l��Tom&T�L  Y��x��?�CͥjVv}���p7-���ll�)Ʋ���Gt���V��B�l<�HR�Y�?�0de���8�+t��
��,�.���q3�p�������+��,�b,��
dpw�� -�c�_�h�>�T��GDG��+w��$   � w  ����}�<b�N��$Ԯ���BC�+P��RњLE*&H����P{2:���40�{�$�ϙMQJ�|Q�)ռ�Ĭ8�w�u���kOؽ���лJ������PO�r�)7���k	WRъ�gv�!wӀ�+\5D�J"Z:�������h���;  �;��q����:    F���u��6�u$  �����/�ݡ��m/�8!�����o�K��b��G��IR؍|D������!�R��b���h�g���rAV�>a�83������{��.�<Ü���<C��s����,KA��b,~�i�y�Z��b�r,a%�F�&}i��Ν���.��&� `� �  C�l[�ե�l�6.��S|?A��
S}��8N7�.����1�n��bwǑ�C���~���Yl`Ⱥp5��J���lSa��YI��b�L��!��,E[C_�]|����֠�����6=�U���������įEA�E��?�.�����\E�  ��|����~m_[[��G�     -VWW���9��gh  ��`��5Y[-Ri��܃B�E���b��,��<Ġ�{X�]�Cdb�����
��B)
��0�m�{QH�{TAVZ>�jlt����~W��� ��	�߀v�=�3�����,����
�?�.�e�Xn��q1�`C�w(	�oVnї�s4vAw  4� �l��}�~qJ�u�'L��Rg\�$F����ıLX�J�R����C�s/@��7,"О��$��a��&�sE8KR�
�o*h���6�/�Un3�j���A%\Q��՝k(^�	W�vwؽ���=�*�mj���f@�]�����;┧�]����n���g�Sm����5�[ ��und��]]E�    `Y3����  `�����e��v��r`���]/�./���,�����2�I>ԎR,s�8GÔ���8A��d�
���M�B=+AG��ߣ{_�������7�r�������лS�%�|�����/��[zk�6=w�h��Yzu�D�U�  �6� ����ǖh�l[<�T�r�z���=H����D�(B�
Q}�f�=\�JW�t�=�8�:O�3.6�l�Ra�~�)h�mZ�2N��%��vw����$\��X�����n�Q���Ղ�/��C�`o�B�,X5i��w�Vw퀻0�#`����;ݨ�)�q��sAw ��byK?��b|     Á�u��V�   ������M�Z���b��>�����C���a�3Tb�<Ĩ�Xq������XL�3Ho�X{��*kY�V����y�6���vUa�n�>��*t�_P���wz��a1V�k�����B�����fe���G4v���e�����
  �� ���](����2m��e�TX[�l)�>q�n�SrA*<�֬����Ѹ�F�=�@{RB� ��������MB��=o��-A+����qQ�v����b�]G�����L�R���;����~�muϻ���"^�P�����b�]lg(�o���wό�Jy�~y�ul���  �K���U�    F�L���n4giw  H1ؾ�ۋ]_PY��hm��kb��bp�ݼ�]+��ON�}Reyuy����3��Q)��K�X��1��V���0긨^a��Ӽ/�+V�]�o��v}��r,y!V�#l�o*=�N�{��|��fw�Pluw���G�Aw  H�  �|�t�ۿD�K�,��UAv�8%�Kĩ>a*X�R�R�!w�O����v�P�y˂���AV�c�̉3/�s��`C|R��(v�4[L�'x������&��A|,_�]%bQ�x%�u+w[z�U�x��:"UG�r�+���ٗntW��VY�]�׷��\���=@�3���z��L��%  �Z#O[��¯8���    ��`�u�ǟ�M0Y  @<���:m-�h�U�v��vo�]]�^���y�q�CYѕ�Ku_r����c=ԎR,���:���H� K��Q<Bռ$|B��$�����m�m���{��>a�z!Q�_���/K�da�v�V�����\��Y:��x��+A���MY�}�hl�<��N��6�4  $�  �A<^�����Ze�j�Bp�]jkj�������(F���U�������(��R&����Qm`�!%)2���e��B���
S:�+N�d�=��%����M���c�"U.@���u�^SC�/��ks���
��l��v[޻��Fw�pp�w����{k��ڢ��}��Q�n��7��	  F������ǯ���~��     �����x��,���  Is����]ܡ�e��X	����(��x�����աv��vm�Ђ����cj�Z�=�0�^-�&��fEYq�I�c��m�QO%��>~�_(����2�0(�.�Uc��ݒ��*��G��W��5��A���[���9;w�^�U��-� �6� @�8{�H_<�IՅi�-�\.�E)� l
����L�*x�{�)aJ&>	U���P��A��m�M���%Zŝ������_��T�9l�S&��ld�#`������9��+�64�
V���������/`��{��v;�O�r�"t�uĪ�L�R��1��:�/ыW�k��9� ���V�N��[�Tp    !���Ưn�Z��	  @B�
9z�R���ߡz�������a���j�P��n\�m��Hw~Rb���}�=Zw�bٛcs~���"q�(�4
�P�|\���0�.)����ð2,=��-Ē����^QV��]��+�W�n��M��d>�t����4�ߢ�.����m5��k  $�  �����g���봱��ry�`��h]�k\(�ۃB�wF*N�UM�J�e!�����(��I�Yx����!aJ���V\1+�U��(a��e$^���)(����V�:��kto�m���U[��os���*���sE�B��'�VW�\�B�]y���~��8�x  Y��p �*    �Q�?�/6���?   �S���K:�5K[K��[,��ؘ�7T4�������C�2,U1�Vȝ���w�h�a�P{Z�XIy��X��%�/��%�����b� +��Xi��g�J ����J�r�}�]�:�_(�{�BwL_��t��7�CW~�d5+3��cT������z7���  �@�  ȁ��p�uy�,'�K�RIj�5-D	�w��6�{*'
N*�*L����a N�>���G9Ԟ��{�96�y�Q#�sd*��=FR�j���{����zawy�O�2��U�}=�*���e{"�(\y���f�^����.���{a_���ͽ�	�_nT��W���4��$  V���"@���     `��V����e4g~w  �I.�K�_*��wis�F�B;��������?���ڃ��@��j�&�X^?д����s���B�&�kc����>�����hz�
��Z��;6ʸ$ʳ��{�a�4jtw�������c�}�p/��4�;�@����ms�	���X���� ��hP~�}��Z(��Wo�[�/�s  �
�  0 Ɗ9�ƥ֝�[����,N��A��_��)�@���֮/L��R�v����~��a��վ0���,d��.�%J�϶8��c[��9_�U��{?A�U�{1����9Ab�L���z�J�����BC���=ls��\K��.�ݫ���'�9���y�ŝ-m`�v �𱺝��f��¯X�_[[�Ç     n*������  `�g��Ra��˫Tw��E*��mm�{��~���ҳ��$�Τ�"ԞU�tl�96�&y����sg� k��c%���vW��x��{.�K�/������r,�ս�6�^������
�
��}y{k�ƫS������Iz�N�   ���;  ��ۺpls��7��r����S��v�h�i^��Q���aJK�j?���)��� C�iVI��3�����9lD}��nf�)N��7�l�IG��.��D��}� �/L��*��\��73��+��R�).C��-G��M���T��b�,��aϭ�Y��x�9:w�~:���^�  �D�i�p��5z�RA�    `Xl]י�����6�  ��O��EZ[Z��R�il���~�|�R�V��.�2.��'C�*�D";�!�#̚?8��Xix{�_�[�e� k�ʱ�'F)�
:v�y��>���zz����W�v��c�W�V����X|�������F�g�Q����2�x���v�>Z@�  L@�  R��%zd��//S��XN0D�
���z�#H	+X)���X��.FyC�Ο��*���!M���ci�c2�tl��q�%}�ax\�
P~L~V��β8%?�U�񠰻)�����U�h�
��,�x%of�	W�x�w����6����h��F�{|�U�šѠFe���D������O7� �n���߿��^�B     `x����w�f�ɮ|  �g�P��tz��Ӵ�,Ҿ}�����=�=D_V��,Ԯ
�{���X���ۃ
�\F�?�9&�q�ؘ���F�(Ϗ���Y.���	Uc�P�/쾫�/'�/��>��:~��/��ʱ�ޡw�f�+�Ӥ�|��S���ͦ�g(��*ϰ�p��k��t��@O\=C�U��&  w  H�����ܩ�-�t�)�u!��u�]���_JP�q����	k^�Ѷ��(��*�qQ�G�cs~���
6~���f�T�y����2�nS�ҝ$^��'����zc���,YK�(Z�3���m���� kgؕ�V��{-�Aw�ͽ����ѽ�t�Y�pj��}W/0
  ���&KF[Zc���h�^�r�D     `8�k�zݬM��&��  
�9�����X�A�9*����b1V�՞������d�C�՞�Y��8�;�d���(��γ}�,?^�*��}.���:�H�˶���Wv�^1�*�����%�9��k���b��ap9֮�G����KZݻ�Y|,�
��0�3l4
T]��O���&/����Suk�_k   Ip ��8�?O_;פ���T[�S�����He#���� ۽-���q!Rk;?	*q�dm���ڇ[��;7���$��ɖ����n�=������DmZ��%�J<O�����D+OP='oi��X�&Y�=�c*�����V��v7���,Ch������xI#C��~���N�����S�z�͠� �a�Z�m;�z}˯�tvb�     �p2w����M،  `B!���^����mj,֩P(z}C��XZ�={V}�y�F�=�=D�kk�Z�=p��X(����,Ȋ~O�'���x��7��vw}@�����G�e�a�׽r,�{�O�b7����cyW�nݛ��Q�F��w�*��/n-ޢ�-�Ɓs��7Z�4  H��  �)�^���}k�[�M*�K�0�J�r/f�E*Y�BP�]���\��%N�!	���T�T�%o�5Q*�@{RBԠ����I�J�{������63�|�16L|��%�*�ٿyK�R9�h����d�Tp�]�����+7��ig�6�Wn��7�p��
�����"=�_�g:G?�]��� �c���~o�H���V��?7��;    �3??o4����y4� �6Ϝ+���}�X^��b��ڮ�[�ի={}�0�0Jk;��u
���C���5�P��1I��;'μ��3l���vq���h� +j�=���F��?n�Y����@����u7��0ms��cy}����+@{��n��^����<C�ݽr��t��w� �͟��nah  ���;  X�+��@c�6�6i�X���1�p��P�6*�S=�J-D�B���s�hI��+L���ݯ��D�#P��-@��v�M�'�R�1}�L�$�)��q�)��6�'�1��T���m
Xz�7���N�{N�����	Y&��NWp��"�.S���x�5}��v�����fw^�p�2K�,R��9z��5v  2�ݪA�}~���     ����5�V�Fs�m�W�  ̃'J���eZ[���b����IWyWz�	���P]�%��ʱ��ʱ�	�nw���Ϣ��q�c�g����:� ��sE��ldE��,�������{L����E���\S{�G�zC�U�U+@˂�U�U�a7̮���momё�5z�����1�xAw  pA�  ,p�x��9�LkKTwĩ1O��/P�.��܋eU�=�u���E�\�8r����$�N:�T���a�C� ���FU�r�0�%J��+J�=lޠ�]�
:&{-�'�hi�U758"��L��W��|~�	���W�6����(\�{o�#ri53���Vw7��y?�{n�}�L���7�!Z ���Z�s��X~���S�N     .�ݻg<�N#  q�@��zf�����R��U�a�K����D�����;4^�|~��3�P�p�z�=k��$��(�
f���(�|��P��'4�T���x^�l���}r�WH��2�0(�������\_н}�ݛ�~a�b,�g��1�����ڬ�����eZ��7�  �  ��`9Ozq��뭋ͼ#N�[ڃ���KJ��`%��u�)�@ej�-L��-D��(X�=��L�ƙccn��</6E)���le�1>�F�$�4�+W�j�X���1ꦆ�h�+okjenhP�ܽA�f�ɽ�iro:��w:"Tgi��p����/��U���w�շ��H��x��V9L�Wt ��z�V[�ᒞ�>;;��;    �2{����*,F  �Q�}�j���7����b%��m�OX����J�0�?���j��U~a��H4�����c�u|�9I�c��K��_��|���b9V�^���_��7Z���x���@�{���;{�;J�p�skR���y��W(~�hhc�.}i�5�����ֹv��e  �P�   ��.�p�H����ؠR�$�dK�D)پn�F�=L���S��vY���s�?�����/F%���*��(��γ}�ax̸�lp�����T��gY�
;�䱰��������
L��$�T*�*H�
oh�od���K��+'��iuw���~�{l�r����'���Uk�����H�.T������m5��5	 0Zpp���m��sss���     ����2U�U�9+�y�6�  ��g��Rn�6*Uʳ78���.�Uav{�a��h����p;���kkO�#���2О��wn�eL��,de�'�g���$�%ƙ#�����$~!u����bI�B��u<��{�Q��9i�]������r�G����ϰ��
�-�L�_�?H����u ��G  0�ON����Z[Z��R�ʝ�1�n�����"U�`�q�]7�N*a*,��&�԰�ړ����:���A�7���y������
Z&b�^����Α헷4���Wъ�_�bqjW��.ޏto73t*W��������~���ze��}j?-�'�i�� ǝZ�����������s     ���;w���`/ ��ġ}����O�v�䴶���y�bs���n!خ�!��/���ů�$�Ο��{��a���y<���a2�tl��Q�$q�,>VZ�(��}^�(Ȋb�;6ʸ$ʳlx�6<�x~����G���x�<������{��A��_�#c9^a�7T�bɼC�R,޷��A��8+@�j�0ͮ�3 �-�@ �&G���O/ԩ6�j�BwIA����*W���{�T�68ОD�=�0�� ��=��{�sm�1g:6����:ϰ>>cC��c�s�<~a*h��*��%-P�O��A�_�\�X�\{�+RyD+�pUp���V��<���7;�UG�������p���t�W�m{{��kS������1�Z�h H��Z�����rA�avvw    �!�?�޽w�x���   *r��+9�/MSm)Gc�����m���a_����c
+>Sp�]ԇ���x���H���1�m�1g:6�s�<�����K�=V�aМ8�⠼°�s��e����D��w�#����������0�нt�z���_X��&�f'����,�������A������S�
=3y�~<M�� �G@�  B(�.l�z9O�o�f�A�r9r�=�y���B�^a�_��lW.%nwft�o����6��2Ԟ�`���8s�8G���~��Ay�Ǐ#L��7�d��MbL����9���{����{W`���|�U<�Jv��3������ �J����/����zhg��|�<�d�Hխ�y] d��+)ݬ���z-�J�677i߾}     ��������&��9Z��  �u��X���YڪlR^����~�Prw�A����w�P��o��u���[�O���ˠ�ä���9&�qQ�ǝ��y���Q�Y���s�U�e+�n3Ȯgc���4���M�}�<>�W�������:�.z��q�*Ў7�ms��݃ݍ��+@�+L�k��r �>� @ O�)҃������z�,yZ�*�J#���������.'(��ۥ���B�,�ޙB$]>О05*�TZ���8ӱQ�ۚ�乒$�H�$&ϟ���gN[�2�E�*�M!Jg�nK�?Ԟ�6���{~���ū�>�=�h��ۼ���{W�j�V����:A��"�ݬܡ����9ze�  =��S7�ί�333���     �67[�m�\_/S�/� �hs�X��=�Jk������<ĠP{��(6���u
��Z+>���!���&�����6�$=6����:gV���F�/�S��Q<B�<�X��M�OL��*�1>��/l����X�~��R�+��*�Ck���?t��V���ݝ�i�ѽ�]���t}{��4�ыWO�k����r�  `TA�  $���/6�6?M[�"���)�t��%���b��`$L��������(�+L���IZ�ګ�U㢎�:'�s�����}�	��|�q�)�s����G��&P��M��A�_|?�2�v$Z�[�h���V�foN^&Z9�M�/���	Vݠ����	�V��<v|s�^�z�^���+� �g�V�Z#G�E�뗙[�hrr�y�     ٤V�9��¿�  {�}E��w�h{�:�V�4&x���P�7+�r��!eXւ��v"��:����_��='α4��1g:6����>�0}q|�0t��!n >J�=�Oh2v^a��$�%�z���^<~�?�������{�g��	ۛ�
�'���7�;+C�aX1V�
���{me�>�_��&/�On���k"  �w  ��K
�ؾC��m*����Z��
T�օ��v����ۉT�Tz��dǙ��2���4�7��>G��X\a*���)��I�v�!^����Gb=�Q�xt�V2�J*Z���f'�����۝��f&gS��{D�B����@��
 �0�
3S-ѣG�Zܷ���޽{t��Y     �dzz�X3Z����~� ��xz�H���hs���K��b,�r,���5�����������̘6��I�?L�#L#�>H1���sl�Թ����5,��=�;�G���T�=-�P6��x������sN�VNr'
�y�����'���]������7��cicI�AO�S�ը��wN�۹��Ɲ: �(��;  t�x�@�?�BkKj��K
bT��������v_�n{�J��la*k�����(c���:'�sd�&�%��|��t�a*j��lއ]�����3�d��Oнs�v×"����OW�R��{E�fG�b�jG*\�awU�]��lk��T���_�=@���{hs $��5���3��M�    2
�}��i�� �'�����p��Ţ�;+��.��>�t�g�p�l������(�'��������o����9&�qq�ę�����ϝ�vn�a�96���qQ=G�s�=����_�<��'�3�.z�;;�^��
;�v{;{��^�W���W�չ��ɶ��D}{�h\��ON��f��bm�  `@� ��)剾~�uA�4M��\�8�h`��˖�S*aJr��d���p��?�`� �����G�ccn��6�>Q��q���sD�l��mއY��3�/39�i���rbC�VKC�P����[��{��7;�j�+Q�jݻf�D���ؤ��=49A/��G˛�  ���,��v����^c���iee��9B      [ܙ�u>�����Vp �r�]z�r�VoSm�A�������՞��MJ��}����s�����1I��Y��8nsL�cm̳5?+�����":ϕ�c����E���f�+;�T��̶_���������n�]r�ݕ��M�B�
�j��=G�K(��f�D+�
*�r�k�s�܁<m��@?��t<T  fp �i��(҃�9ڨT)/��K6�|�T�����ڷ���r�{=��*�qQ�ǝ��y��qu�+B����&�t�4ĩ��Q��Q�����_O��of����0�����w�7�s�}g'/���uG��,A(��ogP	V�h���%Z�8G?��$  �͵�2}�Ħ���7n�g�z�     @v�Ͻ�����fkE�6�  �ΕcE�ܑeZ]�Юo�gU1�y�=x�gY1VP�=�`��g��fq�cIε=�d���8sl�M�\�H���ԏ��͏�-����&x79����U�}��tw���D�Aw�Wt����ao�gO9�b�g�b,Y9V��=.ޠ��x��^;NS�X 0� � ؓ�_�?=�M����-[R0��ݸyA��^��t�T�T�@E�P�T��g����S!V16��4��Y��?�q�c�̱9?��f��?_����cfE����+d�-P�O+��?f{��w�� չ�tW	U����������u�n�{�#`���M-�JK�r� l�-/]��_>N�[9F7� Z �1�V���o�^w��߻w�֫U:x�     �lp��]����L�_v �Qf_���/�+ש��o{�
�P��=ĶW������v�R,�@{r�v�R,��A����8�;&�qQ�ǝg�Y|����ʰ���+�G6�v�]w��8����q��(s��e�)d5hw���{P9V�_���՟���>����h����ʱ6�W顝%���Ezi:G۰ C� �=�W.���-ڬ4�\.K�%!�.��6/t�TS���V�ݽO��~A*���x�L�Fw^��C߇-�I���`�}�8e2vU�q��������L���`Et������ɖl6s]!Klgh��bU�+^��Un�])Z��,Z���c�%z���������k' `��n���TKt�P]k<�f^�~�>��     _�]��2����ѝ� ����E:Ӝ���&�d������r��J����3�{��X:�a�`�^s�K�|�4�øs��dL�c���=?�sQ�(�d�c�3�G��g�+��m{��1I{�6��/�?�[���۞a/��{����O�d5]����궹oVnѷO��͝3��]�� �� �=������-L�N�D山^�=D�
�K����v�0�,0�.�ڥ"?v��Y��$X�8ns�ɸ��α9P�N
��s������{n��T�<�Av�qY������NQ�'t��	U�6��������.���Tb��ʠ�İ;�o,N�__<Bo�=�% V��N݀;3;;K�>H���     ������ϛZ+�Eӕ   ����vn��秩Q*yW|ho�/��-���p{X�]�?�`{V��$C�i��Mƙ��2>�3,�DT�O���h�A�����)��
�Ρ{~�c��#��B�O(�$����w�_�:��7����W}�ns�׷��Tc��v��ϭ2�m�  � �_�\�#�[T]l��ؾ�P�I��^����=�}Ad�m]�X�=������x:�m�1g:6�x[s�<�^����%L��f�=� �\�U��$�(�9&��j�AwjU�	�{����wX��_��	U͐Fw_�]�a�X�'Z	b�����6�����z|�"��u�:4+ @�6
��]�#��x~�q�=���     �����sZ�|铕 ���%:�}�6��`{�/,x�a��'���
�=�|���	���^)��H�P{�`�0�����8�l�9�d���8sl�O������%$��:�~7�����
Î�y,K>�lp�]~Wݩ?���ʱ�<�|~����|�X�����.msWc�x�^8Z���E��-�"  � F����:�-�'�A����Z�����8%�%N!���l�9&�6�ٚ���4Q�([�Tй��G��ƚ�O:c!`%9�fx]��Aw���n#�6~��d�UO�R�34���P�#V����B�����'V��Uo��Wf�g҇[���y�� ���r��pJ/���ܺEW�\A�;    � �w����ϛY/R��'  ���ӟ�ߦ�b�gE1V����՞mc)�C�`�M/p��C�c�u���I��I|?q�>L�o��'jx=h~o�f�]5����iK�/T��k-辻���c�x��'�����������kc����׍z��}B/>x�^���4c �� ���im��Pme�/�^*�7/����@�Rk;��T���ܳl�05�U�uǘ�3g���i�o�򜘊da��D�]5/n�]66�U�qSQ)�����s���"�x,�����KE�]uC�i;�Y�{�O�R53���f���%ݷ77�rs���H�u#O�&^; �\_-�Ƿ�@Q����?���z�     @�8�c�|i��e �Q��ã�ڨ4W|.u���u������b,R��͂�=?�I����f�#̊?��7���hc���o����u����u��Q�ŨAv��$�D[~`ǲ���[�S�C�{�A�X�_h��V|�hs-ƒ��|��4O�*��������  �w ��q�`��rj�����r��Pa�f�v_�}��$���߹7�`�����*X%1.����l�#��e�8B��-Q*�|I�m�u�R����%D��?��;u�
AwͰ�_�R����z��f�fG�
hs���V*�J<.63x� ���Y�Eߝ8H�O�{sX� `F�Ռ>^��<��=��{tee��9B      ]xE���u�y�6���Y   vN�����h�2G�A+>_�����&����!��T��s��ilf�p=�Ax��c���57�s�:�ϕ�5�6?)��d� �°�I�_��o:6�ߚ�C�y
��!���{��Ϣ���V�����g��9^_P��S���=��B�ց�)z�����w�i��6w @�@� 02�r����"\���ݶ8l/4/�	��Ĩ��8�T�°���FU�Jb���8sl�M�Y'��%�Xq����&��l|\!k�*�����kt���t����`�mso
�U���/���Ukk�բ�W��2�����~��	=4y�^���6�  |�R�ǏmQ9�=��G�>�y     ����]�i�Kho ?Nk{�Ֆ��+>b��>����J���Ty�}�����^Ϣh�I��:>�$Α��Q�@��F�1�����A�z�q�@���i��ǒ�U���u���x=D�^g2�H��{�����{�&m���a.��Z��X�����U�����@�,�ʩ��4C @v@� 0L*ЗO���R�i^(�K�p�/�Դ ]RP&P��c���@�+N�.Ȃ�D�Ez2��,	S�"J��l��26����:ϰ<������-aJ5?)q�d�	TA���w�Yн;��B��Q�����n؝H�aX��me��W��@���:�ج��<KJ���}���;g�[��y�V  =�׮��=vt[{���"����ɓ'	     �Í7hkk�x��V�fkho /g�����w��;��*خn���{�^�P�!�����ڳlϚO�5�P��1&�L�Fokn�v�<��d�cD�����mޣx���H�/��h��t��	��P��1��sꕟ�-�'���6��v�{�^�0'������r(�����6�_�;@��& ��A� 0�|�R��nRmu�ۼ���=�
�5/x��~AJ��nE��T�u�tnG!�E,�`���8slηu����fw�r�����l���T�׻m�|+3
y���e�������v~��q��ྦ�X��o�>g�q<�Ƕ_o��ƨ!�$�������� ��(Tⱸ�����W��t��%�w�vQJzw���uA�D�_�r�\�`%�7�FO[�����k�՝�N����Z���v� 0�|�\���ԩ�ӿ���'ND�     ���u�ƍHs�[����  �e���pu��+;��vU1VXV��Ϯ�(��c�o��C�/�"
���٠}&c����۞v,��6�$=��<������������>^T�0hn>�j���3&k^b�~�j�iP=���~���f�]��� ��۾�,���~��3t�c�m�__��.ҫ3(� � C˱�y���Z[�I��.�ۃ�)�8Ծ k^�	TV�)�@E$���.���Y� X�3.�8󢜇C�Z����hyyٹϦ�򶾾N�j����֜muu�9��y���t?��r�����?�9r�y���� ��C������[�>���ǝ1�;v��x��{L]�SA�M��6��q�.P����l���Αl�].d���9�N�-��ngP�Y2�*H��uD+1�rw�)�*q|�r�������q�YA3  �Z#O�����5��^�z�     @�|���/Y���]��� ��!z��R�����+>����
/Qj�c���J��H�?0�/؞�'8J�a�sm�1g:6�sm���A�gdo�7���,�u��X��9~x�Z!�6s��������5�=?>��5�~��{~|���q�x?o&D	Ǉ=�Iy��yI�ޓ
��O�K�9ǆ��/4kt繒����B�~0�Cnr�����{�TM�~��љV����N��'��On���� � @� 0�<{�Dg�����߼�ڮng�I��jkl�
��\�"
n]@�=[��a��-Z���?�q(j~~���t�������h�c�J���b��I�j���l[��|a���k��O�<I<��x�ۣG���Ç�[�?~�Μ9����Iq�)��&��l|\!+m�*��cqC�I��M���wG�L��i-C(��BU�~�p%�r���&��z��5B�+�ڣ 	������5z��J�^�L�s!w @0��9y�N���u�'׮��Ąc�    �d`�lnn.�ܷ+c4X  �i{����X�x�~�н���A�=��:�v�j����
��be1�n��tx=Ip�=�(���3=��������'�X�",��7q�f߳�b,?��s~�,���㍿f=�-�r�𼟏�/Ȟ!�[=�$o�#�g;Ȯ;�tL��z��4��c6�B�s�����=��z�F��{���H����/krov
���
�P,�<CeI�F1o��{���e��;Oo��	  �w �P������˻�Y�F;��q�]-VS�`�\��.h7/P�0.J��T̰�^�j�}����(����>n?���ݻw��u6�x���ܹC�o�v�t��
��ysŹ������Z�b֩S��ĉt��9�k�8 �x��&b�ߓ�L�B�
;�V�]gNRb���t���[�`E�̠
����knmq��2�*ߚ���['���U�e�w�������������Յ#toAw ���f���R�O�"]�5��ߧ�=�     �4[�!�z+
��ݩ  ����<}��6�n�NQ���a�������Cu�����څ-�lwoU���ۓ�	��?�{�$Ǚ��3Gg>kK\ru��}gs��n����~|�o]_���x����0 >_����£� /k�w��~�R,wc?�����<�cϐ=B�UAx� |�P5��WL;��o��%��m��6��݃猪��"4�����c�՟E߰�*���&��V�ů����'/�K�y�n  �� ���S���pq�6kT*��"T_�=��]���Z��
T���ym��T�
���FI�ʒ`e��1&㢎W��d��:��YT���u��u떳���
^�n[|Pc<��r��N ��ٳ��,p�>�d�I�SA�GM�29�t��t��{w�lBU�Gw����+q_�~�h%ib�u6�5���]���V������x����  r>X*��G��l���4�޿O�[�     �.�>��666"���v��B  ��wȅ7*����|Cي�E�+�_�Y�+�7�y�ʍ��~/�~�=Ͱ� �☍�cLƙ��2>l���ݻ����Oq`����
5|�oYO��h~.9υc����~�;}����-�ŕ�����k��aߋ�8>�jl�qA���9�z�6|D��%���&��=J����y���W������W��w����0����=CI1o[�w�;g��[���H� �w @�)找u��^�F��R�@Լ.P�� QJּ`n���i]t�=���A	V6ǘ�3���͛7���&�y}ff�	�Cp-����xs��@�-,lq�������;}������-qJ6�f�=��v����qC�Q�S��}ϥ�����%��D+�k�h%��>��|�$T���s��󸃫����g�'��hmk�  @d��:���=u|�h�{�Gǟ^it     sVVW���t��sE��� �}�;���D;��i�Y�;�uJ��0�d�goQ��K��s�p;�t?��::�2��k�Y�#�nv���qQǫ氷��u��Cd���|;ݺ��¬�����N�7��;� ��/^tJ���;���{͊|O*��+���h�X�}Ĥ���T�;$�� ����r�w�P��W��Eo��)�6�g�����2�p{s��6���K���.5w��� �d�J �4W���ZY�Ri���.	���T�@%���`�b�i^0
��\���S���+�>(a
�U8qE+^��C�lf��߸q�����M�,NT�U{�7�M�����c��}��%�z��s��Z���Ç�E�8�j�iP]gL�*�x�@�Μ8���I&c�	����"U ��'�$Z��uD���{���`���}��<m������4M���hf  x�p�L����`I��`�z���ߧ��z�     @|�s�;��ܚ���JoΏ  d���3]��3��!����o�g�K���W{v��ڃVy�n��߆�˲}�����9&�qAs��daa��9���E�#�}��<��j5�~����_�i���~��𻸱G�-�&�����8�wcl��I��h3�n:?hLп��"�
�Dҍ��������]�Ք����y�g����!~a���ze����Q���1���$  H
� ��O/h��ڨ�hll,P��o�*g�Y�]'ܮ/R�O,J�}���{��='α4��1'��8����wC켱 �K�n�v횳��)��փ>贼s����rn��\$��{*�ɱ(������ݻGq*���]J%T�[�u��^r�+Zy��v7��mm�\gS53�VA�_���Ls��r�2�4��f @��K�U�G_9S3�7{�.�>s�&Z     ��?��)���'�%Z�.  d��w�@���Q�K�COQ��7�~��.[�9�?���7�����]�f�S�o{N�c6��cc,}��}�7d?����Od����/ߡ����G�&¯ytg�71�~��	��{�P56	?��� ��cI��Q����a�t�t���w�+@�eY2�P|W��εD�x>���m�����Xk��da��|�~6��;  p d�c9�օ-Z[�Ky�T�!U�}Ik{Q*N�/+n�݀��(ۓ����"X���E��=���O>��i�d�D� *�o�����¯����裏:��'''��s�P�8Av�q�,PKb�������E+7�޾���$�_+�VA-��}ϵH>��Ag���%���v3�M���������5�V �63�E�[+�ĸ��_k?v�	'     �h,.-���t��[�ϖ�Tp- �.�����gk�V����w���l�n����S�U�j��������q\w��8����m����|�>�d�������$x{�W�}�k#���X\�u����-���$z�Wv���A��QǦ��}/&���]���
�=oP�t���}��7Ty�&�X|�F�N���������U��>  �� �L���"=R�K���n�B�#T�(P�S������rq�+L�8a*P�"��G��+NeM�ʚ05��U�q�a�C�~��#>qC;�����*D(�)�����
��������#/a����#�<�Z������v�=��x,��eHW�Ϻp��Ztw��=\���+]�*L���$����(R����o}���zf�U�^�_ߪ  0o.�o_�R���%�}���駟}�     ���?�����?,�9!w  �"O�.�d�U����CU�=,��kn/����E[�Y�!�z�n���ݒd���m�xix�Y�m�#�8n�f���\J��?��>��g��� -\/�������_��{�СC��9���X�'B���sd�+��19>�~��9�������o{?��o�s$h��5�N�=�7l6��1�0��u|����]7��)�ꌩ.�џ/���s�ν �-p d�\n��������N��cc}��[�`{Ѹ�=8خӺ�#R�n���ĩ���m�������cq�&9���b�@;���y�ZXX�,�����Y\����l�v<x�>��O;"/Y�B[�Z�#,�6��,����e26�}j�ʹG��ΐ�h���xz�n��+J)����J�
Z�����k�������}�Q��	 {���<}�R�G�l͛��Y�����     �x���$
|���J�   kr���y%�kT/��v�g��y�����`{���������C�:x��Q�'��h�x�q��.{�b��-����$ ����Z�O��\��� �r9���,ǲ�T�]g�m�0�Yۧ�7B+@wW��c��e�a{���.��=�X�m�Awɭ�#�-���۹A�&/�O5��  ₀; `��<P�N��Z�"oj�50�7�X�k^nmW�.�ǂD��%�"����)BJ�JS�JC�2�6D����w�	���`T������_���ǯ�.\�'�x�{�1G���,p��TQ���H3�WԲ)h��'j������T�D+U�]&X�m��}�zD��
�����9�hU[��o�>H��N��"� ����2F�i��g��|Ժn=r�;v�     ��K�w�܉4���^����ٔ   S�<����^���"�Je�gh���}�@uV|nߏ��}DF�CtI��`���zV=�$<D����������o�M�����x ����_��Սxc�5��ɓN{��rQ��Ą��5��g�+;��|R~���A��|d�tw���u�A�#7ݐ;_s���*߰���X^��N�*��X|NW�LӋW��/���udS  �@� 0P�9W�s�[T]mP�\V�S%�@���_��_ZP-N��v�p�,��1*q�w�Ɩ85,��A��GE��߈�e9���G�k���Q�j�
A
�Y����̌����K��0�۹��g��Gy�>����ѣG�sl��ecvOJԲ!heI��2/L�ᱲ`�J�
�\�J��]lr��=��h����s9�h��Y�G�=������^f��z������	�Q~�{����/?����     ë5~��G���\��� �,���"=�y�j+M��Ͼ�,c�P����������C4/��R�=K>a��a�s��a��]�yjj��z�-����� �;g����_w6�_[yh.�b����w�B~�pI�+;���8(�P�?��A��ecڷ�/�;�]�Y�7l��e�X�1o�{^����Y�U]Y�/\�;G�ӛwP� �� ��Pl]�}�*���5j�>$pxAG�
j`��ڋ���`q�+T�
T:Bӻ%�>�8eS8ڋ��Q����9��R����hii�  ���#��#.Y��C�T�O>�Y�>���=ֆ�eS��r,��g\1�dl����<��{�p�RT^�tB�m�J\~P��.6��r����U���U}��x��|� -m ��^�v�H7�Kt�`�h�Ӱ���٧�6z]    �k�篷�~�h0�V����  �B�H��+M�X�I��Rh1�?Ю�zC�E��vY�]�;T����]�9K!�a�	m��Q�i�_'p��]��׿���!�����_�_������C��SO=�ln������s��
Îۘk3���8(o0ʾ�1��n�]~��d+@�J��0�����o�X�m�9o��p�t�q���x�ɭ)�����^/R��^  ~p ��ġ=w|���O��O����eb��l`W��t�T��&�_�bT"Uĩ���6�4ħ����b/���o�;�C��.mllh�Z �`��������~���v||�;޶@v<!���m�Qq�'j��q�V�Vw��{��=��+Z��D+���J����{�t�./����Ã��<� ث�v~��ߠ}��U^"�ͥ��I     r����V3[1G�7�����_( d�+ǋ����QY�R���U�X���xޡx_�z�wt�0����3I{��ld�}�tǈ��/d�������۴�� M��
����+�8Áw^������}��s�z��16��6Ι��dlZ�L�������C�O�l�v�5tV�*���M����7�
�B,�/��;�W��k����r�  �� ���D��7o��z����zbTH�=�}A��.n*QJ���j�YV�	��D����~[cm�:'�9M��-/��r����^�J�B �����=������g�q������-P��hיg�����|[�vq��hŻ5��h��T|�F
�J|<qs��p՞���p���`�]�0���>U��_��／�]ٹN�'/�_C�; {���k�����3��s?�v�i���      �壏>r~)0*�WK4[�E �_�T���7h���ry��3������E���;4)ƒ�7��0�Ŗ/8ja�4���q�iyu�7�|�	������!��=��������1\�Łw�	��C��~��I�L�XV�B��Y
��橂��Vd����5��%��ۥXM�o�b��=�0�R��'��	�K��[�
е�}��N�.^�_͠ ��+ @*�r���s�X�F;Ţ|Y���es{�0�me���┩@����Vf�]�:�>�}Y�?�c�㋋������ij��o~��!F0x���������'N8aw��_����w����ε9'�~A+������}��V�k��n�VwY�=��]&\�Ʒ���҃��w!�����w�h%�U|�W�/ܠ''�G3cT��{ {��e��ޠ��Dk~��û�:� =z�     @�۷o��7"ϯ6r���> �AS�}��.m,\�|���cI��cx���v��E����[^�0x���۞��q�eϐWyf����_w<E @z��I�������6{�����f��}�st���@o(	?�Ʊ�}Ĩ~��ؤ�����
Y���	�-,��{\y�{{�[��in����]�P��ʱ�V�n��txm������S�� �� ��9�?O_?�F�J/�.6��,+(�D!���L�T5/�*y�]�xA�ʊ0�Q�D�����v�_��W�ҁ� �v ��������^z��������/~�Nk�X�~�"�nS���?�A�������J��w�6�!��kg�q���N^����b�ΐ�tﷶ��}���]��XD3 {����ӷ��i�dv�˿��ޢ��%��     {���%z���#�竱����N�  `�L*�s����괶����+���l���|D-�0g��s�� |���n��0����4�s9�� �����������˗�r��|�3N9��Ç�ー���IK�G4	�g1�n�C���A���|�S���
���{�a�����A�>��/�$��f���ţ���1�[o  ��;  Q?U��
w���E�1G��5����m]A�ؿ��Z��k^�ol��S�J�b�D�Q� X���fA�������,� 1����?v���t��!�җ�DO?�4=��s411�kK��������N��q�+bV�B��J)X�uʮy��J�r�,�`��.Ch"X���`��A���K�.�/n"��^b��������s�֧$��^^E�C�l
xV    �=
k�|]'����ݫ  �3�Jt�1C�M�(��M��D1-�P,y��'��D����O�1��9lωsL<η�����\�š���M d��{��g��輿�Oȁw.�z���r%��.i����U�����Mƴoy��;�!���6w�TY�9����6w��Ϯ_蹶�byW�z��6w�_ع_[[�Ϗ��쑋��x�  5� �ϯ橸|�;��@�X^P��=P��1aJո��]����)ه��ĩ,�س"LeQ�⥃9���;��+���.  F���������c�=�S���x�`��?�����ZI�mݳj���V�[�h�\��s>�6��҃�K��UO��r��UN4�$M��z���L��N����Q�z���^an�@�/��SǶ�箬����|�Y)%��;    � ����F�z�o�R�,�*e �A���ҷ�Qc��J�U�����a�������ü� �Pk�gwe�;�9/�F�o{N�1�8���Ρv�>��й �����������իN�;�\��V�v���4�B��6�%9�F�"R��ܥmR~gGZ�Em���^�н���]��t�y��a�X������)���K��T���� ���; �:�r��󛴾x���r�eA�ܮ#P� ����(N�"��q�T�
�*H�b��g)Ğ%aj�v��6g�x���B� {�`�+6��O��Ot��ez��睶��~�����f�=��i�)dE���Pq���ݑ�:��ab���� l�if�������y����w����[<Fwװ�  {�?,�љ�:�����B�Bx�]z��'	    `/���~��T�V��c�W�����#  ����g��h����l�lnW�����=C3�PԹt�C&kޡ�y&���?��q���+��o���y��/~AKKK mfff��������������}��_�'N8c���G4	�:��<՘0��G�dw7YA�x^�����=��)��o���,]�Y���s=���c�ze����	z��AZڈ�b `4A� `��
�ľ9�.mP�<������۽K�T��vUk����S�~�	��]�J3؞��d#����:������4==������ ����wy���t��G��;����äh���ߦp5�}��b��˾���Ű�x$�s���*�.�w+Yؽ��J�ۿN����  {��������OߺX�r~�L���m�����    ���no��&����8K�^��O��X	 0��(���;T[�SylL��cu|R�D�C�Ȅ��M��$�؜g�/�Q�۞�?v��z��W�@;{���nm��r n�u�W�~�嗝�����B,.���W�BgϞ�E�P���bV<��-�i߲7�+��[��O�
}��&m�=�p��/��cuW�_�_C�
����3\Y��[�?:Gܯ  � � ��/���i�n}w��T���=\�R�f������SY
�gI�JJ�����z�~���:������ �˽{��?����p��qG�z��gk||�cC��#j��oK��j�]ܗ�hE�%�^��_���;�]a�#^u�)��W�`�����x	^^~�;��m� 0ڬ7��ʽq�����+��u3���>o>��C    0��縷�{Z�����R�n�� �oN�*S�,�P�j���W���ڶw(jZ:�!pg�x|{)�>(�0���͛7�P�3n�  loo�k���l��OO>�$}��_v�|�;.�@��~�j��$�z���]��+��u�܃�����r�^)V�z�BUΪ/�.��s�6��v�.�L���W��c�g @(Z ��Z�yp��+�(W,�>�+Z�c
T��3�*(����/V�Mq*�`{�ι�B�w����g?sD����#� ��~���o��lG�q�ݟ{�9'�>66�KR���?�j�l��m�V<�=�c\QJ%VqSu�iTb����to��*��!/�U��&�6w�`%�V����3��7˴�2w F�{���8FOߌ4��kלא��I    E�p;�qp��*� ҧ\$��KuZ_��z�2�0�?W{�}T���w(���+>��C&-�0+~b��m�;�o?��cz����7���S�%�  q������{��y{�ᇻ��zQ��#*��8b���d���ή^���;����t�A�0�Py��ks�b���������?n���D��� �X�ѷ��h�2O�R��v}��]>0L�R],�m^�^T�ɒ85������8��+J���?����t��]�� ����B����lǎ������hיc;�v���&ъ���w��E�J&V�53�!��@�W��k��EcP��Ks��3��'��2� u�[,ѱr�.����ǟ|�Ρ�    �_�p�}nn.�y��<�:7�����   ��8���V����w�J�t���������۳��I��Ohc����s�����_v6�� ���|���������裏�/��x�:a���B�~[~���$C��8ct���� �~�f�{P�]'��^��"�j�g�5VP����]�ޅ#����4_�/���A� �+ǋ���UW6����*G�*���*�p��8%knW7/�E*&-1*+BԠE�4���n߾�R?�я�
�  M�������ߝ�ĉ�o|���~�i�=��z��Eݟ�p��P��/+��qE)�X�ii �Vv�  ��IDAT�'��A'��煦v�A�����[U�Ly�&�]�7�D� ���6�����t�M��&w~]{�G    `��ro����lno�����i��p;  ]��(��۴Qkt�C�K�:R�](�����a�ޡ��ݽl�=+a����:G�9����*ϯ��
���� ���/~���q؝�P.��ַ�E�ϟw�������uΑ�����h�Cl��Dާ��뷹������ð�{^�N2X���-��o���nЍ����9x� �Up D��tb�&mmR/�..%hԾ���Tr��w,H����$�a��j�v����g�(��o:�> ��g�L��(�{�5���	 �'>|����(��SA��G�����9�P$@Y������d���쓙��{f��_uWwUuUuuwUWu��y���j��!�]}����imm�C=��~3gΔ��g�}6����v�WN�Q��[�1/�V�뎴H���L�J�msM����|�lAw���!w��9N7�7���q8�bbo=Ο7OփR��_�^�W��g�Q��n�h�`ȝB!%�n�݂��������h���B�əs�v6a��Wc��ڮ��Y�!�������;tr;�+���Wnkoo�ڵk��/�7ޠH):�ۑ��w�u>��Haw�N�0Aڧ��r��~a�s8y�ۡv+��#_h�A=��ܕM�F>a�����/Pk˱��R���m��%�b�P�̙����K�H�wBHN�@��u~�5�����d[�]ZAe��,8����H����E*����^���0%�`͚5RS���D@!^D�n�ڵK�.��wߍ�?g�u�v;v�����\ǝ��sB �C��ҳ!v�wY�R�U�&w���rL)L%<�ĵPF;CR�ʧ�!��L��._�E�v��yS�ĎJ�|%�x��A?���W��"���o]L�-^���?�B!����������V��i�®����
��pN=�{��H��9�b�ǳ�bi}B����������[�ͼC�1/y�v������
=__֭['c�������g�7�|SZn��v�x�8��Sq�i����Z��K~�Ѹ�Aw����b{�F�����{:�.y��8�*���"�����1�R��O�_}M����u�k�h��z��͛�U�AD��R�P�"�X��sg������q�r�n&E)�H�mZA�p�^�ݯ���LE����y\�c���l\�&��[���ó�>���BH)!^�6m�$-��v�$^�q��x%ޓ��H���C���0����z$-R����(�ܵM�JqJy-��������u3q��E+����q��Qx�k"�t����r�m ���q���k@~�عS�0�/}�K|^$�B)D��[o��C�|�;+�Qg!�XL���ûn�DeeeF)��G4�[+�Jl7���;tr��ٱo!����ￏիW�g�AWW!�����J�K�妛n��e�/��^(�n��h�ioPw�Wt�C�v�g��^���/YP\�������E	�I�PO�K�+z�2�s�5����}?��WZơ%̔;!#�	!��1.�ϏnA�#��V0ש�vՔ��Tb[B��o^�
TzA�l�T�H�/L���mq�k"T������矗D�>� �R(ū3f��sϕ�$�����[�r�E��g_/R�1;E�|E,���9 y��)������ٚ�E�!�v��z������p����)3��@���dO8����¤���q ~�?�a>��Ϣ"�E/B!�/���#��E;l���	ack%!�X̟�Q���=Iy��J��}D�p{01n��۳�����u���k̎}߿��>��hhh0ܟB���RΊ+���#���B�N�6M��_h4^���H��=C9���˾��K�ŵO,]�������g�cY��f�ֽFS����n��>��F��a�tl9Hϐ�� �?%�ٱ����;�.o�nO/ZqJ-T�R�q�0e2��@_���y��Av/�Zv��9�)�D��$��;{����%K����]j�=��p�9砦�FڞK��h�T�+'�s����O�H����+��63��W_3iŪt;C6a*�%c��hӢ�0g^jb�;!�J}W�C8n|$�sttvJ�����gQ]UB!����ny��w���#�����`�R,N�DEg�w��f+�2��ޢ�Y���C�z�N��>^�c_+��/\�f^x��]�V�!	!�\ؾ}���u�]8�䓥��)��"�w�������R�՞�>�d��XT~a� K.ǒϧ��c"̞��!wq�<�Ae�ݤK�W�n���s���AB��	!��2;�Q=M��3��Z��,�^X��xZA���D)�"�aa�v�Qn�S�"B�+L8p@jj_�l��$����x-ܴi���~��8��3�`�w�q�v+�s��R���;-Z��k�;�IY� %�*E��$V)���T
V�qy�AI�RW��V�\E,�*�ш�G���� ��!�ͦ�J���c�zuww�7��g>�i�7�B!^c���x�������h��5�턐"��pA�0�Z2��u|�|�����:�vm��o�?,�whe�b���<�Xcv�ke��?��ڟ{�9����B��Z�E�L�<Y��>�l̟?_�^�_h4^�n�y�C�z��U��[�
��wU�{� K��jW���69ܞ����^w�p�Px�Շq���x�abfkBHy;!D�/�u񋂶F��T��ve��,ܮ/N�:���I�Ȑ��o^pJ�*���S�g�І���W_}UZ���Dmm-� -�\��(�����i�o�������k�;p7����/�h?��7��9��s���{�߽���駟��c�9F�D���ژo �h܋�U�������z⧾H%#�U�v�f$���V��,m�f�I낕��u/ϝ�'wՠ/�!�o�T�?�G��?�>00��o���=3f� !�B����mۆ��F[��1���j��Oq�ʠя����J���ۥP{.����XZ�0�;4���7��x�}�V���/K�����S����Ŀoq�nyW��ǭ�v����/nݿ[�]~}t���}������wn��)����#�<�G}�{�t3A�3t.��sxe�Kb.��|�6w�����BEA���n���K�����mۉ��&�U�g�;!e	$�jv=mt��Z��4ܮ����3��J�J�0���*�(��ҋx���b�On
X�8W1�W�<xPjk_�r%v�ܩ�_�[	��p�����Ŀq���n��倷S=�[���������bq7����\uu5z{{]�!@	�ެ��ߖ�;�C
�_x�8�裥m��rٷء�\��C�*D�R�k��3"[3�hqO��SXv�*����t+��u|�B��}��i�;Zp�Qx�s"�w�xH�>lh�B��)���:N���������ı��f^B!�D�ܻ�6���Ֆ������Z��	!Ea�� �c\+��=��v=��4�nnϥ��?����&����� ��B�v��F㍍�����-�Ο,qK���N�����n�	�~�n޿|�n����w����׻��>�m|���,]�_��q�H%Y���l��ʘ�=D���XMl�I�vQr����BEA����,(�����%�Ik�B���Z9��E�z.�ނ��+���%�b,B��	!*��&�!�ѝ)P�uY��n���)N)E*��9O+(���Lҭ���܉u���w�b�˩��q����{R���'�p-PJ!�����N��E�p��K��VD'�q/��>�n��.KG��wY��^_�V�Vs�*S���'���7�j"������ ���u鍃���o�]����ݻ����O}��v!�22����;7ڦ]vGEs{-�n'�8�ѓ�8&�/��*bc�=�f�˞�<����2�C=�{��Nzy�l�����,ϫV��o��Q#�-��7��[�L��Э�������oír&���Xܺ��ſy�f~v�o^~�s����wss��>���8餓p��J�wYK����e_/�ڕcv��Ny��u��D�=�#J>���mj�䰻�_6�0�B��n���}a���_���)�oc1!����'B{�o�QC�J��̈́)u�]_�Jl7��ە��l�
j/hF�BP��S�w/W��E���?��c�裏�A!$;�5tÆx뭷0m�4,^�Xju?�ä�N�Q��[,A��qN�V��XZ�)!PI[ �����Vy
B�9�D����"2�L/�P��ʢ	�+aF̉5b�̹X��!wBʍ�+#^?X%�|�U��xk[^[����'1i�DB!���{�b˖-�)��%���բ��vBH�Ҭ F�w`0�s(�H���ci�C=��)���>n�K-�ng����R�],���!��_��^���ӧ����1u�Ti{�~_.�s�n�ѩ�z>��3�
�_�hqG,]�%����_#�Ψ��,����k6��z�a�������~�;_d"����/�ab�F�5�n$NIc򔂚p�R�?z"U���B�L�����Eq�+�����'��چ[ZZ@!�>�k�0�o��6�u�]8묳p�E��c����)F岯ۡ�B�qC�R^%�䰻|;-`Ɂu�Vm�]&S�J�_B��o�5/doeP���!�q=��`�l��!�����=P��$`���BH|��n�\u�Q�K�B!v"�A�l�jk���ߏ��``��1��9g�hk@ ��s
��gx���{��b,m�ݨ���C����8'���W���b�
�K�dB)�.Y���sN>�d|�k_�g?�Yi[�~_.�k̮0|�=�\�C_�����м��ωE��5K.�X��aΩ�����A��	!�@k��/d,P�"U���`%�����b��0��RP-L�7/���d��8��0%��[�⩧��O<a�T��B������+W�s�����p�gH��v�Q�_H�]9�h冈�����!ټ ��}x8-^%�k"�л:�'XAլ _n���U�N\4o:V5�fEHY!��׷T!�c��§�mhlDGg'>u�񨪪!�B��tuu��M�l�1��xy"�B&��Do�^�B��Z�P�?��B�o(�ە�X����R�2��:���
�g�H$��_~�?�8�y��}	!�������O}J���ϖ�3K5���q���]W{���ͱ���/�z���!���ʠ�O�J�6��U�a{=CB��	�|1,�Bo�ެ�
Zm_P��+��f"�6�nl�N5���n�BS2� F1��Z�^}�U)`���S�"���o��&6l؀�K�b��Ÿ��P[[+m/DP*��\��fc^�����ar+���XFSʘG�p�|;�8Y��.\!C�R/}��p��xf�tP�"���ack%�)�>��&���v���8v�����B!�"L����uz_Η��p�`��vB������)]�m�DEEeN��LQ��]��R���!Z��B����u'�)�X�}�ϫV���C�0L!�8lڴIZ��n�/<���1~�xi[���BƼ�!�)沮��^��M�,����{�/�Τ�+���2f~V��H�����r,��U���;�<���̾��	)ap'd�R��_0�=m�����Ys{N��S�M+�c��B�2��70�nwB�rr/��f#!J=��صk!���x�&���I�Z�`.��L�2Eڞ���˾�KvWLѪPQ����Ou�]��'��A1�,65ԢR洃CC���J��o�.Xi���9y��O@Kx���bkG�Ըr¤!�t.��&�U��ۇ;�8T�?B!��KOO6�����n'M�!�k��V!�8ʌ�A�0� z��JcUh�J���?4���v�3>�5�gx�b��X��>�бl���ק���}�B�;��-�܂%K���3�ĥ�^�#�<R�Vo��1'��vx�Ny��!T���^H��b��p"쎄_9�	�y��k/m�=3������ϰ�_�4�u]�����!!�@D��W�t"�ѕnn7jp�&Pi�T���i�]n��(��v�8�Ǵ�� >9%`�y��c���X�l{�1�Q�H�"��.mmm���{���㬳��7���b�B�]����dv�B���x���*!@�1u�=��!v�d�d�]y>=�*-<i���6�w3���~SK�����?�D�^�44��R^l�@w4�/M�E�������x��������̙3A!���ScS�o�nkk��t��#�w��%<B��3)�#�{��B�F��ٌωu���d�]n�6�Q��p���P]�0Ҽ�|���\�����aThѯ�?��;$�� >��8�S�}'�p���KAw'�󚇘�zbL��^!�Q�P��:M�F��2�.�N�T0=��I�azh����[�������G���!z���"�2����h_�P�S:B��@��T��n�Bf{���v]q�`jA����
�{E��ul�Νx��ǥ?�p�BJ���~�\�O=��$\���O��ҶB���Ɗ!d�-Z�+b9�.�zj�,9�nu�A=�JtO�.T��:��<ON���h4�c�0f�,����!���� ��S�/O�Cm�� �x�x����b�1Ǡ��
�B!�m�[��]��z��뛫��!�8�	�C8|`��`�;4��9�7�˱�c������v�{�nc�q����b&Hh���q�FB�.�5���^5kp���c�8�����^�C��1����Ct"o�g�����z��XI�P���2�ҷ�o�K��u|�t94��ar������i��q_��ҁwBFGM���D��^�BrL+J
T�i����a��H���'�&���T��v�� ���� �����[��_���~�iD"B)M��/J��I'���.�H
�k��*�c^�����ldP"�Q�􃪰��\�E)`)+e���P2�:t�ԏ�D�R�+r��߈Sg���;r'�������:���^���hin�ܹsQWW'}>%�B�">kl����;̾���a^�W�����!�s�Tv5����|Ck3>����d�]Y��m�g��v�o���q�5&�w�Ԑd��\������x�������>K!�9�k��M��y�f�J�-��ŋ�2m��X���9y�Ӟ���ɞab�gy���e�p89�s,vGRK7���-��{���z��k:���j����}�8e��Bϐ����!#��MaR�}�T�B���L*�i�D*+�٧��8Ԯ�X����S�8}\>co�������_O��!��>�p��oH_��Wq�gJ� n���R����e�J-V�S�`�P��)��T�)*Aw���>aʗnf�*V%O�^�Tj��us�LC�-τo�7����jp��~�eO��P�uN���ߏc���ĉA!�"���ۇ?�ȑΈ��Aw�_�#�8�9��5mM	/0�V�ܳ��,{����nm7.Ʋ�ڮ�U�a�7�ԟ�ޡ2��-o�M��+~�<��ݍ'�x�<�����`;!��0�5���7�t�q�s�9��׿�ѣG%�^��Ӟ���i=Cm�]l�%���ɰ��Ǭ�]q6U�]Y����Ҟ���R�]�J�DPs���;O��3$�`����is��l�_پ���njOߖ��Z�*-T�C��"�f7�ZPG��
TJaJ�0��b�M^��l���{�n�:
S�R��Aw��p�����K/��+���jW�3�nv'֍�VP���b�[�5Aw����h�ܓ���zPޞ��K73����Ī��1(�Gښ���XY��C)+�}x�@5�	��I��ϐ��7c�[oa�ԩ8���PSSB!��\:::�`{gg�#������*�چB�$��aa����6�[����o(ƅfTh1��7T������=�S���>v�m����>���﵄Bʋ���q���htA�q��Iۜ��<�����5��P9��3���٢��.{���U3?�!��w�IԞar�h[͛�"�����x�	)s��!kSjo�
T��v=�J�r�ũ���B���^w�;�3�ƍ����kײ��BF�=࣏>¯�k�N"�p�B�ڢ�Aw���v㶈e�xc�F�Y�}+�úR�2"q?���5�,2%S�F�c��2���sM.}�{��n
V4U":Đ;!���C��SzQ��o|���8x� �O����<��� �B��A|�m���8p��#���Snn��֎
B��T�����֌
m�]��}�g+�>�cYmmW��V�C�Bz���c�q�1l_�b|�AǾ<F!�;����%K���c����7��ɓ'K����<������(y�g��q��(�cP�"��2ʠ{�3����B<C�7T������s'c��j�3$ī0�NH���/����m/B��a�"d>�`�H%R�����d&P�S����t*��R��<N˫��*	S������BF.MMM�����c�IA�s�=W2ќ�{I�*�����K:�.�Ti�JZK�R�r�	�ʟ|���ޒntW62 }��H%�M�S�U���	�K�K�� .�5���FO��Rn4��ԮZ|iJ�����Z���{�n)�>{�,���I��	!�R����c{}=����H�]3�Ԡ5~C!N3�ʏ�L�D��+nO��z�XٽCm�];볱g�-�n��g~�ȼ�]��Wnޡ���˗cٲehnn!���šC���O<!�b}����.m�b�]9榇X�u�ϗFlO�) ���Y�&��F�a��U�=�{S������ �тf�ó���� C�x:q��!A?�hN=m���4lm�2���4��`��@e���hzA���4)2��9n�On�Q�
�oذ��?֭[��C!�4پ};~������D+'�����cgh��9�����C��^P�v��Aw�p5��F���L��K	U>y0-bA����)D/��!�]�8{J/��G{/C�~����v� ��/~lcpp��سw/�Ν�Y�f!�e�
B!��җ�w����l���A�o�����+�b���~|aL3z�����:���w(���g}�c���skn���ڠ�@ֱ���R��u�|���\��=��n����ւB��E�E�D��q�%���/�)�n��h��Xщu+���3�%���>C�jʱ�H�w�3L��H=������g�pO�D�7�=ԅ3&ⵎ�h	;�B�wBʌ����A��--Pi�̦L�Sr��f�JG���g���� h廏ǭ]����?��;�B1cǎR����>*��?�|���K���}�Z�{���'�ԍ	�J=���F9设�3Z�t�Hn���r��@����RjX��p�<ak��p���!��p��js{%������}Sa�YD���?DCC���~�GH��	!�R�����)�YU���d�}(~Y�n{>� !��Yc�L�D�R>a�A�ݒw���YU��1��j�BM!V�w�?�`�{�N��<(��)t���B!J����t�R�}B�b]v�e�Aw;<�\Ε�>N�����ʞ�hlW�JQ��9�jʱ��X��7Ty�r�^3���3����@__Ż����Iϐ/��;!eĘJΚډpg�Z�ʳ�=%N)��	�Jhϯ�={�=S��~��NAȋ���)�}6oތ%K�`�����}I!�����K��<����
�y�������r�-�ʍ�|.��b����ˈ}���Sr�A�h���O��.߇/pGJ�ʼF�^/*N�neH�����I��cchvv�R~����Z���|b\���G"l����0��1{��esB!��"l��؈}��K�m�D\��~��"��R�Oa�o���b,y�F~az,fן���b,S�P�!3�T�ޡ[��w�\�Z[[�f�e˖I��B�"���`�ʕ�袋p��c���ڕcNy�^����!whf|V!��=CM9,� �<�fN?�g���f���o��3��(>U���3��!�0�NH�0�6�S&����G��]!V���n4��_h�G�Jl�Ƽ�]�%ʋW���zܶm�p�}���g�u�ՈBH����������K�v�Jp�%H�c^������%_�%G�hgPW��(�jdPݡ�g~�1[��Zp�E�T�]�x����/� R�G�*��z�L|D����d(���vk����}�
������A�K["'�D���q�@!�����&��8p��Ҏ������+���R�i�B���Oa���12��Y��c��l�ܮ�e�p1	��}�p�t+��iuV������l_[�b��ntvv�B�t���{�/H-^�W]uƌck��b�=E�B�ꂩL��'ƒ�v�c)=C#����ܳx�)��Z�]���#����Ĩ)��� ����RL��G@_�?մ`�ڞ5�����H��E(m�]+Z���:�V�R�ڭ
Tv
F^��&N��;v��C=$	T��B��>���J��?�y|�[��	'� m+� ee�|'�sc��+�� }$�-�FM�]���ވ�lrԁw_J"S�2h�Q�=��!ZE#�ۉ�)��� �m)Wv��8�s>9~ G������x�ۿ���;�f�����s�͂B!N"��&ާ��+"�WZ�x���lm'���f�pXo#|� B��v�+����`��l�Y����:AwA.ޡ�a�R�
������ᩧ������c�BH!:tH
�?���R1�%�\���*GC�ʱbz�v{���y���I�B�3�Y!�2H�lrO�z��r,�P��v������F1cp*������	q�	)q���o�{t���L�ʵ��,�.S0loO`��䤸eǺS�仏<v��A<��cR�]U�B�S���ذa���/��k�����q�)+�"0��X�v��c�@{b�ئ�����>ԭ�6w��Sb=)V)��uE+�f�J�J��&T�8������r%2�hs����1&��LT]]]x?�l۾3�O���F�!�B���L��с={�J��b�D)�;�k��ǝ!��j!��s�� �5����WhWs{�7L��[(Ʋ��5��x�Z�����R�#�^x�,]�MMM �B줹���r������&.\(]�8��c������g��G�Ɣ�r�]��Jݳa�3L]'����}��P�T�6��g8��'Ϛ�Ww�3$�Mp'��9����vb0K�٭TF�z���p{��y��^�����⒗,yLLu�����.Z�!�"ރ֮]+���;�<��}ƌ�6�)+��+0��Éu;.�c�����p����ԃZ�Ji`-ɓ@ne�АR��6�'���@�'^!y��x��7Q�"d����;kp�aQ?~ �95���/hhl��ѣGcڴi�?_R'�B�s���c߾}سg��pQ�{ooo6W�w��턐�r�\?�3>�cYmnW{��cY�b�c���Xwc1��s�=�{������B!v�{�n�x�X�l���J�y�O�9��>v�ԋ����h�3�:�.��1�=Cy��_��ͼBs�0���|e�\<�T�/�B2a������B��!�����*k��Ԙq�L�2��:-�y
Tv�ӽ���1��#B^+W��ZD{;!����hŊx���)���
�;֒ؤ+d�BB�F�(��]/TВ�ݒG���XZ��1m���he��u��~�ޗʸ�����Oq��ٓ�U͡�9w.�k�`EH93����Q��� >3��k��b������m۶a�I�2e
&O�,}N'�BH�Y'��)��;������Nk%���~#������M�,�C�����;Tb��۵��c���~�_����sz������n�:��oÖ-[l'�RT>��#�p�R���W_�N8A�'����Ct�+ۺݡ����Ҙ}�a:ܮ�'�f���|FAw=�Pڧ�	��;��A)>T�)A�03$M��0�n&R�n�M:B�Yk�=�"\�	�	T�$Hy=�.�5k���;�����A!�xѸ'�V�^����
�-�<�W���i��m�PAKO�I�	)ޞlk�L���[m3L�U�kE��ӂ�<(�82�1*Ɣ�&�>�фs���
V��;�"~��W�)5CR���
��"^K67K�x7n�N��)����*B!�:���hniI��;;]	�E�}x��ۺ*�@!EE����uO��]'�n)�����F�X����>g������������w(<D�	!����o�--g�u���N�%�.��O1<E/e��[L�P�/LݿOn�J��~�ǩ���ޣb<�ڄ��ƪzB�'��p���Z����70��Զ/�E���JY�*��iqJ�	.Y�/��2�)B!���������˗���/�9眓�����v�}
	�[=g!��v݉лr��X��!Mz�L�R�G���׍��>�^��L�*�T����H[Ο7OR�"dDp�7��w�b��>=1��@q��"^S;::��>���'N��	��~��>!�22D[{;�Z[�`�����f[gH
���;!�n_\7�޶}R�]p�cYnn��+ƒ��,����@�ޮ�r���J�;��y�%�~{�}���C$!���}�Y)�r��[��&M�d��S���!�qL1֋Q���&Zܡ�p�Pymh6t�ZP�����,����a�m9˷S�'��0�NH	q����4J��(e RY�������)��*�(7�\�ٽ{7|�A),�FA!�x��%��������xu�5��㎓�e���c�1^Y/D಺�Xb1Y�Q62���Z�J�v��Ku���6ܮ����}�~�ί�˷#�;��@�B�5vW`w8�O����"�����yV,����_#�O��	�e��ц_�!�Bʕ��!tuu���M
�w�o�]�!Zڛ�Cx��=Q�ۄw����Ds���gh�ޮ;۳%�P��=�Y�Sޡ�oX�wX��u���屾�>�\�w�u���A!�x���<��#x�p饗��_�:jjj,���C�3��g���{�"؎<C��'� {��kH��)�к�.=��H����{pѼiX��B���a������ATjHNaJ+RY�ZP�����*U�ݧ�2o�f���d�8���H��M!���l�ڵx��7�x�b\y啘2e�'D+7֋�Ġ�&��#�+����S��<�,ZeG�ϐB�J,CCzb����=��m���ۢm;�p�l�dȝ�Ct�'�>��Qc��?n��Aw�P�5R4�E ^+G���;cǌ�رc1j�(B!�'�]Gg�l��pqfVɆ�����Jb���"n�;�����B,�`{^�a2��K1�a{��o(֡l��*��ipz��;��>��e�=��lojj!�R
������oǪU���o�w�#3@�b7;G�x�z���S�0���ɭ�x���I{��V�t�=��Y�T�]�˔ڟ�;�����.����!e	�B
�wBJ�S���K��CYE����S���օL�*o�J'�nE�*��� �A�h��Y���z+v��B!����<���R;�W��U)�^YY�x���rib�g���xZ��i	E�{2����Ҥ^ =q��(�S_��B��\{jϭZ��*��i���X��84O)?D�}kG���C~�Dk��)�d����Q�0j�h�gm|?�@!�xd���AOw����� �F������Q�C�	!���-�A��`�7̘�9��ڬϙ�a K1�ٌ��|��v�L�ʱ�;,�w(ظq�ܼy��q�B����_���җ����j|򓟔Ƴy}V�)$�nt�z�V�5���3�}}�=C#�0��/��#M����<�wʵp�>,�7��+r'�ap'��|Y��5"J��h`�>�`����˜V�	��+��ħBαm�6����k��Fq�BHY!f#���;�������SO��R])6/d[/�(e�ob,&	S��	�J�"��)e�J�bג:���U�X��*�J�|��a�V��zp79˷3�B�Hc`ȇ�����uc�8f\�Ao4Ɋp�XZ��T�"�.�⭮�BUu���Z��/r�����BH��W�Ed���ߏ޾>�ŗ��O�.�{������a���vB����sD��9~M_a:복p��w���V�enW��3��)��ɰ���|�)�8p ��s�/_��/�B!���[oI_�:묳p�5�uh�=E7B�����������J0�������ˬҧ�~�����X�X�AoX��%��aΜ@��	��~k{���jZA�Ԃ�)��
i_(u��Iqˎ�B�S�>�����?�)�K�BH9"������ӟ���~:���:̙3�v��.��f7C�`�)���u�p|!R�53���LO=�^���
V��2���[��yӰ�! �q����ht���Ǘi��8�L�����&�(�Yg������!������Pb�o�|�VW.�>�Jߠ�UH���a�B�A(�Å�{�h�hm�m�gec�v�g�R,+3>붶k
�|I�F�Z����Q����������$!�Rz�Ϧ+V������*\r�%	�3�h7=E'C�vy��mNz���H{�iIZ|>�b�\��d��g_:]4wV4V!ʐ;!���;!�̹~)ܞ���ۍ2�4�Z�xzA�p{	
TnNn	Z�iᩧ�½�ދ�;w�B)���X�n���
\v�e����Ip�Ǌݼ�m��M�u���)��آ�R�:�9Zt��P����C�]�ʅ޶}��n�7�8� !#�7���UC8z\3k㟉K�5A|V�h�%�B��}~l;T�]���g�	!�A����EOgk�3�!ܮnn�ll������b�5��9ﰜ��Ny�bٰan��6|�� �Bʙ��6�|��x���?��ϫ
�����}��;�^�л]��2�;i�0�ص� �(�p{.�3	+�r'�	p'ă�57��ܱCՠf$R�O/�hoW�TÀ{b���<*P���U�9��}�����͛Q%���/n V4:������s��_��_YY������n���wYXw7����/�[���7p�o^���^��뭛�]6Դ�߅�������o�s�Q�V�C�V��d3C1E)���z�	�im�r=�\z��*��0�}P��>���}XĐ;!$Ns ��Q�a��(�����n�%�BF��}gO��B�@!^�*,�ٍ���W�-��^��p7�吻�Y����*��"C�)�8ҽCyl׮]��?��g�y�_x&�2b�"?��}��v~��`֬Y���͎qc�X�w�=C���Xz���oh�/Ly��s��c��;e�w���#&bծ�3$�Np'�c�3ϏXkSFS��p��@�
��M-�k�B�;xU9	Rv	Z������;���)��O����ߐ�o��n>w��C��u��uĭ�����_{ܺ7����/�/F�߼�Ϳy�z+���{(n�׈�{����o~��Y�����1{��4/����(�z�E�l�I�#�|�F��ɠ�I���he% ���D�R�d�B�D�}�~�BZ&Ta�بx�wB!�x������� �wW`_O�m��R�c��C���0�s�k�Y���C�Y�M}C���^�{q�h���~�����?����ɭ� ���M�߆����ߞ��!����n޿���w��s��r1���.^o�,gr�o^~�+h*#�o���v���R���K/�%�\�����>�c�Z/ďtr_'<C�|��Mg�2���*����Ý��`���Uː;!6;!�̹�ڶ��@����&P��N-��Yim/o�ʫb�v],"���?�	{��Um�
��"�(�틍���p7\:���.~�n�]��w'�n���Y�y��@��ߝ�_�p�k������n����_ĺu�p����+�,X��[�r2_Q�l[�x���&!b�CFm�z(�7�
V�F ��X4�A���! =~B������JL�ƬQQ�3�J?�(%�B�"���}~���t(��a�f\$�+����gd���b�Bʦ��r,#�0[1VF�]tOl�¸K���-�ϫ^�޺��r�-ضm��.�������pص��߭��Þ�Hn������^�(rӻs빋�b����^��x�q+���߼��+�d�#�o>��x\����SO�G?����/J��}f�pb�EY����5�2�|=�Kم�պ���y�;�p��V�EĽ�B�
�	�g�"�ј��	����f�
Zi`�/ 2��S��g��xY�r;�n����؈[o�����kafB!�"�%K��oHm�����Ri^Ю"p�)J�G�-1&72H[��]ĺ��KL9�mf��(e.,)�W�c��'r_|�,���	!*D���? -ۀi5��UŌ�AT���Bq�����A��	aO8��!^�BJ�P���z���+C����À{��Xf�v�w�Y��_)�ם�<�;�C
�U�B!�x���z)�~����.?���B��X)x�V�U���>����%�Վ���X�T�(�n)�	� ��	"d1�n��@��,O-�g���*;�b�O��ŷ}�-[�;���� �B�5�lق뮻N����ZL�<�s��u����d�*-ɂUb�4�`r�Rm3�פ�!��Q61Jo�\X7��ݙf��}��/u"X'��3�rSj�0�:��5����wB!�z���ā� ��F�j'��"�~�lno-0ܮ�j��j1����澡y!V�ޡS^9z���z�����_����fB!��G�X�B*����q�EI�>�������d >�3To��Z�3�B��̛�=r�&������X����R��2'DeW������A�)e!J��M+������/RNPv���書�����B!�#�V�=U43,X�@%�h�y�\������ے{@V���É��m��h��`%o7�ޏ����m/9˷��AI�W�����l�@e �)ՃR�}R� �V��B!��	�����d�]�BH���p�~��[S!�\���`��+�#,c����7t+�N�P=������o�믿B!�X�������W^yE���c�)(�.�y�#�z�Av�mj�0� K`���8��+T��S�d�m_V]4g�7U1�NH0�N���:;�����p{�Ԃ*aJ)Z��T���X�B)Rv�O������׿�U
�`!�B
c�����o~#�V?��1{�lǛr]��(e�o>���<�_B�J�++�E��`�Ijj�*X�#"����Z�\0oVՃB,30��Ξ��*�1L�a��R=�	�C�c �BF:�+`~���P{k���ka���@���EnoI�bn���cۭ��Fޡ/��;���z���p8���_Z���@!���X�n�}�]\z���w�����C�'<A�z!�3�nt;<Ch�ܕ����7L\������ʽ�6�h��9S���C1ݽ!Y`����Ҭ �5"h$PY
��/�n7�Z�����N^�
Y���o��w�!�B�e͚5ذa���*\q��u�SM��{5�^�6��2������lj�$X�MTc�w�e?X�x�Ѷ�8�l<ɐ;!$O"�>��V,25��Tc\��WI-�����8!���oȏ�:#tE�#b�?�b�Bʏt��9=�M��Pr�g3��,��=BS�P�g�`��v1�����:��~�z�t�Mhll!�B
�����s�4#�(�:餓��|���1;����b{�v��9y�����=&�A��3�e���a��=���h�T��>��3��	q�/�aTw�$*�M�zU����������1]a�R���������tHK�,�c�=B!�8�h;3����O�Su�Q7-�^jM�nK��=��_�`���`��~�k4hדc�Vr?O�3xJ���A_|	�@o 5&��C1��Q�/��z�vM�g�?���B����P"����3�O-�h�gԇ�0�_B��@�R.�BO�A�7�z��<��!�h��a���S��a�]�z+�^�av�zgg��c.[��3>B!�m�6)�~����Ø1c<S��]/f��u��3@a��*u�(�Q���h­�pѼi���Rd>7=������4�R��n�ҋ�4ܮ]��)Sz�}�X���X^z�%�r�-ػw/!��<������·��m�����/Gee��"�v�Q��<�l3���	r���Ա|ꛚ�1��PmQ�i݁����S�4	!�0����V[#��*@����z�c�m��g����U�B
g0��4�4k#C�1Ѹ>0_��?�K��uB��I��C��K��k�Ê��!��7�l7���0ܮ��Y`�y�,5�P�ꫯ��#g|&�BF|���G�|���G�җ���KY���^/V��}�0a��y��� m�y��g��:���/�7˶@���OOab_#�`fk�B�2�����J?�S������R�������m�݆g�}�4XE!�gm���_�6w!Z͟?_��	�)ۺ�T�籲My��`S��a&V��V��i~F�v�̹s�\�!��}���sB!�B��n���&�a�����XJѺo�_�%p��+��S�b�g��Z�
�B)MMM��O~��~�����1~���ci��#���~�P��{�1��sG��!//���Z�bѼX^�iW	�
��OLaZt�xMR�@��n0�H�K�=-V��� UB�v/
TN�SbY�z5n��V477�B!�"Z�����K/�D���*GE'���b�RV�ɂUz�A�
�6���,d�~a����۱�F�2���!�B!�B��º�nW5�+�C�ٞs�g܍��f�a"�.}�������_|�E�;ܳg!�R|D��#�<��k��?�!�8�U�*0�z1��J�3�b|Xnp�x�>��Ɏ/�Vk瑯��G*�Be9V�n\0���g�)!V`���"P7>����Č(���)u��3E�@���Xe%ܞ
�g��<��	*ۺhmS
�Y�&34E!������=�܃w�}?���t��ˡ�!����n�Jy_Z�Y�J��vYf(X�o�����s�~C�B!�B�H��y��q��Vh�B�vP^�%ܮ_���!ʺ���v��@��׳����`�ҥx���B!`�޽��/���>�_=&N��I��ʹJ�3��"��T=�P���5���ؖ��=fҊe��,�_�uέ;O7𚎐l0�N��L�ǿU��`t8����^�H�R�ۃ9���1��v�He%��T���*;�|����?��o����B��ٴi���.�/��r隭�����l�[��1����u��^�)��{$�	}M���s���(!�B!�229k���M�R,=�Ь +�p��;4���v��(o(�C��� �~��ޡ@���b��B!�A�W�^���~����NS]#y�#�;��x�����ɞa�i]�"�3����s,��=�0N�}'N;b.^��b,B�`���P�ǉc�1��)����@f�=hw��0����/Rv�Y�zGG��<��� �B�������ߎ�����?�9���<��`��U��N+���1�s?1�O�Q`���O��[(XB!�B!#�/���ѐlOy���(�L۝	��c	2�C��K!�n����)y����B!�E���p����O~�1c�x�#�zl����l�v?�v�3��Vy�:!w��1�M��Ġ�3�~t6��Yuxu=CB�`���]�ǩ���ۯj`40�/�-��@rQ�18n�n�G_~�v��ٍ�mذ����� B!������ޒ�ܯ��:,^�X�heE�Ү{A�2ڷ�m�VYZ��*kX���%�J!ZE"�߅����N��B!�B)|nz�5"Taɞa��K��S�	?0�G1V��v��(�ǯs��J���!!�R���U�V������~�3�x�Ҹ��v���� ��y���@zfA��+����ZL��tn��%�.���i�N��{9�3!z0�N�T���Ξډ��1�`R�2�V0cIݝ�'�ţ�n�C\*'�*�c��0��n�w�}!�BJѦ��?�7n�~�L�:�VQ��w�ڭ��H�R��c�[�@yU�j��R?����H�W������w�!wB!�B!��9~J����t��v�0q;��ݩp�<^.�v/{�����^�u�]x��08H݈B)5�����W^y%��?�555յ�������m�z4�&<�t�=f0�]!w5�׃�XƸt�Dpxd�;�l9Ȑ;!Zp'�fB������쒚��۳TF!��U�p�|�PH��\*;)���-[����MB!���<�6oތ믿��~��*�I�^��U� {�����{��V=25����t��t���M�} k�&�%<B!�B!��'GO
b��.�|~�`���=�GLy�����z�a>�v�~��v�ns�X�uz��BHy �����c�����/~��;.o�P�^�л�����Tz�Z�Pr���Y�f׊�q�pnl�&�BC+C�(a��	��=/�ۏp{k�(�jo׈U����L�=d/�p{�)+��YѺ�d�����B!�������_�_|1����a��ўlb�����ؔ��!X�"���K�,��|n����-����)ڱz�0���#�B!�BHi2�� >�߃��Xf)����u}À�?�y��k~���a4�#�<�;�}}} �BHy�u�V\{�������/�\��s�#�;֋���6������ܕ�+0��2Wl>à{bc�0r?.�c�cOg�!D�wBl�º(z�&��m�!��v�@�h�t�=!J��KZ��/ܮ�Z��p{1D'�)��޽{�����úu�L�O�B)m�P�裏J�K7�p�=�Xך���`W ފ`U�ԃZ�.ٲ�2ȏ5��1����c�=�8oj+��B�z!�B!�R6L�ǿW��`tȴ��7�C�e��_��v'|�R���;w�č7ވ��z�B)?z{{q��cӦM�����ӧ�j���sٷ�<C�}M�r�=���	�+=@Ց
�0�3Ln�D�8a�r�gBdp'�&.��(iۋPEe�H���Su�=�6��?��n��+gE��"Pɷ_y��z�hjj!�BF|����i��ˤk;7��s�׭m^�r")\	V�XJ�J$Ī���CX8;�e�U�K�B!�B!��W�ǉcZ0�Q5��b�����@@�˟Q�e9ܮ�GZ���av��^xA*���� !�B�����k�a۶m�����|Eu���G�]�gh�g����)� 2������}5������	�x��?"��;!6��#��5!2hn�,�&��ͦT�T��S��m_�m̥K����CUU!�2��
�/�}�ᇒhu��{��!��d�Vʂ���k:�} e+��`e(Z%�*e+CO�A\0o�o�1|O!�B!���S��+S:��ݗ�+4�Xf��z,�����b,˾�N�]��nw��#�n���Ӄ;��V�B8!�BFį~�+�������kQ[[k�G�]��gh��U�0>(y�6c�/��_,�1L?~��D�g�����X�{4g&#�	)��N��P#�������4��$R�X��kU>b�����V���!�BF.����G}$M?x�I'���`��U�UM��wu�ݬCA��p{j9�����ƹus�t�$�B!�BJ��χf�!�ѥjnW.b��7(�c��n/�?0�p�֭Rk���Q��!�2�~Ճ>�M�6�n��������J��ݾ��g����
�����[1�2,e�=�����pW'Q��*��>2Ra����?9����T�Qs��􂁌����`6�`��ۋ-P9-H)o�RѺ�?�	��� �B�ڵ?��q�%������4��ӢT.�C�2z�vVv��3�\���к�p%?GE�=��mo��Ś�!B!�B!��X8o=�͉p�N)������>���J��K�`1��B�z�'p�M7���B!җޮ��\w�u��׿��t���	�d7�f��v��)=CO��r7�˖��9�y���ә��� ����z��ȅwB�dƸ ���Ɛ�o:���(�����go`�;ܮ�(�v�����-�c�����?�O>�$!�B����'�����_��f�rE�2ڷ�m�llp"�n$,%��n%��J�2���E)^�~��*�Ww�������}QB!�B!�48�}�{PQQ�[�U�e�g��{�4����#�nw𽥥��z+�z�)B!�����J_~۲e~�ӟb	���v�Av��x�3T�+�%���B��f��,�/Ly������8�nVs�g2Ba���<8�ڏ��6c``H��]!PemoO�SE��U�����^�r�WL'����~�!!�B�X�n���j)�~�i��E�b��!w-�s
����6�~���T��ah^t�i�*D"�݁����e�B!�B�6_��P[#B�
��v�G����,��r�;���+��o��&n��F�޽�B!z<��3���ǯ~�+|�S�*�g脟�g�\�#�n��kו	��jhm�]{\�_��1��g���]��ȃwBr�*�Ws�����%�t*K��z!����Y��R����*�"C4��oVvww�B!�
��Iܿ��o��k���/K!Ȟ�6χ��q�t�=��{RtҊU�N�5�rQ����#���š�S�����B!�B�W��� �:��bU�x��Y�����Y1VΥX�۶�ʱCCCx�Gp�m�a`` �B!f������}|����e�]��{��f�uz���,���u3`��]}ݧ�eQ�<"������!�~��}\�	�O����r'#�	Ɂ�/����<��FPO��k`HTV���{6���v
T��zzz��=�P�vBH�"^c���v�z-> CA����GͨZi���ae~�AFq�x�H���h���G�]��{/�mۆn�ӧO/�(et�B��-X�r����Ě�n�ߖjE+�k<�K?�X3=�B�����{Éc[���$t��B!�B!���	AL�	_0`\���;�bɋ�g����c����ۋ����oGG�T��z�jB!�X����ӟ��Ѐ���7n\^�v�˞��s�_^!�gV��L���tP=��R�d�5~��F�YC��3~�r'#�	Ɂ����ڒnW�܍��u�uE*���I{�R�A��bTV���Ԅ���wظq#!��xݭ��AeUe|��^�+*+��V�ە����4���� B����_�gE�D�����'9,��M۶c��G*5�+_W����2�����M4I��F㷓�`��il@�9�9Ab���!��o���}�{R���'��(��y��=�b����ۭ�U�ǣZ��R������l�F�����W���=��^E!�B!�x���8�b/�P{���vc�PY�����e�0�R�R�;��3��e������ZX	!凔�P̰!f���X��t��\�3���@3jg�w0*�@�L��4kphC��%~[�
�c���I�9b�eBʋU�V��?����㎳��e_;<C��s�wt:�nt�1��b����)g���U>�|��qi�Qc�[�~����0���ȀwB,r�<?z[vJ�G�p{����:��n��2��:�
�C���^x�������B�7a��j��֢�v������&L�~VƷUUWI�fdF��r��xL`��	����"�p{�>~K�S�:�Gs�����c�QuR轿��}}菠��}�۽�=���	K?	!�k�.\����kp�WH׊^�̶�-X���+䞥�A{=�K݂�҂�,N��*�sd܇R�J��ub��*<�!�B!�B��j?Nӌ���~1��K�g�W���٬ˬ�����l��W,˗/��7�,��B��xm�Q��,Œ���vQ��L���m��6_vlo�G��nD�]�`� ��s0����0+"|¾~�,K�?E"�m�	�6"����@�,X�q�V
��ٶR�[E}�S�?R�v3�0t��(^�O�Њg����8)p'�'�b��!-P�U�Z���T�`ZA����z�
&�%��X%�eQ�����s�=X�t���hBH����ѣ1f�Ԍ!�T�֢������ޝmm��ݎ�8�8s.�����:���`�O��=c��q�`{F>�����3��}��Ĩ�@uu��(w�)���8F_o���{z��FO8�t���>��L�Z3:-��%[�lI�|sB�$�����'Ɇc @��l`CH�$˙d�KHv��`ccl�C�-[�uߧ�?�=�]]]=�#�)�ߏ��S]]]����zߧ��BgG�QM�ID|`A�Gy�\17������ډ�@=Ҳd�b�kZ��*־��0��f��^�?1Xe	�u����
7��{�⼅���n�AAAD*��Θ݉ޮ>�Q����)V�)t�,nW��r1_8�����Ʋ���?�0�{�9�z�h�M����'`x`Eӧcڌ�F��B ������Y�	�75cn�<�lp���^�Q��'�E�9ϴA����Nlذ�!���P��Q�0�<��^���]���E���w�%��g�0��Ӄs�s�B]Fu�:� &$p'�(,-���Y*���W)pe���
FPq�1 %���a�^&��
J%3� USS�q���o� ����/S�OCaQah*��:u�1��v�gYu�'ڳ��܉Y���򱺶k�B����]�D��O*W�Tu�n��v�Ƶ�jY(*��T:{�n�8�í�9�ww���ۘ�ԝm��n_�}�+�����z�_�˖-�{�IU7��7&��OGu��=����Y�*�# �@��Víu8���5�� � � � ��������{��#Mf�0�0�
:\�#���<��+���s����&2��k�.�u�]غu+�H�z:E�#M-
�M1{�����MF�q"���s�g�TL������=l����'�:2L�j�H4�~���Ǟ={p�m����*�B�X��Ĝ��>Rΐ����!�tqgm�?C,�0���?{�y��|!��;Z���xi	܉�	�	"�Xlݔgy�<��r�*�pmz8/d�w� �,nw�08���hq{�T~�W[�l�w��]�߿SB��L%��>�N�j�3#�1��m����x��|�#�'��������y���yv]E�#���hi5&��J�� ����'�vĀ���v�~���툡}�q.u�e�mس�Cu��]�]����YZ�M�fL��0�-6�!sy�7��P���)�"��y��˶/���Lض��+U��T�֤�z��}oll�5�\cA�v�ZG�$��D,K�z��܍��A����Z���;X%׳�S�IX��b��jlmAAAA����-�F,��a�#?�qo�M��s{,�X���&`)��1V����)?�'w��?��0�jkkA�]ۘ}���(�65,d��E"9�� v�٤b���0�b�wf���م���Щ�S�DeӦM���G�|��8�Ӓ*d�2��X�%K�I�B�џչ�pNWN�/�G�m�����?���^����-1q!�;Ax��v�Z܆���q/�Reyܹ�=zpJ��Bv98E���.c�o�[�������x�G�����|�L�ʾC��w��f�&�M�Z��=UwC웛���3�iƌ�z���Q�k
Zp�]$�vsŎ�6#xR\Z�lג�;�o��ڝ�P�d��<�v�cWu��B����5��]��"a#v��,s���\vp���cdt��������n��H��R��g�<������d�lh�T>\����[F"���y��nP_��׌{��:1�gY&�"����J�����>��k;28�9�U�9Ȧ�!��>����n
XAAAD���� F[����>�"v����y�9COs,1o����Oq{"���<��>��Sx��ǍXR&c��S*H�)X*Mr�w��G�� '���5�4�2��S,�Qn�#&�#̭�Ә�
s"���0ͶR@g{�v�Iɶٵ���C��	�Fax��9�s�X����=n��L`fY��YOf3��Il�8��,�|�wફ�W^i�W��3�3��,�����I�.�
�����v{9��y���G���k�a�7�^��ʫ�N#��ALLH�N
؏��UC�m�����s�-r�;��r�N��385���P1�࣏>�'�|2%hD���U�%31-,dg���mX�x����%]|c^�t������vE�B�csm�.�R}�I�\�v��_0�7 �ӽ���>y��]��ڎ��Z����o {���t�4��Gttvt������>l������x�	c$�o�%%%)sb�� >�+"wi���o�%|�F�'4����r=�r�����������L��ȝ � � � ��� ��j�)?�0�r�y�0`Or�19�;F|����D�c]��Յ�������;L�Y;������"��`�4��G�K)=���PR63fcFq1��^�%�=t�	�S�PP��3�W-�Iɶ���q��s+�d��u(�7���bn��mm�H�̬�e%�+��y~O0�̙2a��z��� uuu���PTT4n����D���5-��?[b��D��ײ�z,�Y�ݭ�3�#�DAw�PpA�������؜��Ђ^�Fs`�<�S���� U��R��Ǻ�СC���	�P���o�Kf�����Be��{��'���jk��bjM]�ol��k�[d��k�bM/q{�]�5��:�-/�^�i���E�\��ܖ] ��2�G�T��*{�^跌��W�T[�����r��-�hi>�CM�)u '�t��#��ۇ���cٲe	��uY:����͠�5����D�r�E����wk>��n��9��So�������]�AAAAĉ�),6bd8�!f��7t;��e����۳�|����#��eR�L��`�e������;�i�&�`v3f�4�졉�
��P�{o�D�D�a�SS�O3���F��vwv�����	ߓ1"4Ad2����iܛ���(g8�u8E��?�W.r��Et��F��2K�6��4���!��9Mh/���>2�"&$p'��0�R�����:�G^P�`��󲸝�s2Yܞ��۷cÆ���A�	�3��Y������9��Zᠹ��{�\۝�jaA����Ĺ�;�����]۝�v�k�)$�kٕ����+�O܎���k���hn�r.��hj�1-XXc������͇��Ԍ��0�Bg�H'���7���r�-8�3"o�rT��,�V��y��~��Z�^�#�<��W�JX�2+��T!z�����C�=��tM>^�Mw� � � �HyAങm���4ƒ��y(�۝BvQ��-j��S,����[�kN/��n����o��;���� �MaQ��C���3Jf:�������UF�3���C�����H"R���lٲ_��׌�ᩧ����a�e)g���M�s-	����,��T��l�9C!�444�O���o�O�=DL H�Nk��۱���w2�T�۽��5����I�nϧ>�����xTlH�{��b� &3�:�Q%����M�"�`܀K�񤺶Q�]��{��r���%nWu�[^���M�i���������暳̽��ޫ�]&���u<�]-++Ms�b�Y���M��`�7���ALV:::�`ss���+�{�x�=`e<X�kµ���Q$G��y���]8f�pq�Ԧ#���C�`��-�pFu5^�K�^AAAD<a���W����!nF��b�@��m��@0�1V &S,�9�w���3!?mi�������}� 3�X\Z��ٳ03�ʜڳs�A�B�s����a�nAkhb�A�W� �C������W_�/|����3��,�y�t���푞�Q�a��W��K��ς9/׭bĜ!o�O���:qAe>��C���ā��bZ �G��H�%��]5A������r�eׅ�C
�Yܞ� ��?��{��"&%,�T:{6J�f[�(M!�v~�Q�Rܮ��we�jܵ��\ۙ[w�I��n5/��p�R��C�c�O�vCt.��vy;^�|Yܮ��Q9����\�y��]�pIhZ�ب��ى��8x� �����L��9~�a4���k�����IX1����K��]��DsdP�sF
XY'ɕ������X���ű�5�{#Y2AAAD����im�tn�:�s�����3�&pW�b�yC�cw�p"���������������1�	f���-S�ٳȝ�H:�ww��9��`����:�d8�3�;��d���=���ߏo�����O��a�6Ɠ[L���|�ոG<F8�Μ!ˢM�����y+��� �		�	"DaN�+:���Q��#�T�<H%����/A*y�A!h%��?n��v��.n����<�_��W ���f�a��}��2)�)�زf;�k�umR�,h�צ񺶻���������e�T@�ڮ��?��:s�8�ݧ�Eum��O�v�k�k���'vV�<�N���ӧc��%FQOw7��1�{K�!�d�����׿���q��c�ܹ�@��%ӱ!=D�Z���{l��]���|����M;`�Kx����01w6��ˇ��2����&AAAA��ӫ�l݃��W�З�]toL����Y�ܡ������a��!q{�m455a���x��A�v�*-��Yef�pz�G� ����r�lZS����f�55�dlHL6�}�Y�fݺu(--�؜��z�[_���u�6	���f����eR��Fݱ��i���X���"�!�;1�aOX���Co[�Z�*FR�������T��ݿ��ʅ��w7�4e��
DeJ𪹹w�y'��׿� &:�S�P~��tV)��k�
YܮKK�VU�v�[!G�\���Q��a��mJ�E�ф�*!���<�i7��.��Usbvmw��%<�[�ԩXĦeK��{[��1��Cc�~]�u��J���z�~��[oŲe���m�o�x�#��ݸJ�j��*X���z7wY�΍�y�	�@U��d,���!�ݖ�����AAAA��e�A�u�"̎*n�ruX�vٹ=K�ǖ7�l�%���q��"n�G��߱c�!���AL�u���g�)S�bDf��Y6J9���\n9��߈�����C�BbR��k����ظq#�,Y��9C���>{k��%�U|�g�?�3��(n��C3����6��ۆ�-?Ӵ޽X4sv����DfCwb�s~����C��풘ݽ,,l8�ݢ�,O�����\��LM$q{�쑖�ڵ���W�����C��T/Y�9��hjQ�ڈ�k��[X�,�v��.��Hb�q��]�V��M���8\�M!�%׷�E=�]�8��;�������bgE�sAگpG�,s��1��N<h>xuu�ݽ�� ��FCC�����[n��g�9�U�e�,r���D�R��92DO��nl�2^��Bw��*���M���8g^>���3G� � � ����)YX܏=�S�)���{�3��g�6�r	�yC���63!q{�˘(lÆhooALd
�LAY�C�ΦS,��TD�����tک8�Ԅ�����1Qٽ{7���:�p����>��9C��'r�Ж[����q�Q���P��l-�r����:�{c�X�} �eh�;��TH�NLjN��P�oq{80)Pe��;�����p_P�0�^��@9P�Qd���,{��׍�)@EL4rrs1{n���bny��TzE͂��Esmw
�!�U����xK��Z;�k;�`��O�./����-�wtS�,�v�~�H�k�(&W�_���ݵ]�ɵ�т���x���4E_���<TU/M�8��G[�a4�գv�^���� &
�����{��e�]f�c2��#QcY'^"w�9�M��V�ۓ�ً9��)n��y�*<���ۋ4��ƹ5��nAAA١?�O�Չ��G�0E�.`��Àe�������b���y���2"��)'���`�z,���s��_��_08H)�ă��O�6'-[b�~	b2�����U������4��lj=�QgC�HGG�!r��w��K.�ĥ1�w��O��K���s�G6���{k��?ԅ�!,)�����l��3fwㅺ��1�������,�D�@=4/a{�@U �`��K���[�.�g�F�Jp\��VV�څ!Q���(n� 1Q�RT�y��7>���R��[M�\�5$͵])$��!nK�����'�N��brm���
��p8�z���>j�5��?��]ؚR����cum�����\:{�1{��ho���z��p7�6� 2���a<�����;Z���%T��Ht i,������k���<�U���)Xe��%G�p�<������j��G����h�A� � � ��˧�G���a�ۃ1��Y~P�Ypo�k�%���ڕ�X^#?G��SN0��,_��� �<�b"���U6s�S~A>�v�!q;A��:}�1-Y������C���݇��A�3������~|�[�2�s���F����c��?{߿"l�%�c����?u�0�н����)�Kd�Ed($p'&%E�YX3�	Cp�ڃ�80X�����`���^�A��9V�omtq��d�G�ǞN{����SO� 2�¢B#5��ųJ�r[��丶C!n]��]˔}�uy��?V���b|
ۍ?_����G ���~Im� �0.�v�X�k��,�k���横�u�;����j��>i�:�eF�cZu����`_]v�܅�#��D���kmm5ݧO����X���^�ږ-r_����=9X���,h���#ݟ�e�m=h��EΡc�JP9���$r'� � � �h|rA�-���*a{4q{0 ��v>Q�3s�ޣ?˂v�(K�b��+n��l�v?����ꫯ� &y�y�;�a�U2{�k�I� �0w����tdt���ذ����& �_KKn��1�#-�$���XE��,nמ7���/�e�%���=gȄ��������QD�Awb����]ރގ�1�����T�H���,�}AZ��ۅ!ҏo�瓵~2����O&����Ad*�)r�bC�M��Xf
xn�.|����н��pmR��.��ua�HZ.w��!��ro'v�P�]}<��L�k���p=ͪ���Q������%�:ˋta=sU�Q��Wy�uW?U뱾O)���+W����kOcC�|��{k1:J��ǟ��'477���FEEEF�)r�X%���Э�2V��TA+�����n���&v�PY�����S|�e���c�4���]���AAAAx��,�����|a���XcS,o����yC��a���bv�}��.ng# �[�۶mAd2��3o�a�5{���8�
�V�ߧ��ߊ�v�������� �L��:�6`����3�:�j�6������϶���t��v|��ãAv�aiI5v��DfAwb�q�B=--�����Ә���<wY�)@�r_�DA�Ӆ��8���Bܞ� �I[�~=6m���4���	�+��[��Z�'��v��]%��E��>�;�h��p��.�)�s;��Ph\��*�v���X�ǵݽY��{?uE���mW�4Kq�I����5��4g=(]��m��fwGjk��ݵ_�J��>��jj�v?}���E͢E�480���Z|�m���N�K�]s�5��}ɒ%��g�Q~�%#x�G�.���e汓]ܳ�C�����*��'/�Z�T��}���*�ŋ�S0��]'� � � ����� *�F	�an�	�CY��*W��f��M��X��!뵙/t����D2A�>��`�z,fv��"w��D�b^U���>��A��;sV�1�>��nAc�>��v���� 2�͛7�;����.,]�4�9C?m���]Ŀ�=��0���ʣ?k�|a�џ�W�9V�������j#�����X�݈�eh�;��H�NL*>Z���ûMq{����)@�}A��n�?�p�h�vU��{��;w�4>{����-���A)��la�7��ڮ�%nwmZ�����M�D��C!�v���%$W���Mu���]d�]�U����bn�wm/ѥ2�E���͸����4���|]��b��T��#�]l+7?K�/3���>���aǖmhnjAd�~���&6n܈�N:)��u���-r�
j�E��u����B���)�ٞW��ay�J��6|M�UO{έ)�ov� � � � �� pjq�z�=s�^��\��;4��bsn��s��2u�0��t��*����q�w���ĉDf��UL�^Y����<�onI�{Ǧ�����6c�}���QAd
,gx��Wǜ3d��`},��K�.�����o�?[�>k�Gfx��l9�C0Â�<!�
���ϟ�Յ
1Bw"C �;1iX83�i�{�%�������C@p_���GT���C2b	R�%($����X�mݺ��r�m�HxP�9�3���h�)��\�3�\ە��Q��x��C�'[�m�K�k�K��,�v�$��C�����n.-(���+VS{{;�|�;�mGWg'"�imm���_o��]�6�n~�e��ݹ=y��!9�_u��U��������v+`�R�S*j�AAAar~�0zۺ��v��ݕG�	�R�P=�stc�,���*�x�c%#�7���/����Z��ߏ��<D�îs����s�8rA��3���9�nj6���cxx���^�o���K|�l��d�/����{�g���U��6ms,����'�ź�\!�z��p~u>^� Ad$p'&�9Y8*�4Y J�<ە�(�Ђf`�����Q�`U�;0�zn�%m�{���-(�����Ђ �t�}�K�f��f�+*��L4��]����#\��+;�ʞ�v��
1��>;���>(���z���+8廉��&�jA�?�v�v�;��G껣�(_v>�y<� ����}0�������u.������]'Jߥ���˻z7��ǟt"�;��:���w`�@�Joo/֯_o<�q�e�������XJ�<{�;.s^E���M��W�";���(#@e;h��G�{�f�աrz%�;FAAAA���k���r 9��Qs�*��@8wP���X~M�����C4c�v��)��&Q9��l#��D���4�x�	<��#�<A�3�PV>�q{ @"4�HW�o�9e�4r��ۏ��z45��J��=������6r��A��3�I��ݙ/4J�yD�8������N��r����=���tD5���[������������Ĥ`mE?z��L���k�A1Xe/p/�Z0�
Hy��;�ܮ����|JEP��:�c��K/�� E�)�S���T��j��
F3�º�D��b]�Brg�\��^[%�p
�]�AW
�=��Z�v]�w�k;��O/q��OBr��v�L�hS)܆[����.��E��s�\���v}�V�&���/������2���vg����?q%��Q��z�a�Y����}����� ҍ���>�������m��fZ�*m�E�Z��Sts���5� "���*�"i�xpJ
PAz/���"`548����g&(^EAAALbV��{]#=��Jq��;:r������vA����ܡ��$k>�ǫ���z�!<�� �tf괩���6��|a� 2vO0A�1���������Bb�HGX���DSS���jCW��9����D�>g��X*���Q���P��jΛ���rS�.��8	&YY]�XZ� ;SҐHoH�NLx��d���	���� �/q{@b09@ɅAv\��VV����L�.�t	>����z~�ӟ��G��(�S����WV`��j̜Uj��S����n\�a�9�k���n��K�n����#�g�;wS��/C)��ݵ].��)���x���tm� ̏�w��;�k���¾)>����?_׹��O���Oe�5�����v�ל����U6�KJp��?�Ύ��`;>غ�== �t�g�A__n��c8�LX�m�$B�n��o��!W�JzPu�|u�2��O�X���Ἢix~7�� � � ��Ɍ�,,�:��`��J"�H�v{�g��=�1V$�v��nq��SHD�/Q��T��\I��>���7"������
TV/��Ad>��X�t	�Ο�C���{j���"�x����ڊu��aʔ)�y2F2\�Ǜ'�wn�k��̈́EJc,�G���q_�#?��23g�p�a�;/NG#=[�B���h̝��A݈H_(�MLhV�Ά־���AQ�.�\�)G�J�#/�e�|�����@�xF"��J�:��B6� ^� ҉¢B�*+��WA*�x�]��f<*q���) �����ׇ�k�R��
���߮F#��K�g���)X���FT��p	�!��"�ve]��]*�$lw��r��U�N!���x\�UsN%�Uյ¹#tTފ�37��ӵ]:?<��l_��A�i�g��SN��9	���a��7��;�V��W�BOOn��6et�*��r��YƯQ�u����C���#92�a��`�����Lv��.��ҝ�v����gTW�ս�0(AAA1���N?��=]C�e�>+r���k{0<�37�
�D�\��K%h]�Ŝ�#�0���d��Zv��a�_����@�Ƭ9eX�����!�۳1!�RX����}՚��߰u���pS3"����~gc�{�3f�4�7�u��E+r7s�,_h��f=��?��k!	ݝ�A�K*��/�?����}xn7�C�/$p'&,��C#��vPJ�<��f���v��rap
�Š<�qo�ma�q�_�1���u�S�������/� ����[1Ջ�pjz��q�?��nV�!��k�Y7��Nնk]U�L�_��J�,���r�NY�C®�vH墛�&W��ס�U]�{;Ϊ�|Wg����!��?wW=�a����sQ�����z�黠]�� <���Gw�qm�ͅ�	�+�0��2t=�m`��� A��W_}�8�����dt�*��,�m󺠇����<J�`��t�2��w���b��U,XfMB���w�bYi5�Ӱ�AAA�$��ݭ��	c}��d���s�����?�"l�h�%�Y��i2�����x�8p 7�|3�n�
�HX,oμr̫����� br�tGl�61�@��=�ݵC�� �t��^õ�^�{�eee���1���*�mE���l,���������򽬘/G~�-�r�QF���\���zkk���rq'��ÁaN7���� �jxA��/�T��])l�>��%hU� ��r�e�It�*Ձ�X�a����/��2"�L)*D��E���Fn^�Q���k��7����}�����Xׯ���:����06�vsYl���Ϳ�-�>��t�]�U�Nq�s\�U�w�p���q�k8ޮ��j�YO�w|����[y|�z��X쥭U=� ձ�%���*��w�S���vT}�M���?�{҉�W[���mAݞ� �T��o��o�ƍ1w�ܔ��E�!x��d���,|��$w-�������]�y��+8�%rwM�;��l6��,t��	� � � b�qlyC-{|�U9�@ `���GV��,c�5Ų̱��!���D��D2-��ZV[[��n�	�v�A�3fc������Bwg�i�AĤ���:�h�X�
�5b��8t�	�j6o�l��+++Ǖ��[/Y"w�D���2�u0�^.�zޝ3�.��{��{�-��<�V��s���A2�"�����#90��T�/$q{�����~�t���v��=U"�T�bY����peOD*)+��E˖a��2�rݧ`]7+������;છ@�vQ ,���b��sA��(�D�b}I��Aֱ
k�>~���T`k�������w;~��ȵ=r߅�9�>G��R�n�9�]�-U5ա�---x��M���mA��M�6��3VUUU)�'*x5^�
���(q.�.�n���Y�tqĠ�3@��9t��+)X580�O�����|+�FAAA��)����E��=j�P4�
�"vU�p���Ǳ���.��t��ر��744� RI0;��U�Y��fLA�����ü�
cjomÞ������#$4%R����q�5���{�ŢE�&��=тw�����}=wq�yC������_{�gu�P��a�)�/�G��`AZ��ɝH/H�NL8�/��P�n����y��tl��UkR�kxA�{����u�ReZ *��>�[o�o��6"�?6���\�b9�N���c� B��}��Q]�b��B��|sQ�Z���[��^sl��j�����;�:ŅΉsmw���G�;����]W�K�k�]�9��^:��}u�߬6V�vm�}�W��Jq����wն�����8�3p��>�w����|=�� �d��,`�D�K�.��"���'�6:��.�7w��IRq�����΃V^�`P=� u=~��ނ��U�ov� �� L����n�<����t����-|�����=����Q:����!���>�ͻ� � ��?�O+mG_���;������v���+�)�h�%������#1Qr��e���[nAss3"UL),D��X��u� �/l���N>��;�{���m;���	"ٰqX�����ի'��=��]d<"ws���P��,c�M�<F~�9Ax�ew1_(
އ��p��.�X7�d�E�$p'&s��3T?f�q!���C��CR�:��;h�z�Y�-tO|`i,��td�߿�֭�֭[A�&� Ջ�f�"���zֳn`�����f��7�����}���n������rmג��W�5�~&ҵ�YW5����;�ێ�0_�^O�c�x��;���� ��d|7�Bv�>z�]�^�w���ꃺ���C���T�q<��煮/��9��>
{w��;}�(C$���:#`u��wc͚5i%rIa���?��wV�ְ@zP����yQ�.��T~�Vb���nۋ5sb;HAd8L����_�I�+��\{ɩ�^��[~�rҷ=uJ^h�y�Ȱ�{��/���¦]� � &7��9������*�r�jq����1�����ͱ��He~1����o��a��F&�T����-���J��AD�d�dc��%�M��k�N:��H6���V��Nr��&�V�8E�F�s���;߮<�2Ĳs��s��\�"g��=m8�����HH�NL�C��S����sdLjq�-f��T.1{�v�z�=V��OA{�Y�w���7ߌ={�� �Iq�Lí}���)Sh�f�����)6�E��b��B��|���qvm7���S�\ەhH�k���ǎ��졦,soGCl��
��b.~��vU�s��~s��zv5]:���y�]^/��[�v�O"uq��.�=Q��Q��o,\��B���Flz�]�ڹ�,���p�u�)V���K K-r���]l���vq�2DzP��u�I�r�<��+�F4̡a	Lx9<2�ށ!&��9����	A������'.Kq;����C=����"�L-�ų���"��` sgNE:��݇��A�!/'�iS��G��>AaN�������A)o��/��@x�g��=�O�9Cٽ��ˇ{�ʵ����a���Y��#֯_���>D2a���h�R�,-AD<a�s�SG[�!t�W[o��	"Y��������ߎ3�<�̰b�h�e�+󅬢`����s��M�n��,�'��z�4!��o�����0�W}�����r���vu�*�s�g���i��L��S2��~�!n��444� �EɬR,]�e�ч8�Dn>�9����]ۥz��Vs�e��D�������$�b�Lخ��T~u�^<\�]
k��Bl� �%����>v��x���oG�?�vu=W��ǵ]� ƶ7�����8A��r�7�r�q��8?T�tn�rm׌o�e�,a���}��3�s>�WŻ＃�����QD����7��N�+C"E�"�Xi�F���ӭd���]re�T�,��;�;�+X���*.v���a���"����|����՟Ƽ�i����v��?���^~ã�/q������p�E�`IE�Q�x��<�[����{�������5�t����o|uM� �xS������4��휛��	��߂��u;��3QE�9�<~��q�q��4�t�[��k|�	di��O��`���������{� �T��x���9�s{0,j��oc�H��	�`����^��Tc%#/q�K/����CC�02�<؃35K��y�{�$� ҃���8���`嚣�k���ڍ�!�ɡ�����s�!3,�nc,Y�6�
���ݾ���<�w>Qe�e9��^K0�hv�&�H=$p'&ǖ�߲'������#�b^0"v�tj���ܹ���۷�h�w�	ڗ��pn��8n�=�����˵=\S^ٱ~b\���IqmWvJø]��n��v�f	��#���\۝N����w<��=|�|����vݟ�|.H;��|U�u���\�}w(�.�Aq��e��d��������q~���יQ<��uN<�d���&��λ��!X�[�w�qǸ]�p�I]��(�u���T�\ /���W/w��O��U�+COG+�V����{���|�/W:���@��=w}�l\u�q��~���܏�E�����Ū�2Gyy�4<}�e�����g^݄tᴣk��-�ή����<�t�U���'Q{�/����۾��WT"a����ع�0v�o&��=����x�p�'�������G��g���*���ጣq��V��_���W5��	�0a�>�PԊ�^&Bu;�g�$n
�v/��(�l���!�R��X�t�G�;�����^0��### �d���ՋaѲ%���AD��/��QǮ1t�{�b������h�a����/L+��H����m��Y2S$c���.���o�g�Y'��<� �2�/�a�����~/����)���Ǒ��}�����=z���|��k����#���T���|�o������"��]�����������:�ͩ�����y�+�ӥ:�C,+�U�g%��/�Z��k�����v�R}��^�vYoK�Ocpm����x	Wv�[���?q;�z�sm��bu>פ��E��y���4i�]�����:b7���pHW�]�V��H:�cqm�z@zo��E9&��w-�]),,�)�~Ǟp�mق���-z�H(�����l䀳�>;�E���r������ŝ��_m'w�#C@�Ƞ[.�^w�ɝ;2�ߏ��a����L�/�����ϒ�]dѼ�������x���b�s�'��_?��x���q�v�6����kj��͗b�te�̩�9t��?Ǉ�� �.�b��8n�<d2��9x캋q΍���~��D������D�/�u%>s�hh� ?J�O�S�.�ы�#K2��mW���W��w�A��_=���N��Q�}:�[�C������"ve���m��HA{<s����Ƴ�>�x�F�$��.\�Ջ"+�FM#br��k.]b<t���;�lCwW"�0��~��ƽ�E]��o�C�0Q�_���Bwݺ�����W1O��G�/�&p�Ŝax����[3���H)��"0��i����9�vo��� �ۃ.q{��r�da�+P�)l7zQ�H���x�O"�dmٲ��777� s`�Y�KV,Gn^���L���^���ZU"�����z*Q�؀ ��pmw����4Kծ�
'x=�X^(W�5��:��a������[E�K
!�s��um��w�&��u>w�s}򹠉���k?� �U-Z�P����wm��>o]�����q4���+y�k�q'��k�`�����EoO"���l�ڵ%r�$xO,���H.�r���ێ����`���Sl��t�.�la� �rg�{���Ŋ���!��0Q���L
���Y�)n��/֦Z�~�1�>���vά�xq㕸�'I�N�&X����ql���9˫f�o���=�"�Đ�"�t�s�'���*�Ǒs���m_@���u�:~�iB�� &='��F_K��7
yC��}�v�˯{��/�G}�̱&^�/��_��x衇H�N$���%X�r9��+OQ�� "2잣�z*Ta}v��m4�"�8��9L��\�/��Ҵ�{�:��QK���Z
��x<ͱc�F�{��BW[^��7�hID�H��AD��� zZ[� U�����]N�R��L^0��X�ڼy3n��&���8~��
?�=Y��=RE*�Ͽ+�D��l~uj/6��b����PԶb�ctd4J��TXnQ��ha���O"X�����кYf�˷���@ +����/�Gپ:W����*��έ;֮r&?�qe�dl�튦��pe�3ʎ����!5��.��-�V�s��c�}��������h�Q/�_M<��ύ=�=:��uٵ�ѧ�����st��}�L�;~�v���xpB�3��GFGB��/������y|�4i�'�Q�d�R,Z��v~����d&�o�����u�>�,`u�w��\W��H*K����%����Uve��T�1�e^n�^.�V�:��;�n�= ��!�	"��1���s�-�_|����@"w"v�P�?��,.�D�SW�/���?�"1d��=��&r����=�}�H�>�_:O�r	��� ��Q�g�S���ͱ���ͱ<��nc�(�����)z�I�p݋t�/2X<�'��~��1�A��	ۗ�Za�	� 2v/1��Ҙl����C[K+"�{�|��^q����$:��Dn�)r7J�eJwV?��{��a�w1�(�ٲy��7���d�E����~��������Xbv9@���G�J=���s���r�2cx����z��w�~�z��� //񀋾R%|c�3U�r�l���g7@�ھ����;sV)f�)CNnz���)���#�L�<���)L�PiKU4��H˭m۳�ѹ���$J��zh��t*�u]]nm�7�Gt���׹f�?�v������sn0�p�[��k��
:mvN57���w��6]�Q=M1�t��@cc�}�v��Z�>���j��v�w���]�]��<4ڊ7��ѫ�췣��A���<T>x��$�ϡ��Qt�����Σ���a�w���C~~��7ԇ�o>`�\R�[�ީr�a��{����=�������k�g>�q�"zR-N�׼����o�f~sٱc�Qte�B���:U�3�틎b Jpl�
XqW��ĂV�-qzU�TG��Μq�"<~��2J�αD��;� �2mJ���
�h.&"�|�ll�sИ�Đi"�L�s�1'��I�>>}�r<���d�o<A��@�o��fu��+�Q��	V�%n�#B���Ja�%^�"w��-ng�g+Ѣ�L�/2X��?�)~��g<`��M*He<����~:�RU�/�6���a�̙�����?����m���a��;K�~e���;;12<��޾�l?��>22����m�����[�J�N�}������$� �������v�kH�'���s]P�̩ؾ���T��c����x��=]��ݾh�%�ew)o��_�y����/s�f.P�e�%����!�1����;��,(:Fd$�9YX<��р��EG�H��*W��3@�v`H�z<D�j����2��;:��7��8�Ͽ�/50�z�����qO�O�;��=�D͒�X�b�!d��o�8�۰�݀�|Y�`֜2��)zSiX�:�RD��jn�����d]^5_����&D/S�I՟��A̫�p�Ŷ\}���y}���6��n�Kf�:��ɵݵ?R���0*j�؎�x��[��b��ja]�ٵ�%@W}nBف}�Q8m*�M�f�I����Z�Spc�ك%�,Q�Gҹ��y�Br=j������e�<�7��QM�H!l�I.3��֑����ĩ�lۆ���/F�<Y��]��}�@
�����;φd���.��D�>E�&�`2�ijw�`-oG|��#��:�+_�V<@%�1�)�]��P�F"w�HG�Б	��1S)�6/l�"��	�0q��q���3�����g^���A$�L�g����D�υ��>�����{t"���Oĝ_:�tj#"&�� =�m֨��>G}���b�0(�����\�?�v�������;LF~��rK?�����c�!��8H�rWl?S��#�d�w�}�:˙^\l�SJf�J��y�:'/5F1욗�m�z����ܜIy�#,қ��g��HY)2"Sw��H�hJ�_:�,t�Eu�"��p7:B�J�f����բ$j��o]�`#�����+_���l��э�4��Frq�m�r��]����`0���.	�{�[pւ*�~/��ɇ�DF�v� z��M����0����AZ�.� l�����ʅ����XĽ�؞���7�4�흝� �xR�x!��^���|K������̑���w?2�K�m���y�=����-�b��^� ؽ&�r����B�+mǫ��-nW�ý⮺J���7��ۅG�C$��ˌ}�e�U�ե��9=J=��!��~)>_�9C ��z=�}W
୾kR���P�� ��)nW}w�A���!���p}�=X��#��C�m�yM�X�6���^�+W`������ X@��{�5~�>���&$�$���x��}����bpc��/��]X��Eq��R�1����#8v�a��,��h��A���v����c{=��	o&�s�HU�<�������8����;�»���=���s���ƫp�m$r�C0��{��W�},���Us�1ں�l;o��Aר�YR�0�-lW�`��v3�ǅ�$n��>�C���?��?�x�>����	�X��m?�s6U�O�3X��[Lоb�*���Nڶ����x s�O���l۩�>s�RX���))�~*�}xh}��O����;P8�����T{3ޯ��;?��Ҙ���m5���E*���>k��ֱ�'C��x��G��x��ER��׼h�e;����^Bw�C���rѻ�kR:���A{ ���K��acɅ�D�qFuݭ��ӝ�ク�A�1808VQ�����)��+���T{,A�M�6��[o%q;7�w��r>��gb��eVY,�	�u�"x��J[���:8���C+�ϕ���m�I ,�����*�/oRզB��*��+��
�=l�s�@\W��Z�c��OA#�藏�x�]�k����R��q~hb�z����s�}���Ƈ��k������Ֆ.���<���v���n<5i���Sף�	o����x��;�#�(�R t���c�r�Jl۲y���O��91�`����ϸ7fN�vU�Iu *�~���G�"�����1�n�VG�E7w/76��t��ixiWj��$��yY�G��ف��4E�W��۞$�;�dza��}T͜����p��y�F�+V��*�YT>�6�?y9�|�����z���`^�Z�Lႏ�0��~au��r|����y��A�Ω�k�ܙ�{S�ܽ����Ǯ�g���9A����jЈ�@�!l��ޮ���g�F}��da�Cܮ�ٌ�̱�C����x�b�D�ۉ�Mn^.V�Y�yU ��,̞;ǘlw6���/����_�*���K�n��R��~A6�b.�����B�aV �0�\6�R�#����+s��/�����N$�E� r;k�%
�E�����2H���m�AU��^��j�/�x��A�͛7�n@kk+"̚S����iӧ���ݖ�ݿ���e�zItm�b;
�xF��{��XW�)���U�-��]MK�
vَ��\��\m��ޡ�������.w>w-�����j�N9��z����U���p=���-]%Z�<�����{��%$w�]�ﰲ�C��(?��8?T�)
��ڮE�>z���òU+���w���H�S��ą��ٽ�\�T1z$R#`����i���iJ��j�A���ܙ��� �{�H��E71`�xN���_�zA��	^x�EJ�Ι9���3'��A�EL��E��.������������0~ے�>}�e�Ȋ�q�s�?���w�ǖ=�*���u��[d
O����������9�.N�I��1D�w]��n}�D�
ʊ��ԭ��t�#��Y���>h8T}��l��W�7��\�y�P%l�m�gL(q�L<�eq���G$n'�ʔ�)X�r�#q;A�����yg��~�nڌ��D<`"wvo��/9a"w�T��3��3�}��������n��ϑ��9�5�`�5�߇s*���n�Ƀ�6"c�]��+:��^�rk�
R�V��=R� ��u�[�.��T6*��4�2���֭[q��ד������kV��d�U6�]�òXw7#	��6����>"
����Cخ�OO�v�G�J�v(��k���[�n���{�]S�E��.���<����d����Ӫ�j�1���Oa]���＼|�t��X�z�z��x��M����������kצ��B2�=X��r�5�};��,8$�2�`���۴E�b��^�D���2x
�E'!`5s`f����"U|�����5!��#*0��Kw]e�L7�N'e"uL/�3ܵc}��+�?�?����w`����Zw)>zԂ1�ÄΏ]w1θ�1����{�s럊Y�Μ���+R.r���vN�ܙ����uO�����e����m_@y�T16Ψ���	9�Q�-�`��=�s{Б+�D.q�۽G|�f�%��+��I�_2�*q�O~����?Aă��,;j%�V�׺]{@1�a�%�A���P�{/�oي��~�x���7��ϯ�⊄��3I��c,9_��K��9Ckh#ox�a�%�]9C�,<�۲�V-�kud�E$�ù�:�Z�� UPREpa0�� U�%n����rb��0q)n߾};n��F��h�T�X}��q�}�ĸ�×^�*d���&صݵ}�(W)�7�
!���{
x�y��S���S,��K,=�vc[.���?�O���յ=�~T�v�s
1��<R�����������wK���h��~�.���}1�)��Q�x�ßk;;��_O��y�MZO���0�h*�\�)w�	x��~�1V���p�=���g�yfZ���u���M¿��¯Ztw.xw��Eѻ������� Λ�-w�jpp���๽ "�\���x�;"��!w��ڌT����:��پ��f���~m��K1s���X^5��:�]}�|�/�iW�]���q�ݿ��}��b�t���'��L�����-�ണkb^��W6%���[2߼�C��&r>����'�ߨ��Ǐ�ƿ��9��=� �FŴ r;�Q�-a�Os,y�g�e��˿{;�	q�r��H��=��S�����1^�)�ңVb�E�
��w!��,�{���QQ]��;vb���1<D�ネ���/��҄���
ʓ+Z��͈�X�\�c,ކ���'s��˞Wb9\�]Y9��S��S�p��D�D�!�;��.b�ew��\u�*�C��
#�ۣ;0h^����C:Γ|�&ng��MM��&�{�s�ꕡ?�9n�3���) ���%���WJ��rgOm�K+���Gj4�vQ�X�tnõu.V�g�]��s���vR�ڮ��q�\�5Y �X�5�k��ϱ����{�:���Q�X�� ���8]��:�Ee͋�����3�q����	���?���Ac�9��_���-��'?I"��+�$�j1`�_�C�^�*�2_�XY*���!j�WG���8����`A$�>���gb��t�"���J~���xrݥ�W:��:3�����3'�]��>an�/l��p6�˾C�t���ݘ>�	L�~�]����\jY��U�:���8����&r����йq��"��͝x���0kF��u�/�w^i���o�d�g����v��� M �w�	���ߣY�X�ܵ=�)�רϼ�;wY�M�nbF��=��X� ��E�xꩧ���?��ILl�w����8z5r��2� �h�{��+W�z�B�ܶ�>�a�.�X`���c$[�az$�3�6�r	�a�y;�+���e�.c�.�G�xb������씙�x���8� 	܉�gJ���&�cR��vS�΅�{�,n���1��Q0� JO��]�ߵkn��8@	kbl����eK�?��sW@���S�ڮ��U��.�c���(���mE�;��u�rY.��\H�k�����>j�e�rx;Q]�5�W��<����|���õ]�S�Br���N�{��יl�r_�k�k۪��~���z:7�v�mM<n�`hB�xϘ;>.�WaǶ�x�OBwW7"Vp������~�� R���ɞ���Ќ%cv���@�s�A;h�P^NUx
t֢r�Է�ȝ ��g>���Ӆ1�ߘ`���R/ngl�kƙ�����9|dE����M�ó����p�&��X��-]���'�{�104�+����8��cj�9d_}�)����A�'SD����������_�-e�v�{�c|�M��앳g�^oIE)~u�U���P{&_=�Dl�ҧ|�l�͹5:z[;g�l��=�)V�Q�M1��Q���+_(�Ϳ�U�X��K�y����'q;1n��+����)E��#� Lrrs�꘣����mނ�u ����J>��q�|�%�P�з1��8���ce)^���9� r���]vr�r�R���gWO��{�A"����H{ήF[��
z�Da�������gx�D;0D#�L����L�~�uס���D��"k���/(p-�/lO�k�R���{�`����v�8�7�\�\7�MC�?V�*�v�=�������r]���vm7�";��c��O]Ѧ����'�ZW��D�*�v�8[��v�1V��5���_
�����rm�r����޸��������L�]ۭ�T��{Ͷ���X���,��o��7��W�� b����pr�����'��cB��H񜏴��ί��;�DvPR�6mA���Õ!�ҝ.�`�J���<�㧵a�4�R�� ʅ[�G�sᘜ��E��i��3����y���վ�3D���L����Sgg&~�KS[7.�����s��G�����Oo�<>y��1�qř��__x[�!�XHw�{�:��44w��c\3w����+1db"w�;1`���^y�y�� b|,+b�u����5�s�����]��QG}vc��Y��yD�����yղ^x��?��c��d&V����?0KA�)�:'��QZԄ-߄��vD�����z��^p����t��z�)rg�Ǉ������ +�1�S�.�ܭџ�������a�5�V��3`w�("Q���HkN(�FoK�ہAZ���a�{�R��^0]b!��6��ۇ�n��x%�X�1�kN8ť%�S���<�/���F��õ��u�z�׵�-���k�������k�S�<v�sޖ�<�-��}S|��z��{��K�%ӵ�%�������1�]U�e~��:�P�v�?��%lZ)���j��3�r�ǰ�c����M�����X�n���pL�<�(<��X�k�5�"m�[W��T���=R����]܍���+6�vv`m�4�v�H_8�h<���M�HGq;�	|�������&����|�[�����Q2m�����w`�o���?�:84�������ŧNX������;�$l��+ b#]E���.�x������������^����B�{��?��"w�����v.?s��A�r�0�;W�gyC/S,[�p�����G}VO���W��I�y*��/����^���8����)S��أ1��AD|�5��<�l4���w��@?"���q�=����sN���W4�:Y���smAX�ȷ�����2��]��|��34���B�Φ�ZP�>��*� H�N�-�Y(i�/a�5p�/���'�C�HT?>�;���� �X`�,?zj�,v����k����*��"Xq���W)P�M�.�]��1����f���
a���K�.W��EBre]���SW��)�v�I�Tۚ���~�Ӑ�Õby(����{i����.���������/��5g�z��q�qlT}ڒ���Y�ӵ=�-���En�:nN!��������?sHe�}
����_��)����g��+�Z�W^��6� ���ى�o��pfX�bE܂=�h��v��|�}ݓ��<`��BW���̕!,xծ�a��Y�j��KKj���Fx �x3��"?��7����^w�!��^��i�}�~�Y3
���+Gg��ߥ|�E�_�9���#�����ǿ��9�u��׿�S���Ͽ��J$�J��ܙ���?�3�[�Lܾ��@�q���8ƿ����_�W�6n���'��=1�m�y��p�G�� ��sN��[��������b���AK䞌Q���1�<_:��㙻����+$n'���.\��V�]H�B�(ؽLeM5�++���رu��B��oܸ�����'>�+?���x���c3Ɗ$t7G~s��P�=����B�nc�t����nDB��|"m���>�����T��]���],a{��)nD��ہ!�H��g"�[o�;v� A��}�Vc�Ն����ο�o&�z��,zU���F=����\݀-Z�k��O��X-�w�G!(�ۊ�w��ڽ;TN�\~����vI�5+� 
�ݮ����v�}7߹�Ϣ�PO~����ӵ��٫�ݿk����D�&��#�Q��r��9]�=�7�nWQ��nh�����k����O�;m��ֶ�����:��D��r\��/aۖ-��W�����)< �{��[n1��.\�Dw����@�S����,(v�nP�vrgx�ۙ+���]��� U�`��5�<� j���wFDt���_?o�9|w7ο����KQ1۟ӯ!2]�!r�D��o]tJL�v�??�g��·�4�h_��9������ĥ1�[���sNZ�g^�"v�������W�~�������˱���ҏ�� ���19�?��i��.S{����^�������xn����>���������y���A��5s���9��]�����}��>K�X<W��!�W .�.y����7�����o��"��+���Ea����� ����^���*����qp��_�~�z��OW>0]���cTc,�w��	Bw�����\����N��������qpp���KQD��X���Ob��~&��t{A�[�%ƈhc,1�رDA�F�*R�(W����3�3󴙝�{��7��vg�y�;�3�;��g>��/r��Y4����Gk�z��3�m���D�!�;��;(��[}<����]������#M�x��܌+��o��&���AA����&O@�JU��k{x� m�iT�vYt*��U�f��W�;"DU�tEq�{��vS�S'��t`����)��6<��3Ko���.t�6�v(�T��\��퐘k�鬔�&��YyU��ۿL[�m�m�.l]�\_�x�]�FHȵ��ݳ��,��b���l7�!]�w���~�v����E:~ŵ����د�|��P��CǍÐa���/��7���ƍq��c��0`@�N�����䞏7[�҉�M˝Nuq����w��}o�����c�@D�3{<n��r^�n����;-'�ic���S�%�<��Ex��u r� ��~��^@G�9��w�#��_�btt��$�N"��j����{yp��������^<��ۗ����v6��7�y��l��������xnX�+N�Օ���l��H�.%��p R,�ꆶ9�W�woq��	����#���d�۳I �����ۖ1ց@A�\Qa	����� "3�s�c�ƖM�-�{cC#"���V�����=Ǝ�qy*E��ZNl"w��S7���\���C�k���y'w�џ���&�|��>-��V݁H.$p'��>!�7m l1{�����=| ��*���&���T�td�(=Y��]xW_}5�.]
�BiY�0jj��>����G.�X��ڮ�s�k;08m�fS�ڮ��%��,'k]��-�C̵]��H�Y����/���W���_D�����Z�ݐ&)��!L3M��w\���"��W{l�!�w���&����1y����\��,��]����	����sg���I;n��Ǔ���VD4V�Ze%���{uuu���{'��dw��g�����*���IX	.�19qr߻c#����ɑ� �����<��0��W܏�ߙ�o�41�<�J��𒯑�=�a_u���/l�]h�M�?؆�-X����|���<H�DaN�]~�"�Da��{~s:��0,�y�����<��;?����)������'�=+��gcH�*�f�߇杭�{{W?�����v�{{&F}�T�.Y$3��?����џ��;���>#ǎvrbADfa�i����?���>짛ֈ����㷿�-n��&6,�&S�ɾ�����!�]Ï���|��~"w��.�
�ڠ�fȮ�t��}��avM+]Mrd"��Ed̩pz�.47�(..R����RT�;KL����{�	�ˁ���N�"V��9s]�����3π �0pH�%n/.QݱbumG\�k��?v���ѩ��K+ί���?T���	�u����$mw)�e�q"7]��<�S�rrf)T}[��W����M�>��m�D���
R<�45v�g�sm���ziں�+�,~�v�_��4B�X\�����ƦG��͵]Z��S��Ը�ێ�rLr?�^��.�e�sl�~}���V��.���������zp����ҥK�D��{=���C�+a%'��iz��;�`4w/�;��P�M���7�Z:�А 2Eiq!n��]��l�Մ�\z>ٸ��p៟Ƨ[�qŷf#�ɛ��o��1�����?>޸�W����L�~�����O�>:j�U�v���,�8L�~�s��G_>2m�<�������ث¹]fQ����������4s;g7=����Q>������� �Ì�B4�Xg��\$�ci̱��aaH5�*�ܨ�:�������֭�DM[�nM���}�����Љn� ��:�o�cF������[�|sn�m�Բe�\t�E����z�gb��t5�w}�������K�n��lJuC{���X���1u����nv!�	܉�b����$�Nܮs`p���v�J+n�=Q�i�hdCRJ�}y�z�X�d	"]�Ub��I���y���T���n��b,z��]�Mh����µ]GZ]�q{j]�݆Fd�I.ں�Z��<-�B1��kE��Ivmw7��Ov?_e_T�3|lhb����n��˓��������'v�Q���4h��cCwA��k; �d"n7S�F]�׺�?w�˖�uΝ��C�7��sO?�O>��ǲeˬ�����Z˝+Ӊ�L�ٽ��"ww���Vr������%r�Vm\�JrP��p0򷵥'؏���@q��\�\�����c��:��_A��Ҩ�+;��Oִ�'�����̺���3�x�۸mθr!��4�Hmi �<2�<�*�v@q����q�϶�����K���]:� ��P]^��{�[�>y���3�r��B���:�F}֑5�T=߼y3~��`��� �h���4� A�ݰ��w4�lڌ�����͔� �Y�f�%r_�`z��l�fK]�����sK���!<j��߰ȝ5���S74#uC}������l݈ne��s/�DI$�@YC��!�v�C�-h�PEA;�����ݝN>y��u��с!R���Һ뮻�׿��}G�א���e*	*��bHص�PE���zi��S+a�BaE�nǭt���.	���Ʈn]Pn�h��3K�$��݀# ��CX�n9nGB;S�N�{?K����Z�ݐfW��~��V��]�u���c�������.�3"q�X5��u��<������e���Ƶ]]W�7� �y<��د-l�	�v�S�<�?Ye	ݛ��@^�����?L�Ά�tB)�DO�c���c�qc�V�����}���7��NN�D�V��'����L!A%'�t���1��P��e?�H-�(n���۫��܃�.:��v�m��L#��+��B��D�?��c��z�r��Žۿ���p��`1��l�?�����n�%�qh-��t.+A�cf�&4�jci��^�f(�a�<j�Y7곎l�'򼮮���Z�
�;������nn!� :lԍ�_����a�G�� �X�r%.��b�p��֭��N�-uE_c,��uJ[�S��k�����;����Z�%n���k���[[Zp\�}xd�G��@w"+`����w�y��$��^�Ђ��U�A������ rǁ!�.�'���w�	��W�>?e�u7�������hFo��k{�m�|������kgֈ[���Z/���N�̉����e�:���Vl�퐦vm��k���ѵ5�.�C�/	���.W�|���D/L�vm�֋�������F�0v��7+��!��)��=f�� �D+$�C��u�)qm�n#gk:�(�+�p/���uس{7�\�:'�|UUU��l�^��QM�.�;Ye�ݳð���_YܮzP'r;3r	���#����Α�~�&|R�����@�䞧��Iq�ͪM;p���]�>�
zq�So��O�u��v���g7?�K�z=������Z`ۮF�m���v��Ȝq�a�tH�8�~�1��O��BHO��F�ƈ�jD>s��B4�oEqI��v�qo����υ��]��T#�,�9�"b�z��ЀK/�+V� A�Qٽ�5�s�U � :&E��7�R�寿E�X�/o��6���J\s�5�ԩSƅ���S�[ߠ1�Bd����o�g޵ݒOp"w����ꆼ�ݳfx���3L�7�6 A$
	܉����B4�ׅ$���h��"r���u�Ar`�|�ҥ�+���/-���.hƎ��Çjߏյ=�`=�ފ!a�vM:[����sm��wm��Iڎ=Ů��[�tN�,u��v~}LCޞ��r�յ]��1qmwo�5�6е��%��$vg�ܿFH���Ǖ���<�=V���|��Cjd W]��e[7���eC>�	s�X���%ر=wExDb��~*++q��
��Չ��.?G%a��5�]��I,�����E�vM�ud��T�ߖ�V̮iţ�)�@Db�j܋3�\��ߙ�o�4Qy��'�Ꮛ_���l�����Z���|i�(��Ó��b��:q���IY_v�˵���<�
���; �|�{�tٻm�EQG|V!�9V<�CY؞ͣ>G#�u���V̟?˖-AxQXT�1��Ð�Җ$� RKe��8d0���������_�~/�"�N0�<�%��X�)���s����t5C[����n	�պ����]/��lDeY��K�=�Ty&2N�J6 ��]#nW\�ei�A9)�� /�����_Q�9�2�-�� ��{�=\}��طoBG��}-煲N�a�c�#�L���M��ڮ���յҙ�S��.'~�vY��N���r[9N?�v���k���q�֬G������ns>����s����1Y��F�����`�ُ�8��v�����NM�6����k���o��$M3�s
��	m<�ùI!�k;߯rc���v�y��E�~���e������Ժ�%�[n����8餓2��ʤ���ا��KXy9�&�9�s�FU��{[�폃���;6��>C��r�%"1lÅ~m؆k�;���������%���_v7�� ���S��?��u��~~�Q��YG'����p������@pl�f4�<6Ɗ�����{{dZH�%�#=�C/�v�G8�ٱF}�F����7�|3�~�i�=z�Ąi�ѹ�ADn�~#}�����^{�?�
���F�����?�AJF��l�%�"�0�{���0Tc,�����}�5B� ˴����B���]7Z3�---8�_�1� �gFu�w�(..SE>	*G�n'�
݄��P��+Bw;	%%�\�d�w�JG���?��S\xᅨ��AȰc�9/5B��-l,n�,��hPvM��kD�B;,��mՋ��0Uq�:gx��Fl��.x� %v�}��#t��CS
\��vnx40M��Fb���JqM�(���>_Av��fx��vS�8�x"�;���k�C��]=���}�8�Lӣ���M����ekjL���4�6P�p+����\+��ҝ'����,"W�>m���ۇ��L�y��'}۶RҊan��Ȯ]�bڴi�gR��{&7_���M���9NL��ΰ�m��=t��C2�����G�������������>߉�f7�;�F� ��'����jވ�u�L����V�قo��;6m�� �i5�h���%���vχ�s{AD��ݣ>g�Η,���~.A�(*.��q�bȈ�q��� ����i������x�o��~*"*��s�U3��׿��H]&�ꊉcI���b�e�4�3�3_#�k���=,n?�u�(.�RݐՀ�vlƤ~C��f���Cw"�[BC�������$�Tn�AA���������ޮKT%!I�#WE�۶m��_��>�!ӧ?��D�>������ 8?�����+K�P�v��FT�Jm�\�����R��.^=��r����hp����'͵]3��$��.Ϋ���.']���x��έ���F��ڵ���p��#5N�硉=�k��=L�6�����!hc4u}k>s6�����n�/�{]R��n��r>]����������?�^y���	6���_�?��=ztƓK��MhɎ�C:r���eX�����$�=�nPv��������=�`�_;iղ�'֚xl��v#������A0��H��J�9|��˯�(O���}~vڌ�����m�Z�� �M�ʲ�Z6����1��=���uuC}�0�{{�G}Nv�|��O��nA�`B�#�MF��rA����Cѫoo���ױ���	l�g��>g�dS�0�uE[���ٵ��Y�/,������eq�m�řbEj�Q]ܹ��=�_�&���FSK�o�%����<����F�����'�d��B;!%&��\<U��v��&��T*�E�HU�����%}��G ���b��2	����M���GK���DU&��O\N$BUt*�����{��.�vy]ൎ^�=��J�N��Ĕ"�vqY�g�r$ߵ���MH����'���ihb������n�c��#i?T���i��I����*�V�i�Mb���~m�ѵ]����E��~f�6��5�.�6��q�/,,�Ga���x�n����ĒV5559�tJ�o_G�?�IX�N�^Cڂv1iŹ4pN�m'�X]��n_��zÊ�ɑ� �H.e�E "��9n0�z�(.
!�a?��~{�;yr�}����w>��Ͻ� \f�ۋ���(f�X��~�v�n��e�{ �v��%��k��T�ԓ�_:����K���,�F��)*.�������A�Iy��8*���������TK \��0w�\TVVb����f^�.��cYF��g���Y�U+��c��p}P�D����h϶)�麵{���hiiŜ�xtU�獈�@w"cݫM������so�%���۩]NT���;���v_��Ƽ�G:D2*���~X̛7���:����O�6e�ʴ�̵]'�T��d����ku~3�O��P�nq+�gXCTl���4�^+���k��rL�޵=��Aq`�v�ێ�ą��ŋ��vIvm��|�l����x�ͮ����R_[ǆ܆#p���"�,��(�caߐ��X\�}���F2�����~��{Ӛ���ǋ�΅�;s�}[l��4ͱf۽D��gajڨ󙦦/ݱyC���F�z��y?�>^^�b���ͦM���n��&TUU�=�ēM	-�|˝[��uN�;2D��#��B�;a�qqg�!�-���-�!� �e� "{�2������~���־��_��g�O���;q�5b�*� x�(D��uV�Ppo�e)�nX����������9�5�l��������+�w�^O��}0��)V�pݪ5 � 򛰛{���kؾu¦���]v�5��ȑ#�R�Γ�Z��1�S7����j��z!���L��Q���(Ϧ�1�3_/�\ܛ�o���C��gt3;��u$����P��%�Jr�(��]v`pU�DU���˽��a���D#��)�J@�}	����ǳ�>��a����b��C�?��ƵP��V�4��k�j��rm�Ϥ�[��Z�fZ,��i��fDTۢpZ�'��q����������a;�z��Wi�Z��1��%ϵ��A�凧��ڮo#n� Br;ص]8^4}����d�m���9 �p�2�e;�aM�_ &�v��-lcbE�cf�!Æb�#��k�.c�ʕ�ꪫ,����ҬL4Ų�d������pn�Vq;2���&����U�ZN���܌jM,Y� �H�:�� ��`�!��eg�Si*0����7.�>X���{���A.%��z!g�U$	��q�[���fXќ۽��M�k��HG�q�����K����&Z� ��_�;�c�YX���x��w��A0�o�nc1�{���3*f��Z"_���	9c,�nh8}�źaA�^X�&:����{,.�������Z����i�[Y�6�G[a�ց�NJ��0�!7Y�sm��W~�����;0���]~�h�"<��� ��=�0q�TTt�}���sj+
���?�y�6� ���z�`��5��b�J� X�����{	x�������v�^��˵J�����!��4Vד�Hk����"i�]p�v1�3/�sh�Eqm���nv��&����>֔��v�җ�3�/��؅�H'n�쳺����Wq�VH.k^Bri_�ɵ�	)E�����������&��u�X9S��h]
Є;��j��~�C���g�Λo� l�o����o������V�]A�����'w;a���OVX�GΕA�����5����Q=o? � �HU];� ��3aD,��l�����
L�~ӏO����p_�y{5��`1�[@���-�[ߊ�bo�vOq��n�������Y;��4��&�͑���T/��ڙ�}Æ �h�C� �`9={��/��]�;A�O?�W\q�U7���["����YK���	axG����>�uP�O�fh/�]/�k��������Q3tD�]7liه��U �X �;�v���;�P\\�80��0J�цԹ0x����줔����7a�QPA�?�������`��gب�=�P빌�&?Ln�v��+z��"r�5��e`!�03�mլc�iU\�*�U�OMԵ]I{��)n�c������ ^v�T���P����sC3���څ��<vg�;���S>y_0����Wi�{6���p޹��cP���\��(m��b�v�uyz�}�\�q�ǲ�󰦍�/���.��v����h���y��&��)'c�C��Ë-�g�X�x���p��M������X�s���WF�I����	���'��_7Q�2�ޮ��<����Xmt����	� �Օ "���/=��r_�^*��~�U|q�!	�u�o಻�����9�_!�v����ݯf�<��a�X;�cy���bzs,F*�:�%z�g�---�7o�5:A0��	� B�KeW{�|��J|���q�f!r���~�_=.��2���h�'�j�:c,�t56��{�uW3�E=|%��,
�M� �K��y���5�o��
	܉�rx�"4֭��9�ǽ�ׅ� ��B!���/�&�d�v'Q��b'���T6ٔ�Je���>��JR��O_8й��fi90�H�k{���sr3Sjc��T���V�_����R�v�vN��S{
۵Bx9&/�vS�3m��ܼ��y�rm7�MWT�l�\�5면K�k;?_$��������M���=���.�^��|e��ej�U�6
�Fخ�l/Z]���Q/�ר�Muy~}��L)�aÇ�����=�֭Y"�a���7ߌ�}�b֬Y9%fO�?��gw�92�U���a�����JT����M{vcVmw<���AD��Mw��$cj{㑫���Υ�u�
C��W_ŉ�G&�ρ�m��g�i�2��Q\��h	���~#?�$Q{ac,�v���˵C��fMܞ��]2�H���a�X�� ]�`⴩��C� ����6u�X���o��M�� ���z
}���~�m�,���d�Zy�K�1_?T�^�B�z�-~o3�a����m��R3�����Ë�⣂�8��	܉�Q2P[���v9)�9� �P����ON9mb*�$��l����[���+���$��kpđ�QTT��g���#�Dm��H��R#Ƅ���sm�*��
���ڮVUQ�:�-4��5XO������{��n��bqmW�����׳���@\�<�}AZ/����^��8_���}Í]�A�	�vV����;!%۵]����Rn^�z#��<��~�w��q��Z��i#�Y��&���� �'&n�WL�qη��7^}�~�_օ.���$��W_���jv�aJ̞���_L�#wHE�����:���î�+����c�As����-AA�0��'��Bh�O�)�nF���!�a登~u*�L�P?���;�?����A�9a���%%%��ݯ~�{�"w�+�׫n�-j��Q��G2�?���X�h�1pH-�<�:^	� "^z��Y_<��&6|�q��Z�?�r�)Y#f��|-�U!��0v;�n�U3O+����|�P#l����u�����mj���xj� �`�U�6N�5�I��(��B�D�΁�����5�톒��$l�Da���6�}Ē�
����f̝;�V��߰cm��0t���c�ۃ���E �-�Ř�����R[�4l����g��=��i|���W��!l�
�5b{h�Ŗ��(�e����Js��d��r;թ\��@r]��J� ������몾��5�h�Ь��.�ؕ�Hڷ�Ⱦ-�$��G��c53�5r��Ҿ�k; ��S�=�,+�k�܋�Y��6r<��uOӹ���s5'l��n��B폩ӧa���X��Cصs��eϞ=���Kq뭷b��Y�tJv�A�K�#������D�)
܅�F�~P����bz�f<�P� �H��]:�'L����:�H̹��W��n�/n�TZ��.:3�M��u���׮Z����QAxQ۽��ִ_O)5�"��aa�S�7�
�J�0�l0_Cd$Cl�|�&z_�t)~��߁ ���0~�D�� �H�eҌ#ѫ_K�~`��3ƚ?�e�u�Gvx1{���ͧ7�r�u4Y\ݐ��}��H�P7��j�e���Ba�g��}�z��Z�M��&�Cw"-��Tk�����E�CH���%�x'�{Ȃ7�t%���G���KP�X����H���bd
��0t��� �랬嗔�b`� ���a�⛖�Q�?�ٽ-��	��HZO�v��TC��=�h��k*57�D����ؿ�}�[���գ����O���ʳE&�޵׮c�cj�=kk@umwE�{ڗ�a���K����߷�ِe�564�M�W��5=����F��~'>]�Z]��צּ0M���D�s��0;����U���U�3|P�T���X�u�YW�ҲNڮ��ZYe���M\���G+?�ϧ���M��YF����8p� �����J�~���?A�,u�l�|+��mFqQ�FA�?ނ�cžt��[���wV�E�(�;���G��Wb�σE��ߊ� ���%���v�܉y���n@EEE\	�lJh�ۇ�}��;~���]N\y&�"�v{�A�V�����$�l�;{�P�S�k�� � �g�%/��F�ICTD:8lH<tE����vљ����}���p�Ջ�}W��îa'tى憐֭������a�h�ŋ����џ�ڡ"|w��:q{���td����?�F�ۿ�����=�,b�
AD�8����y��W�4�������+��m�݆!C�䬘=�X|�P���B�w�f�ꃦ��]�ٮ!��aj�n<�;1�!����H��D�@�
*���d�ށA�k��n��?I���ʄV�E���]w݅%K� ��d�޽���*SɶL�{2�_;|(ƌ;���'�k;;�*�wCIiI�"4�N�e��rϙ��_� �S����.�T�B;/�mX6��}�7�ك�޽�]ۃ��v���J�]�d�oݏ>5���((�՘���]9������_d���	/L�Ɔ~}tbg��4�bIl__Wg���^]-��S�)��/�bl��#ܚ9��(�����͐c��ئ��������C���؎���L�|�p���6nBE������n�m�{N�nY�2������6Kx����X\��I��`wӰ���}Vs\��KwR4\�;�n5��PVV�����0�e)��04��x��3q��ч8}��*����I�o3v�axoŻx�ɧ�^?����gɍL�ѿ���vg�e�~c���[�+�W\Uȟ.��L�!��;2��aDqd�v�MV(�*�mD���=E������"�:��Ž���[� "�`�֘�Wv.��~x�%%"�L:d ��,Tt���x������Ƅ����k��G��V�ͱ��а�><�s��X�C4�rM�x�,YԮ�*Y�ꅆv�]L��U��m߾���<\"�Xl�|^��Z��,w�	2iX���LpسOo��|����n�d�]u�X��e�k�km��;�2��Lo�L.����2�*̐^&ם��1Xk��'̌���5�F ��ٹ;c۞��z}Scfn�ϥc~��a��V���~߰ߏ�]�`��ڙ�ms�)�477c�ܹ�1ssOTp��Qk�"FDN�j-���Y茱���a�F��,cYm۬�a[[�qs���ȝ���7������xe������H9�*t�T��B,I*>A�&�D����������O&D���O~��SOY�d���2��n�Z~&�=�峡���:��(�E��X����c5TH��G�*����l_n����qS6��N����[�.����X�P!��k�5Br� V'�5�y�27��{Q��l��]#�Ո��mUq���`78�Ķ�J
�#M�־1EVH�*h��l�i�_�|�Y�)��~������w�I2~?Ҭ����\w�v�s3���`��=�]��=���~h����y��^�$���qG�Q�8Ӵ7}�/��|S\\�OT�e���i����#�%;��ISnc���k^�	� ��,��ذ�l�N���-Y9�h�=J;gy�1���w���.&��]���lʄI1�v��B�ؾ^��I��=oǐ	���駟F���q���	�t��y��G��ud��
?
\A;����+g�A3�����ĥƑ��ef״����HA��{{u�OO�x��'�w�0w��M�����/�:�e� ������W��qC�&�σ�]�_��8���B��v*KЩiL�s{s,�^�덱B��]�:���t|�TW;�IW/}$k9LTĜ3W�\�Daۖ�ۛ�23�Eii�e��X#�dj�������f�u*���G�g�^q��Ď��A�X����򙸞�w�v����3��3��m�}��]*Щsfn���3���Ϸ�oMb7t��w��R�<}dr�3S��=����2Qr�g��[6m�[�,�jxe�J���"S���]���X��2�K���u��u�]g-+��l�%��X��#����s~���ڡ�o�Ż�[�Y[{h�nئwp�k�e�{��z�&���AScސ��H),IUޜH��@IX�C�n�!u�*Q�0�'�d���|�Nt���{��L&v��R٭�=];�`Pq{�GS��&� ��풟��<���j�Zi�-�V����}Z�US�S'浻�������eA��>�~==]�u�$6��#�0e���i�5qX�N��%�E������� ��ɭ���&����:�t�{C�F������['nw�<r�r��M �k��e�x�����k|,��&����3&C�a�۵]\VP�vmD�[�ӝF$�ۛѶ��t6��Yj����]�������K��� ���I'���	(��R*�QX������k?x7w�}~�A'iIJ��q:'w>QŦ�ݱ#������@A�\s�QZ\��}iJ�y�����v+^�p�H.G���/9她/n�TZ��.>3aq�_��~{�S��A����;Z	�)Vpq�X7�넺�ew�ڡ�9#���#֚#��_�`^}�U�K�^=1y�4K�NA�O�~�u�X��˨�1�"r��^z	7�|3~�_8f���w�Z��1�>bu;c,�f���G�cq5C�^h_��uB^��F�=� [����	܉�2���cKR�%��$����5Ġ���/Dsqg$C(K�Tӓ���m�p�UW���D~2pH-�O���Im	���v��@�v�8TO0�vA���,G#�׵ݐ���SbJе�#vOq�S�]��ͥ��JJ�cS�·�Sd�$�t��5�a����(Z��h��R��NX]/����@[������~�ˎ�9���.���m"��uN�Y7eWn���gB��M�bM�;8��X>�F�,���pmW�1�x�y���Csޓ��n'�>������d�x��+�"<�ȗO?�C��ǞH�]�D���_=jjj0f̘�K@%�_,��m��g�5��p���>䄕��Ҹ��!A�nZ����'��e;��膃$�!� 8���s��R�S��}Q� w��8��w㳺= "9?a8���i(.JNq�݄2��d#e%EXx��0eTb���ث���� ���[�ƺu(..�4�ҏ�vjwj��zc,�v(�<j��kH�v���&���x�KWmQ~�p�B<��� 򗡇���G��� "�uꄙsfa��w�����O-Z�A���NK��=�����u�.���P�������=�wq���ᑞE���!r�[Bw� k�s(Vn��?���D�8�O!wĞ���U�%IŻ1�ɩ���DU���:�)1��7ʇ9��Y�D�Q�~�>ij5C��,�  ��IDATE�c%���t���m��M�!�k�( ���%����Jۣ��C����DD�o�s�ļv�IrmW���5b{@���ĵ]#:�����.��u>��.�vx�3�?ޟ����	�qe>֥�!]����ݞ�)���daz� ���y�S�lϛ>4�A�gbqm�۸=z�$�1#;�|�̵]�����i��j��1I�t�y	���|�Ï8�z��C�?�];w��/��ك+����z+z��v1{2Z�����ב���V�k'�����i'�L+Q��3��� 9�7�ٍY�Uxv-�EA����q��p��ӧ�^~6N��/�ݴA$���q���'n_�����g����"�`�F��[}"���+����� ���2��%�EL��b�Y������ uCK���b@���^�d��1_�k�̵���n��0�	GNA�� � �l���;~��{��W�ak+��㦛n�D�'NLj�'���xbvtK�1V�=�1_;�k�|��wqgӬ�ad�g�-d�#uD�^��a�uÑ���Q���������H	�@m�s'I��P�T�D����$��\��R`�DO:����J�KP=��� ���z�t��߰��������h-��#ҏ�o�u/�{S��TH�)��2=�k�6��N챴���J(�vm��]�j�H�k��/�����{�csmOf쎰�;f��� �C�I�.�9�gݔ�]+$��3��O�/̔��v��)����;�%'������,S�G�G���q��/�v�D]������v~"yq����o�~��O~�G��0>��#��ڵk��1���Z����U̞H߱����s�{�g{��9	+{>Y�n�������`��d���ɨ��)$�G)Qe%��l@U��knAA�l�~��M��[�2L?�6�<#j�-��s�=��-�AD|�2}4n���(%���~Z��pÃ/��0���f1�����g��v����@D0Nl?���5���4\���7�*�������ꆱ�cE7��MKU=1��R�ߺu�Q��A�Tv�)3��sEgAD��w@w����K�M�Xy�޽{q��W�[n���B�k���1�^bu;�n�W3�녎������a{�������=�=�
O���!�Bw"%̮-@s]�%6qSEE1&�ć����tI*��#r�%���ǻ�T;0����~�G���0i���;F�۳յ]�Ih�*}�u@�>��6&�=L9v����R���O������f=3��.
�����c2ܵݾ���2��ɢ�d���䷕�@�]��]����b���rkn���n�����7ͨm"W���M�umW��T��G�GD�R<�,?�k���L.ve���K��w��ƞVVV��}�,���X�or��7�.]��o�?��O�"`O��=�>�ik��&��s¯���k �C�V^.�,Y��c"{������d��� 	�YA��-X��A���z�����s0�`�L��貳p��Eh�Gn]+_�9��)I��c�'7/��/�D6RԾ�w��T?aXB�0�>��	"8}��@����D�VX�c��n(
��ڡW�PW+t_�)7[�^��$ې*��%Rglhh���۶m�1�M<�:�� "[�ܥǜ8o/{֮�_lܸ���x�(//�j1{�5����uR�>��Y����.����P�V����C]���Yvrg��ףW�A��H�?"$p'�NuyƮ�(��'�
�$�޽]��RD��4p�����3������˗[_�A��D�0b�(�9�0�QX�\��sn���1j��]����b�T��+1�ѵ��	����n@j�^�ve�힀�n��`
�A�������]���]d#���PHn�o��_sG�rw��o~�!�)��y��/����y�@\�1�VL\�@2]ەs�&�hm����g�a���?������~��1t�P|�_L��=}�2�_[_G�KZE^��ܽ\�CQ�U���;KV��mڱcz��[� � x��9W/£W��1���3u�@,��k$r'���	G`��N�����mg�u�X��H���-?�2�L�P?�=�<��δ�=h�m��B�l�%��5D^���������=�\�H�ks��MV-0���u���_o����?�LĠ�C@A��:�����xD~��o�w��.����@&�&Y��CG,�X&���y��puC��F�Kg���j��Ԋ۵uC� kF��x���Cw"����;�@�v�Ђ�I*�{�_�� @�J&UB�t͗H[�l�W\���&�CaQ!&9���h�	.l�V�v�V�_/m�Jb�B1E��d*�r+Ź��@�J�ib7����{�[�>���z+�k���pcu�[:�]��5�۩�kYo��ڕxwve��m�
kyvu�|��z��@����Sb�F;חt�"ޭ+ƙ�k�!F�x2=����$$�nK�k��I4�����I�C9~#��H���y8�<߯���=� ��TU��S��%�h���x#�܆��G2g�s�|�	�۷D~����Ϸ�<�0�F�t;+��G��qd�q�Ǣ������n���.�z������<�$��d������莃ts
A!��iκ�,�曨��=�<L��׋����=h��	���'L���Iж��-��Z�1��f#L�~�_���1:�~n_����9�I����~�8�s s,�Q����'n��V�0�9#�fX:�A�~�����'�����S����� � �����Cѥ��zeZ[�!�x���1r�H�~��I�󤻖�nc,��ϲ1�+n?��!m�PW;�	����>C����.$p'���>E�'�u(.�$�4.�k{t����T����&��xS�p``B�y��aÆ ���8��е[%75",n��3����Z y���\�j"���b��^��ٱ{�'ku�5�ve�FDx�!n׶�b�tm��'2As^���B;S�W���-�� ��Ϲv�]�֟(qn����Y�(U����	���τ���t��qr��#��}�����T߯f�����g��O2�c͞��x�����ԉ���J�y"�h��K�Qo�ќg4Ǯ��nu%�@|��7D�������97��m�sy��U8��YX��;��Ï@���͸��p�M7�gϞ)K@%Ý!��b�Y���ܰ��-p����{$��u����&�tɪ�s/q{$YU(��76����z�Oi�A� Be��F�v���ǵ�B���@��8�O���5��ذu���N��_?.)}����;�!�j܋l�����/��3�$��#K�#q;A�HQ�@?s���B�ݰ@��۽=h��5ȂS/�oO�x=u�D�x�p�w��/��}��(�T� ��0��'Oć+�Î�;@��^XSS�)S��]̞�ZbPc,C��o�E[�S7�����.���1ƒj�^�?����E��Q�����B�$p'�F��$7�x;���Cz%���T���T�k�_�*�O�%��ξ n��v��� �^}�`�Q�PT�������\��`RC������Q��$�?�صB�@m��99��V�]ۡ�k������	��i��p4��r����	��i=M[�-�Q�m���@
\۹�=ۄ?y�Fÿ_g����.�F���}�����u#��?��ǀ�������G��ˊ�՗�[�����#�"�>F�;�#��3�6����N���E8���ťK��g�"?ظq#���j,X��r���w�lrd0�O®u��Wwq�'��d�=Y%	��뢦��,�]{I�NA�lܶ�]�7<q�7ѽK�@��Wn�!^X�6+�ܯ��9l޾�	���_�1�<sfR�{j�G����b_�d#l}�K�9��'�Ͽ��?�y�.%I�s��=��������O�.�]���b����k�D�X�f��k9p ;��Dj8�GL����� � ::�7�I���O�n�Z�3x������?����O�=��X�K��SJ�5/����NB����v[�λ��5C/w������{0���]K5C"	܉�q\�����J�*T��IHRQ�T��y&���Ɠ�>�{�9,\�D�0b�!3~w�D��������3#?���L�k�����ʵ]��K,�YN���t[��mL����k��[�,�6�yU�z,�G�r�:�k��;�>V����.��z�/.��D�y9�K�����	��!��)��=�k�sN	Я���C�ε]�&�6�va>�yB#���qΝ�r�c4��ؿt�H�k�f�	ʹx]����ie�6<��cQUU��=L��<��_�=�܃��??�T2�b�#�mE�3���a�C��*9a庸�n,q�0�bHVqw��jmi�1�Z��j*�v�C��\�\��� Ad�6������^�������0�HyY1κ�D�	��y�bo�;�|���,ڲT��~������&$�ϊ5[�����e�H�����ϳ�`"[�.o��ܵ^[+�3��?D���� 2ژ���U7v:Oo��#��Yɘ/H̍��֨�uuu �v̌w(F�� ��%��τiSн����U� r��۷c�ܹ��{YYYRM��YK�Jc,�uC�Ktq�G��j���{[�������,6�{��o�� �;�$����a#��!}�TZ����$�d'1I$+I�7�d$��90\w�u�#.O`���'`Ȉ�´����\ۃ��|��ѩ��C+��,��*a�BaE�nǭ�+N��[Irm��h�S'׋r����ůlcu��}�79������v뮄�>'ӵ]�A\w�h|h�C��R��4B򤹶s���G��͵=2��i��9�v�db��=�~ma�N //[�ڮ�[6h�����c�?ǻ74yl5T�6�,ʷ����N>��c����j����D���rfΜ�Qz�	� ���VLV�� �uU�+����?a�9-Y���Ѓ{wlĈ��x;ݐ��̙4��kA������>�/?��;�}����ҴQx�@���q�_��G&.\c�+���߸����o��|ab��6�V�s��Ջ~��ϕ�݂�?���[����8@�w"C��݌杦�)�}��m�%��l���!{΋/x�,��Ea��CetD3�x��{��?�˗/���`��3Pݫ'� "W<|(:�����^���V�ϛo��;�?��O��'��*���ۖSRn�Pg�Ů��i�U ���5��\�Cj�PW/���5Ö�ݷ����9`"9�^@$涷�����Ib�un�=I�ﾐ�$��lIhu``��ܹD�S�~|������``q;|���l�c��ipm���Ԭc:]�MgN�?Y쫛�����"�u����Q�61�vW�.+�r"+��k�</�|���wm�9bhe_��=r#���P�Ӻ�b7�IB�n�����|�������;����y�Br�1e��k�t\�; �ṮBnmL�^�Nx�yB#"��qΝJ?�\�u���H�]�����D�^�+�@�6V?���>j>#Sl��{�޷__����o���Dn���ٰ�������I��=�>2�6�#��h��{;����N�#������j�U���Nu�����|EA��\�s�y�_�5K�ۑ��'��k��q"�t�T��.>SGL�������Ó�}�l�s���O��|���3~x?�a��e?�[��u�|���x�h޷�j�S�ƺu(..I�n(��,��Z��������uD/�-t��|��O<�ŋ��JJK0y�tTt�� ��uz��cN8���456��}��~�9'�pBZ����RUK��'��8���n�g�e�Y�Ю��hk�|�P~��6�؄��C�c�=$p'fXUa�IELR�
cb�@��������^I��lpcHgb�~�7bŊ r���v�L�m�n�f�Gpa{Gvm�I�âO5LU(���N=\�#B_^�_G5vu��r;�E���Y�&��z�4���c)��v��]L��:��*���<յܾ�h+m�f	��K�{�إ�#(q����׎ݧ����c^�8�-��\�+�k���^q"i��J�\o^�����˶��:�������
�})�qͶ6ܘ���cW����� �����m���.�ML�*++q����<��>�n�8[�l�n�dnc�a��ΐ�dT��+���$�,�v.i�'r�'�dG���<g���wafM���dA�����Gx���+�����r�����H?x߉���r,��l��;�v5��7�y�>؀l��g১N��a�!��&��a���xqŧ�M6��A�~%��&�lCKH?�s0a{��@�!�G|���YvJ���mRe�K�d�����`�� ��=�0t�p�AyE�ʮ8�s��җ�c�6��G]w�u<x0���:`�}�2_<m�5ƒ�^5C�5o��j�^5� �X��{�ctY>&c����D�VQ�����+A%&�
<W�JR�Ȕ�=]��K�,�D�SճG}���`܃����c�mg
��ԋEe!�!�e�Ipm�W���ڠb{��Ib_i��Wa��ۃ����x�����5�����*�1y�E,�qm��	sN�´d�����MSE�q���}��G��h����cwmO�G+$��3�M����ř�N�v#|�����;u���(ˇv�|um����v~ZiI)���x��g���/��m�z�-�~������c�T$���B�j_;B�J��b�k|�*,x��ŝOVَ]�mFyqo4��ʆ ��f��+-��?��� ����Y�[��/}D�QS��۷}>Pӫ]~��p_���Ys��M;����� ��
0q� ��3����t���;A$����\׀��OS,�;W;�j���=H�PW/t��<�l�K����k�.̛7MMM r�AC�`����]O�|A�Gq��ԣ�?�{�u�_�)��f��ݘ;w.n��6TTT$\��Uc,G[y�����B�Цs��ŝ��"�B�fشg���zD�Bw"!f,D��z�����ޮ^09I*��,&���Lґmn~mW�\i909�ACc��I�1�����"xF�sm��k{X�)k,U��{`�v�O,��ж�d�m�M֌j�4؞�1�z�v��sU�,�vA�m5zP�D�]�kcw&��sq\L�إ�Ҏݯ���L�6�vs��p0²�}�Ǫ{�����x#��<Q$��C�GX#m��<��ˀ��s�o|NL]��`�s���]��/����~0<�H�F_�憄X]ەx4�M��>��P٭;�||�u�L�.<� F��9s�dm2*�|��̑��~}�����b�����l'��]�-[���hii���6,Y�� ���W��K'��#s��'a���:�h87�/�v��VQ�\gdMO<x���SU�p_l=��Eؾ�c��t*�/N==+;�+�G�>��ӽS
wo t�X����X!�~�=��\3,p����X�xj���'c>�9�Fgu�?���Q���-{�� � ���q�������� �T��trl��/�8��_�k����c�]�����ۣ>����vq�j��QҼ	�%}��B�h�Bw"n����ʖ�8XTNJEN81����e��D�Tn�JLR���$U,m�:0̟?��� r�cFa��q�s���AT�\���M�� �����������K�mg>E������{	x�NW�����sm7x�4�^P���	���_�.��\N\ۅU7����J;e�s�`�Q�cMn�Y�Թ��q�?M�q���n��\wAc���wԘ<��A]�M�4�<�]��bqΝ�r�xLu���2���2�ڮóo�h�O�.ە�#�N��O�|�T�����އ��� r����a����R��e�#��*<�;wY�F���)9y�VV�#sa���n9��~#�T�bK92A����k�Z^���6���b���3p�/����	yo���CYIr���⾋�L��{��5��u�qoǸvb�oQaDp&2 ���8㊅ �D9�o+��ڒ�ޮ�٫n}�g�:��mfX��M�|�93	xꩧ@�6�x�|�4���AA�a���Ν��˯�1V��裏bԨQ��W����'��bi�1����n�����cuq���1����8c�-$p'�f�@���PR�{{d[Ĺ=SI�l��:���p�7bݺu r��>y"����!�p=���E�:���*:�y�`5�{���0Uq�:gx���k�(�Uc��ĺ��9�v}[�@V�Ƒ�$ͨ�@���c9�LM�d���q�N��0��Iqmw���&�ؕ��?v^!�Ǥ����ʉݧ���L�6��Ո����r_�]�ݾMi���p+���h['��E�@�GHν���~m��k�]�x�`��"q��(���nM ��k��:-���r;!��wذ��q����{；n��a���q�UW�O�����J*ś�J�X=X[�#�;��ǫ}�A9ae_˙N�J������{6��r�$� �s���-A���4�!}�,��7�}���"
��\p������|r�3{�p���SQZ�x�g���W�=��;N���I2&� �H�!�Ѵc�����¨�vYܮ�ٮ'1�E�{�t�a�fX~m�����{�����`ڱ3QU�AA��T�N���_�ĴD��4sÇǘ1c:DM0������ȝ�Y4�j��"w�nh=صc�vȋ�[�7�o���l��	܉�`C��7��h�qo�ەU|��+I�̾���4���F{��'-q������=��)@;�]��E-f�\ە4m�����3��*����rm��DZ���]����.�uն�A@����ۅv^�튃:\��?�2-ݮ�B�L��+�Y�)e����CP�!6�v7$�����ӵ�_(Ǐ�qmW:P���9�t}A;�r�34���t��!�h�+v������<�6	��kcҋ��i��~��sǝ������a��\p�1%�:��Bl}q�+ұ�;�	�D���n��udЋ�cuqo�ۂ1������AAѸ�/�BE�R�5k:*s&��OO���~	D��ѵ��W0��Z�_;n�����?إ�����ぃmh޷�Jsߩ� ��û�F���+Ƚ]��5�PLuC�A��{�,��a:��|uuu��k�?]{�2�+:c�qǠs�
A��{u̜3/�g)���@�&��l�ܹVݰ��2�z]�u�\3���a,���urg5Ķ6�����l="�X�V�cM�n��{�+!�;G�mž��R	纠�{&�
d7uhA]b�Oܞ�$U2O:2����Op뭷��]���t�г�����҈��֎\��刂u����]�)\۹?�4u9�ؕv��]�]ۍ��U�����d��]�7M�b��f�1Į�7�b��BL������N�4�X�n#n�,pm��,M�.Hm?���~���yا��� ��v;a���>1Y���<b�&��B��34�|�F,�������h�u�]x�j;uuPU���ɏ�{�ņ��A�&l��C=�f��ɨxWA������
7�we�sc'�l7ޑ���῜�]��PIRr	+[�>���� "�{�W�?�n�8q�HtT~s��X��3<���s����NEuebfL,�8��ɘ��9��Y������#/���ʶ]�Ի���i��H�#���~;JJJ���Q놼9�ƹ=S,�fh8�<��\7-�a*L���]w�����~J�X9L�U�s{Ii)� ��KeWs�l��ߥ�U�Dn�j�*K?w�EE��udc��my����� �ˮ�uDo'w��\��b4wf�5��P��F.��	܉���^���Q\\�8�j�vI����E�^I*х!�I*�rcH$���@�7ov��"7��f��.]���;���Nx����.���R[�PU��5�q���tI1�5�A��^^�/%v>6a�V�/�����9�05����>4m��x#�rx
���������z�,C#�v7��s��K}mr>�����)L3���v��?)&k����X5�۸�MwS ۽ɑ,�vML��¾i��ڮ�kjڨ󙦦/�k؇�ԗ��F��Epo���U!9��qo
Pۤµ=�	�$};nZ���������Ea�W�Ax�#,��#0`���AAخCtd��p���=���]k���>"w�I�vd�\��߂��]'n�]t"��]�8r@^��1DeA��O�N���%�y�c��v�� sm��Ÿ��3p�������Eq�g���[/�2���l�k ����4��;+)N�?��	d3l���۳�ݓ''�מ�|{���һ��#��?�q��ǀ�ܿq�C �x	���lG����ۣ�c��v�K?�3/n��{���H�Y9u��a<}i�H=�G�F}&r�^}�`���(*�QM� "(e��p����ŗ���- r�ŋ[�X'�|rR��T?�֒!����.�b�i���Bc,q�g��]qr�pqY�]ú"o �;3*�XC�B�0��ɩ/q����O�ŉ!LbI�lvc�4I��<{�=k�*�}�-X\R\����qڙ��sm���k�4]])��$�ڮk��̵ݔ��b�Ȋ����z�����nM�m���,�k;�Ů�7��r���K�C�3���ʾ�d�vg9�}��� b{�BM~P n_�Y�ޯ_ �\�=�o��R�����(�SW���a쬯���Y��^D�m�6̟?7�t�u��L6�,��69�-�dM��΍3�ލ��^��$��aC���wqw�T�=�yz܂����� ����NDM�J��~�FlmmDG�u�A�u��a�оxಳPեS\��n��Wp�e�D�Dl����?�N�6*��%�%w=�%�|�l���7���2}t�}}^߀��.���~���O,�Y��a`/rq��֝�8����n�sLm��{���$t�Ź��ꌱb�z�cu�a��~�!n���ˠ��1~�$�!� "6
�
q�13��+˰��u rV/5j����<����1���\�ЮF7�r놊1V�=�sHk�常kF~nڳ�kz��ۨ���11�O��m��U^"��M�Jp`��r\ $;I����1<���x�!r_�U�{�Ĵc��~`ǂ�ID��'SigJm�����'nk$�pm��r�vL����r})��ӽ\�S���_�I]OS�N�=bvm�׷�=�ߵn;G n�G~���^�k�kh"��E����+}i��z���k;�:�k��wy�����q��7����웩umc�m#)#�vq�Yv4��i��\Ѻ�	�vZ�yd(�bWVO�����6�4Sm��k{����ݿ4�Li�M�rک(++�KK_ �{���k�����|�C$�R���U�9�~����v9i����&�Z�)��]qq�$���}{�0��'�^C?� �c�|�g8�����o�sY|N�SGįΜ�k>"8��;u*���p_��⻞���|�J������gb��~	����8���sf䀽-����G��:B��{����_�g;�� ⥴(o�����#>s�>茱���b� ��l��������d ��Dnrȡc0zܡ � "~�o�I3�DIi)V}���c�Ν��k�?Ym8��]��e�1�Xӷk�|��K���������q;g�U�j����]?�j�Ņ=�J����D`���
������U�ƿ������r�C
&H#��@�QP��S���g�)>�PCB�"�  �#%��!���{��gvg洙��;{�?���3�9����s��N\��	K��T�4���O�>�k#U>�1lٲ^x�u 
��	㭡���pEO�"5bL�[����նjj����\u��<�N�wm7 ��U!E�����VS͚�#��7v�>vfitm��)�Gl{9Z[����J���]ە�ںK��R��:h��@�|��qb�?��n'�w_�{�;Iǵ�-��R�_I���vn�X�	⡖e���;�dM��o�d��|>Mݵ�;FW�x�|��q˷R%q{�\ۅE=�M�/n��}�|�XT��#�D�z�jx��X�paV���J�q�<�g�ȧ~#�����%r�l������g?G����.��Ka6m�ЊIh��� "��q'�q�_p�/NFiqr�����R<�n#�[�1���z�|��
e�wy�G�c~��A�����W��ǭ�8���r^�7�~y��QH<��&�ꆇ�/��Rٟ���Ӎ��ޅW�ߊ��݊�ތ�#�%�H�L��U����^���]3곟1Vq{��]g��Hg`����'[����/�Q����þ��AA����棢�o��D���k�����g��e�O0�r�C��}��X?`d~?'p��u�w��P5�bn�:q�`�I�ܻ:;q��"<@�X��Y>���!K$1��0�E1���qJn����O��7R�ȶН���Ӄ?��ؽ{7��c��)Xx��@C:7#�5M��dE�š�S�1De��!���O�k{̍ٔ���G˺yj��J�FخYO���Nщre��k�!����
�5�Ǘ��y��+��垟���Υ���޿��^�w�ܪ��q^���p���I���k��e���Η�
��:*/�8�m��d\��� [*K[?a��fjˆ��͖&�v+I*�y!��������ǉq�L5&����ǎ�ˁ��hH?ڑG��AU��]w�(,���q���[V#G�L��(Wb��920��}N���b�un�s?��he=���)���Hr�ˑA�Gһ�{q��^ܳ���&� ���>����}�8��x�:�.����{�X�T���A�(/-AMU��`>a���!����DZ�`��﮼w?��¿�>1k�e��r^�e���f����f�}/ZSX��W�����,��zz����]X��v�۰�Y������� �DUU����US,Nܮ�7���dq�W��W��o�YB����0_�}��Gq�]w�(<�>>�"L�1AA��}��FIi	ֽ�J\�>����kٲe���D+��X�'I����7����ɽ�3Ų�ͦ-V9$r���Dei�5�`�ƹ�n��f�Ht_�i��+nGLX�����ah�ґ.�믿�>�,��c�'f�����"��q��J��T]ۙ�Zjߢ ҍՉzUQ��d�fK�Sa��	_[�-��&�ij9�
�ڮI�|J�k;��)N�}=�=i��Rݳ�ڎ811Et�]�U1���-�w�B�Vl��|�����]�{�趑��̵�Y+}y\������8/���}�G�.��umO:.�^�{	�z�k�o����tt饗ZB�d��<�l�JG��|7]�n �sC��m�*�9��#ߣC��V��{d�س����Mt,�w>ޝע�t��bƄ� �H�;{�ƍ����4��x�7_??��>�y3��3?�r>�e�(+G ��*��xmJ��PUY�|/���Ŗ-Q�3AWw/���w����|��%�q��?�W��?܁u3[;@�}�]xw�nl�Q�rg'��a�]訇�oȞ�>�?��5��v{�g~����3��)S�fX^u`m!��F}.<��h�L�<	AAd�i��DYY���t?U`�������=�O����ڤ����?�,���K�3�r�<��#{�*�&w�g�~C��	ݻ���||���D�Cw"GN�GO]��+D������SQ���f�~��H�x,Be͚5��`����ܸq�`)@��V(c�Ce1���t�vU���k��)��G�:!�*浳L�k�$�t�5b{x�����
��ɔ����Z,K���x	��q�:j?�~w9-Y�v�����=CSW�u������J^����oۿ��{�u7�^���h�m��҇,w��B����u\rmw�SW��fj��c�8M^ʺG�Rum緛Z-7ͫ�Z!x�'�Tc���n�?z4L���$�>r��s��o��5���F�!
�x |0�=�ج6Fe��)����J���ЃZa��9�H�5�`�5Ԡ5G��92�D�asS�����������2���'��� ����[ǾG�S���'9�?�:^|g3��>�[�@���_�Ýxr�F�+�{���C:��/����+�P`���ۺfY����*A�M(+/�>��vI�^�هX��E��8�3�W(��E3,�Q���X6��G�L^Ab�ϬM�.��={@�;d�2�W� � 2�ĩSPRZ��|���
��;w��/����#S�X���1�"a��B�o�1��:�s�>�t�Œ)��Y�oh����L��Y���M��� 
�qVY4n��0J�^������UR㔟����@��F�t��ә�Wlkk+.��tuQ�D��\�g̊�L��ߜċLݵ��_�ӶjjSqmg�+u
�k;':W��b5�t[�-��&�i����Tѷ>��ԕ�Y�v؛Q��z�{\��X\��G��!�����z����b��}��H�rm��;���ә���f7���;�^M�\VԵ]��d̵=�(�J2<c��Ja��]z����k;԰��l���g̰D�ׯZM"��������2eJR�B��ؔ��h�t/c����]��.�C�UE�Zq��Ƚe�N�=o�� ���3�t����0{ʘ��g���9e9���Z�aOcN��-xs�N�#���w�_�Ԃ����ۛ��oEkG7� �e������v��]/rWG}���F{֚bA�Fd��͇~�t�h�-�܂�Da�\d=r9F����	� "[�N��G��=��WQH<��c���q�'��'���X��%�1�)�3<��Ϫ1��/F.r��t��Z�;3�ڊ����!�;��zѹ��奊���E��B�V��%r�5Xɓ����'�	�����A���꫱~�z�żE1�3}c�փ�����kD����WY:��r��sm��q4���J���R��V���]ۅ4�'#&&���|B�!��7ky	ĥ���4ݮ톽w{�]ُ�};]�u�y)�ȶk�������SW��fj��-=���f��F�������>X��]x#n��f�1�um��(w*��7�;�������6��Ι��ի���	�0hhh�^e��S��)G�l6\%3_����� ��&7T�C�V�C_�5�`��Ƞ9Ȇ�7h7Zͩj�ۨAA�	����߁G.>C�+^����`Ѭ���6�^6l݋��>�Հ|���מ{�Z0#-�=��&���ۭ}� "Y�Ֆ��a�5�,n/��s�X¨�na�ϰ8��]~6�3��"�}����������w}�pQ^Q��>y$�
� � �˨1������z�d>ZP\y�8������R؞l��L`c,��19c,n��1�_�!��yc����3f:��E.�	�	_�.FW�f�Qʧ�J7Ġ+t/�:0�6P�'���5���T#T����?��S���;A��}f�wb%"Xg�M�k;4b{��7k�������ea�.�Cܮ���-Ŧ�ڮ]ayC���)�Bq]۽�n8�
���.&�:�r)��[q���u{�uϪk���),gW]�������1Et�\ۥ��s��v���͗o�?��o��:!9����Z��Z���o�dEw��ȼk��y�u�J���#l��튰]:���(����RX�eh��q'M��g~��ttt�(�}�Y�q�8��Ss��Hl���3�}XkD|��� �2XS1/lw��9E��~��ū;�� ��w5��K���?;�j�L��?{0	��̿�݂�~w�ۑ��Q�[~qrR��:}�|�w���:��H�ie{��]�����>�"{�g�ɝ��B������C8����ܹ�:?yy��گ.�����絎H��
��$n'� �2l�p�z��#���D�CKK�e��r�JTT�����?�Krp����XŜ1V��+�_ا1��c�X��ϳ5�-T�(\H�N�r�.t���T��*a��"w�Aѱ��ӵݯ�J��S��r����'���*�V�v���,����Ҝ��Ⱥ���oTdaӆ�R~SCc��T�4�����zl[Kkdj��J�bB��8}��nR��O}�"��G��PY������V���ݝ]hkmX
Ww�j�~$C^>Jc]=�wMAЯ[V-�õ]�َlV��:������TѺ�v�W� 'ώX�}�޽H�7�����{��o��]󒅫]��8`���ڍ�ֽ�U��_�3L_��6\^M�MVC{EE�Z��e�x�H�y���k�N���J�'xd���ղ�q��C��=��9���ȿ���_����D���&�M�����m߲/<�^����,�!l���:��ް�"1�d~	��D8d�x��/[�1O����MUUn���}?���p��c͚5�?>fϞ�5a{>96��U≺(�o��*�F+~�Ag�A���;�Aލ�5^M-݋W1A6yy���s��	�&��g��VaOc��">w>�ι�>���!�5y.8�3?�&-�=F�v� �Ē��hil����>Ø�@��Ήܭ��?��9�~C�Y��/�Q}�:��e��o�������
X��]n�����\�h٬�}��Q=x0�R����a��~��}9�3s��l�9\��o���?��{ֶ���ތ���9��t�����6��|fϷ�kj��#���OjG��=_�\��{,��_~7�|3��o���	c�`��r���3����X�Q�Ց�������7dϗ�џ���b���xe�y*$p'<�:�m{7���<�Hk��5R	UE���/r�7X�7R�+v���F*�h�b�/��R����J[[n;�rU�-~����0�A֝��]���L��1M�R�:3q��ӼJE&]�wnݎa�FX�Ysm�����L�9]y�.�Zw� �v�BN>L���Ԍ1��i�Q�u��tm�Ҹ����6�������L��~�����nHu�%n���'�f�StVVHR��OV~_&0g7��ǎլS�������ob��k�w��vLS�Ѭ�]'�uҭ�[��Ü�x����K1ޮ�R}4y��G:lHdqE=��bt����}�_um��c�AĲ�󄜏��?wj���I�N�����7���s�㜼}�ĥ9�}�����x�"���A���� ?�Z�M}����>g	��$}�����ƆF�ܱ����, mRbq�.�5�_���Va~.��}t��g�v�����o�/�W_}5��N�l�,�3�D��tVJ��*^����M3����1�9��e7���,�8�m!w� "|\p������5ytB˕D�����_|D������͏��>�|�	�%�i��_�l����=�)�'"<G�����BW�?��3���F|v��ɣ��K��=ڳj��?+�Z����^z	w�}7*++֮$.S�|V6ۿX�D����ee�g�t�6�XS��������}�Y�֦f�ز��%�sU~G{������rA��}.�omi����93���[�}.޵)S474�쏶�\�ߤ��=9�?��|�η��o66���b���{,v��{,v�+c�T��ڵk-c�y��eM��Hl����}�����~C3j�U�:�������џYڔ�x��Y	�	OkE{��@%��{5R�SBcU�!}��O���*H^?�0��~�;-[�	�'i�7��2��}dq�)��R9^"Xi��|QZ�r+���uub���Ԋy�,�dK�*��v�zz�(�׏��\S�=b�)�X]OS����-�*G#X�t�B�(*��d@�|nx���3�P��M�ۻ�iĄ˦�&T�KS��q����)���M�:Hߝ���8��4���
W��ԗq�}YF.O�y'G�:I1^ǵ!�7����+��'l�XE ���+����F~�+u��XIܞ���;Ǝ�
�uy�j7��po��`��֝8����G���}C��(���z%o��c��[g���/���"��o��n�g�yfʍQ�uIHn~b�UjC���{.c������n���F+ޑ!�|�r�o����{)ƚ�Pl�@_�:d� "Yz����5���_}%�e�T��H���|���亍�w�%ng��_��/$n'"->��-(//wG{��Y4ǒ��,����Xq���Z��T��G��н��]t��7l[��FC�6�o���)�E]��O�m?��
���rnO]�h����	���~�����,���lD��!Æ�����wo߉��T���Ps��=�=سs�M������n�qֽC.��g/U�5�`T혜��K�۬�oǌ�'~�a���{,���=��ٔұ������^k���������J�h����u��^����ϱ���س��6�*��-c�g7��{!BwB˾�Jвw��HU�i�����8��C�'<�[>�	4�F�x�ݰ�μ�oߎK.�$go����-=�G�ߛ7N/rԔ�����cz�y��{���8�|U���������q�,���1q�R''v�����^r���bE�v��'N���5�)��[w�:��py�N���ݽ\�Mn�h�*І�{b��鬻#l�S+���� .�� v�:u�����A��&��þN+y�/����ߒw�1�'�;�,#u�v]4�=ͱk�I�~��Sm���q�D�^yi�K/����M(i�tm�.�[sm�>N��P���ر�cq�����/�\qr'�ɚ5k�`�|���llJ�|�gc�ΫїO��^�̱�k��>G�ss���!��*{�A�(�ڂe�F㉏��� �����51o���Dr�ߴ���;�yW#
L��_�]�t�DD�C�w������r�a�=�Ї���L�t��'p���+��>�Db�%�_�r%>���A��jv���ȝ � ����<��������BG[�D�D�x�w�j�*�s�9NZ>�zŦk~��X�6Ag�e����X��B�h�c{�r�X�1֘~f�5���
�Z��nBG3�@�5�7�`�ƅ�gx���Sh�JW#V��3%tg'o&n߳g��c��'NQ�^uo��To��5�v�d�_���2O['VS^RS'KY���g(�|>�P7*:��IYK��5+��n/�U�d %�v�X>&�Ӳ����CF�Ʀ-�6��r�tm�rU��vx-�y)@�}�-(�sI��7�2V�Cm�tǪF�ĵ�9Wh��������rXk���<U!�['�:qQ�!��Ju�
G�.��smwʉ�D���v��.Mү{<�v'�K=z�ɜ�W^"�0'	v}�uס��:m�M�#\6_==��bG��|f�~����8�n��F,ٽ���F����QZ4=�I� ��y�J�㮜/�m�i���n~��N��cC��������GGW
$n'"�9�u(��pD�}����E��%n��;��o(bpSz��tdZȞ��֣�>����� 
�ʪAX��$n'� �P5�ˏ>
O<�:�;@���n��2�:��CD���|Ay�|R��bi��B���1Vt�g�K�7dZV�+j�Պ�'��c��-�� �;�0��-��Q^^�
�97uhAۅ!��λ�;�ũ	�E�g���5�/���;{�1���ŋ0i�%=�`�9�͞k�Nڞ]�v��Jz"���>'v$��k�'nc+��k�!�%�|�Õ���\ۡIc�ޯ���eε]ZQ����+ʏe��kҴBr�r�K|��P��-(����ė�r�r��6�|����`<��N(��A^w���O�qm�뮋ќQ���~�E�I؍���]q��e�e��0�]���V[[�3�s6nX�D�ٰaV�^���NZ�\r�0�W?1Fj��~�~�jCUl�Aٍ��_�;Ϟ�#Cql�����)�xhcn�'b���D����<���`F�e�*�@�=^]|Ǔ�(2�iv-(H�ND��*3Pּ��!����Ms�
�~� �vm�!���Lp&�\��e��P7�޽�{;QT�Ï>U�� � "0�����'������.��"̞=Æ+���Ԍ�T݁�o��1z�2�*�:��L��џ9c����(-�EO� j ���P�V^���R��ʫ�J��^$4V��z9/$�ޮ�a#U�n[�nŕW^	�0�w�BL�!K튋�/T�ȝk{t�ZMS�������㺶�����i��XE�K׊�ݥ�*j]��b���zF�ޮ�J��8G-ĩ�kY|*q�:�{�J�a��Y\Z/��=�I�ߚP��먩;�]ݹ�$�[�K�\��U���+˽N�|��a'���.�\۵Ǌ�w����Wٯ5��]���ï�]v<����
)����IQH��ɣ�@�y���������4�������gƵ]9���89�HԵ]�&���ƍÂ���g�AgG'�ps뭷Zn�-�HcP���.���CN#,�]��*�y.d���	�9n�#�0�"iF�VT��GٸA!�/O��������F�$-�]8�ҿᡗ��@���Ad�����n��X�7��;,Ҍ���%�<ڳ�g�?���k`����^q�زe��SQY��>�Ճ� � �p��߇}$^x����?����;�<'-�����w�E�O<c,]ߡ�o���
��Xa�g�!?��-t���Ċ��H�B������hi��1k�
4̠�&M��P���4�ܔX#�.-�������@�&n���L!-�`�9Ƌ��,UѦc�C����f��V=]�!���\Oq�R��>A��'o��]+nW�6�sm���n3��{`�vy=bqZ!�	�0޳�r mw������|1�:De����]KC�����v׋�uu��@��v��܏!�4�i�u҈˕�b���դi��r���\ە��p�7u9��I�lJbwnI��ג�r�r9��S*G�Cp�vC>W��v���k|<AzPѺ��K����v^���4���n�Yumא	�vS7�f0N��Xu�U���^Xc�e�]�U�Va��#1�� ��l�O���{�Fvc���rC�W�#Ck�*
�P�>wu��*�� � B�3olJ(���xw�n|�wb��z$H�ND&Z��4}y.����"w��]5���;��GQZ��ӥ�k�������?����O��Cj@AD8\S�IS�ཷ�AwW�ps�wbɒ%X�tiF�s-l�W?Nu�!p���}�|��)c1��~[�����)�bYi%(i�F�X	�	�q؍{�A{� �E���=��X����v&8O2B�x��ٍ�����#�<"��p� nw�D�*�g�ε=&DU��
��yJ��zK�&���IF5�d>]��<�SsrfY(�m�vE��H��89M��f[���k��fH�خ���%j�����u��i�>�Vwa;p�r���A���>ism�21M�y�A96L��Rum׊����~KS�����c���C����+�,���.�7>�9�xM�8'&���n7ϼM5&��Jݳ��nh��0#}��n���S&��3���W^�����w���7ވ��:K� ��Ʀ�6f	gc'F���=ܠ鸷��EG���{�v�A;�Dh��6V�i��'������ � ��6���vf/-)�s�?���s`݋�������A�d��^t�����\�3�?�+l/*�o���H�_ȋ�S�ӑo}���֋�D�)�(���k�AA�ƺ��O=�(c��G�r�Jx���1V���ҙWN���?�zO��P�7����r�����E���Xv��m�%cu��������
��0���&TT$6Ġ3��5���D]2�H��F�d��*k��ݸ����E�?��= 3f��T���k���#�e�]�����Uŭ\���b{���x� W/KzF؊f�L2���+�Պ���W���o�m�vC�#�eҵ][^��k�sw�<�����vO��'������:�i���C�ε]�&����u򪳝&���Q���~����2�_���/Ɗ��>�c�P�Ѽ��)e�v�r�1푷t�s�RqmOPoh..��	�,4?�u��ƥ۵]7u�}��3Nǟ�����fn��&ˑa޼yy#<ϖ�]l�RNx�=�t�����z�8�����E�؝�t��1w���n�:bp�� � �P��/�:�1���ƿ�݂���ćD���i�)��٘g_�7���h<��C|������ ��3�����3,��P�Ct�	��7ƲӴ}�|?!�=��ܤ�/}���O�~��p˖- �MYY;�H:AAC��ң����z=��e�B�>��իq�9�8i���:?k�XV�~�g���;T�M����+�+�����mS,���Mh�F�X	�	�q�t��C�Z�R�Hh�*�3uapO��T�\��ǫS���a;w�n�k���X�]�P�傊���v^�TH.�n+}ե�� ѻf�.�N��m��(N�N��m�_G~�N�˭��zʢ]N�,e���x�m�nw?a����k�����B������lx1-{��B�|�߶u��A�EN]���Hu���3���$]ۅ�\�XT�|�
��.}�v>��])KSv"������Y�sm��A�;/4yl��b���!��m���k��@0��',mǩ�]��m�;0�/i��3��"��3f�?��_�a��A��q�%�XV����,���wi�V�Fl�5ܠ����1D�)�#ϓ�1W��"}C/r���d4oCu��vӐ�AD������j�߹�^|��>+e�ۍ��v����`B�E�&8����6⫿�]��b-A����}�CB���1���@ߡ�)����?/�}�٘��3���{�n�$��8���AQ�9K�<O=���+��v�mX�l:� ��0��X��D�o��w�>�s/B��X�����w�s�������� �;aq���65&��n-�5R�\	ۡ;щT�6Rś�o�P��?��x��@��I�L��E��A��1^d\�a�;5ǜ-����<E�nih���=Ĳ|^��;�IU���vN�n��B��M��qZ�v)����&�|�����ٹu�_e_T�3zlh�$-���\']�)I�����>�����)c���;���%��b����/�xݺ�ǉz�Y���9E��[�����Qʇv�@��bz��O��UwUH�َ��-��ڮM�^�
˵]'��s��8�?���o�DxY�~=֮]�o~��ƞ\7,%���26q��F-��
���*Sh����|�L�Rc��p�ݥƪ�'��!	� ����G���^������-8���h���_�Z������^�@��7��ݎN���V����%c��"Y�n����N7�����4�J&�\�oii���^j�N���/Y�#F�AA�ɈQ#���C��O[}D8a��]t���zTW����?�=c,Q�K֐��X�)V��H/p�0�b�@���
�㍽����:18�TE\#U�\���xRmJf�\ͯ�����p3�f0.Y�|�aTo�׵�O��!���&�Kл��BaE�n�[�4��J��L�T��@�rrf)}�^ +ocu��	�!��+ǀ��Ų��-�v�U2�P����h+1N�޵]\�%��y	U���F �"J=eq���,\2�ڮ�G�� t�'���S'S�K��������u��Bs������=���8q�N���M���_�v�N	���'4%�OqmWҌl������ �������DxY�f�.]�ٳgn�����D���rc��A�������"O��wc�VT��G[��p� � ���RQV��"�Z;�?��⢤���׏A]s{�;����f|��w��� ���|���h���T�c��j��=kj'p��<�����L���W^y%6n�"��}x��%3�AA6��cᡋ��g���&��lذ���;�����Z��	c,y~\c,��t�c1�����y���w�
Y���7�r��&������X<�-���8.n#U��*��ʷqJn���8��H��<�=��������A���c�`��I�}�(���9Ƌ��n�j='6S��U��q�A��:�3'���5\OjEܞ�k;�tS#Xw�)�]%q}]YA��pc��Nŵ�]uw���^H˵k�U��.ޏ�u�^s��G+l���따k;�oͱar_��BSGSS~����o���I�g�U�kFr���cM�;�E��=�d�e��<�h�9�+ŉ)���#o��ν���]�+yk��� "xum���C�8.ۮ�"�[qԑ�����>"�tvv��/�5�\���2+-^�O&�g�1K�?O��nP�ˍUѡ�}�u.��'��� �PAw�;Mm]��G'��,��v;򧳎���Mx��(D�z��[���� �L���{>v���
}�v?bQ���еܔ���L��|9��^��w�"܌?�LAA�IS�������2��r��7cٲe�;wn���0c���ÐF~��2�*v�
���c,��=f�U,c�l#c����ס3Q�v������C�Bwم���J<A�T�\;+d"� �T�=���^�e��X�|��%���7<�]�%ѩ��*��h����D\�U��	5S/����S�����j���[2��.�O�n��(˺	��,�k��jƅ��Hٵ]~K�g�:vE�}���Y��R�ĵ]WwC��Oݝd9��\+nW�+��>1�F2=b���v��5�����oH�k;���q��
�w���_�#l���C��h�Τk�����\U��W�ȼk�P3vĩ�]�R�Zk��D�Еk���m"�殯��L�m'���c>�)tv��ǟN֭[���'�|r���1K��3��*HW���+w^�n���5V�V9HA����bTU����׷�^z'�����I<�<����J"�~���ذu/
�����6����A�������k���X�;���n��eO�����퉎��3���u_����с�+WZ��Dx����}K�{A� � 
�i��DWg�~��G�+dzzz,c�իW����JK�+���cI��ee#Ic����ݚ�ѕ�����
�pO(AkSC ��"n�x]#�ށ�cx��❴��%�L��Lv��Hu�WP#U��<K�8�q��#������]���Sqm���=���!=�j9�n�b��vmc^#-���++h9�|��2G���z���(���R�'�ڮ�]#����ѻ*u��S�{h~7M=u�U��Ǹ��NH�@�c&]����Y��Ԥ%�ڮ�C�./h�Kε=&$�~�x�������R��si��)�A�������}�hlh��^>�����.]��'�B؞�2�Jb�i���<���L�o�*�L��+b�T��U:��&| � "d��c`��1����ڇ^)8q�́��%��;0����~�����R���C�+q[d�������ЊB�����_�B�v� 2JM����͊s{P������-&����/t�3�E���>B��7�x#�}�]�e���a��fa�R�A�@d���������p�~�z�y�8��R����|.�u��E��+��G~�`1a{��	ڣ�����hَ�����8�	�8��Б�{{�F�D\Dn�|�T2�dc�ڵk��*ĔW�c�'�@EeE�Xӄ�����ѩ��*�o[۪���T����TU����.
x�:z�]��b�?�sm�qL�+kF'\Y�OS�1���.�)u����k�f����[���-Kֵ=u��&�����;�V���1�Ƹ�t�!�/K��Z~|�v8y��v�Ÿ+���>�y�C��mq��[D�������ܥ����#l��+�j�s�\w��HU�_�Fx���]Y�D����.ot�?q�u,l��~q�l��]�ߓŴ�qn�j\T�{�i����|��Fᣱ��V���矯m�	[�S2��k�29�{"�U��]h�*r����|����^5o��*� �����|�q�A3����O�1���=�k���es��`���9�z���S1e찄��8z(n������n�(���{p������Ad�#&�讋���7�>���Xv����v��]���dK��}���n��&�e��i�oށ � b`3�������?N�1�a��)S��0]&W��ɩP,
7�3�|�?�}���Ϧ��9���XEE�M�lc�#&�1V�!�� f��R�46�<%�v��a�I�*?7��$t�����*İc���Q]]�g4�k�c"KU{(ƈ�T)6�k��CJ�햴j�ᬧ�W-'�k�R!hE��t[�.�BJO̵]���5qirm�Y����|����-FYAF�,ʽ>`h���d�j�f�������|�#���\ۍ� �?��j�Ǹ��NH�;���:i��/n�wm����(P�v'��Ƹu��]�#n����Sz��=��Jޚ8;6��rm7�8S�(����f�!V�k�5�V^^�o|�t���Oؽk7�����bŊ�TOk���^BwY�n7^ɍU	��G����:qsq'4� �PP\d��� ����������t����s��ĄM�=h|�������W_���D9`Z-V��E�����/�/�m�ی�Ͽ�� ��$̽��qK��Ŏ1V�3��ϾCO���gܽ]G����W]u�5�3Nj'����� � ��`��ֽ��;A����6\~��袋�}m�"l�d�d<c,Y���=S�c%���&2�
7$p�L*�k���s`���{;�He(U^0�*��r��#��T��r�J����l�?��e>r�o�i��&�dq�.9�Ft*���*Tw�̸���Yqm�V�R_)�]N�,����n7���c8�ʂ|�ZN��J����v�����0�:����'C���o�������'Pwq'��;�꤫���v�D��G�n]ۥ4�~X2�ڮ��-����������-L���@��v���$���/����	๪�/�CxT��	�v�\��k��K��:�v�hs��z�Ĕ��Y)	����TUU���9�^t1��@�v,���bȐ!����g�1˿��m��j����CT����{o/�^B�UD�2a�JK�-���&c��J�o��w<��{��Yh|������;��9h��Ə����]��r�g���,�eZ:�0��Њ/��F�����h�Ą�?r�t�����\q��o�/�}� rCԽ���	��q�X��X�s�"l<���M��ԇx���駟N�����-��}� � ��-z�G���"|<��x��q�1�d]�o~>c9#?'`���yW��)VPw���rq'c��B�ʂ�%hi�Gyy�{p�xQܞ�{���
j���X�T��Y&Wn��w�y��d�!�0v|�oLT�/����+�NI �um�3Ј[�<�Y	V//��Rw>�C�.�Vź��v!��v�صH�k��D]��
*�&��.�"Ĺ�u7��w��K���ڮ�ŭ;��h���Hڷqm�z	@�N��vy��5�cZSǴ���u
(���F���oajb��,�1���+uJµ]WwAH�QwUH��1�KjLJ��X/q{�8�е�[�ƙ)�A���k�s/96�:�L\v����	"\l޼k֬�w��]�F�|l�J�2�J���X���[�^�U�96��P�:#���I���XE�5O���>��
;��d6~z�
L�.�;b�4���[��f���?s���S��o�l���C��-3zX5���C^��m��76�v������ϗ,�z���'{A��;�B��Q׌�2&�����AD����{���X)����Q� v7%�ޞ���t�w�^�^�D8�\m��\RJ�� � DJ�J��#�����D�`��W\q-Zd��曉U�c%��n�)r�Xd�^�	j�2��%��0�:���*�{�,b��C/J��*_�t$�gCCV�Z"��7� L����|�"'#K<���p���Br>Nl�5�vM�Z�n�2�xq�R'U�kIU�FH�k�4/��d��٭WC%.��	q�&.ݮ�8�����O��ƚ��i��I�k����u���쥮ʊA�T�A�(��|��wf��?R�^vC�3"����n���F�����r�ܴ���a]/���"��RkYLyd~wOtxy�sd>�E�|K�����:��Յ����Չ�Ύ��N+N�}ma����7Y�vΑ\�7����k����|9v�&F�p\�5��@���k�V��#X�]�]ۣ��_�L��k~�X}D!�u:�
у
�����Ԏ�ӿ�-\u���y���z+V�X�9s�d�a)O�,��XŻ1��X%���t/�;���k�*nۆ��q���n#�0��+��y�w�����G!QY�c���N<�&���Ԏ�{~{��˛�~�.�AO��('9#�T��e��a�ܓGUEb�팦���bdGW��f~�Y��&���'-���͸��u 2Ϥ1CqǯN%w�	�O�\������"��=�v�з�Px�4�I%�����o�5�\�]��8����C�\���
1�`״ʊ����#�GG�g�[��/Bww7����Y�_�kA�GEe%�F���#��۶m�7܀s�9�IK�p*���d�e��ߓqq�ͱlc��'�$c��A�ȬQ%h��k5R�B ~�AU����ۓso�?a����=�XW_}5v��	"|L�1���㷟�"�Ћ���/:�c��G�v[L�&�bY7O��Z���]+��딄k�����Ă�����tû��]��J�ڵ=v\xם�QL%��++/ð�!�\��j+�4#7��0��g����hmnA��]hkk�&&�ʦM��أ�"U�5���
���<�G��¬�k���(vg"��Hݙ��n��o�p�&I�k;�����	ۥ�D\��"yE%m��q>�����B�8uW ��1N�Fx���n��d˵=V��T�q=���j���3�A���k�{��`�ҦϘ��N=���D�`��]v����:#�vdϖ^D�:ȍU@��*/w������ϭ����n;2tuva��"<�)��� �@iI1�;�8�ww��u���`�	��;�Ì	#����U?:KϾ
Da�?�L�ńQC|�>�p���i��ooC}s;�ʲ�Zn����:t����/��-8��	-�ne�x�g�������g�ԅl�g��5?>��� ����$�ִM�;}��bw/c,�_���h>C���X�\���ه�5��^����7���8�kj@D�(�\�BU� TE�V�~���43f?w�6����L�^QQ��.�0��?��\��B���	��2����c��e$���2tv1s��h��i����s�$3
imo��cvt��=���j���#�ӏ<F�X!���o����Ν�R�\������3��xc,��P��{�������cՂL��	� �մ���k��pq����f�wg�wo��d��6P%�Ho~>�5x���q�=��#ǌƼ�j��+�hĘ�5�1ѐ��\�*"��H�õ]�rBaW��;* ��cˈu��s�Z��<ëRV���p���u��f-�O�n���+��,ȧ��,8+$9����3���nW3���\���q�=���bjנ�(Byi9fΜi��Ʀ��>t��[C�n��c455��"�_KK�5���#F�@EI)fN��\���u�5p�76���YݟyA��ES��.��7{��=�@<Z��#�+Y���N�tm�
�u��g���+���=�v�pm��P�Ο������K�̵�>#��;�#M#n75q��=����>"\���+���{q�����)��v��J����� .�ȝwq�����]l�������B�1
}q��"l����Ɵ~_�Ƚ��?<�0�}��(�ܳ�9y�s��үn½��_qŰ�g����N��-ؼ�ac�Ա���'&��ۼ��n� ���ꆇ���??�Ȅ�-�l�?��%|�gk���p����G�ˑ}>�h� q��3��:��O2�]߃rf���z��}�Ŏ{{q���a�3��M*�b|��2�����^��'�S�`��������KDn`��Æ[��!CPlĞ�b�����1�x;Z�6`g�KH��9�����[H'���̱l���cƣzpuԔ��D`�^L�2v��5ԣ�'���D!2j�h,\�/=��p�^,Z�r%V�Ze����vI�a�&���X�wC2�R��l���X1s,f��tr1�(mlD�0&)Fk��ȉ�<���o��M�Нo������*z��n�bd�q)[�$2�=D0�D܁���=$�|���˘&<.�<�8Tc�1Q�~?��n������n�K������H��׈�=��Z!��E�(W��ӵ]���%.�k�X�O�\�_\��������u���/�_S��p�;�k;k|*��Q#��'�fo_�f�DC}=6���%`���F$���������%�c磡C�bܸq�6aJJ��@q$�Mm-���CgW�}�R���>+o�[�B�ߵ�s���]Zέ��c���iA��k���������v�sH���wu���r�6�+���83`�U�4��L�v7�[.�=���Ϣ�����e�5T-[��F�J�q�{~�]�SYƻn��"`c����m����,w�"K�9h5RIn����V,�P��P�QxT���柟���x7|�]����N���>3'�Jx���R�����8�o����Z]�;m���������>؎�0�v8n��)<�<�对�y"���Y��w������p���2��S����=M�w�
����8���ȝ�<���?�A��b�De�N���(#>{	�3���L�&�YT&_D�:�чx�-����>��;�&N A��]�ƌ�qc�b�0vl-F�n5�3{�޽عy+�m|+�:Vg�_��齵Cf����&��������"�Vl߹���"�L�g
Z"��;o���"�[��2�=���.\�7?��X:w^��cY.��X�n�1����=��E�ZD( �� �Q]託��i���\a{L�^\H�.7P�����T�¼��.r����p�޼[z�(/;(�x�Rum����
R�X�|;w�Z�-4VoNLmy~by.ݳ��v�Ny��.J�=ʉ�P�\�c[͐����T�e��C�>|E��+���*�[���j��N�H�غe�Y�&����������a���GCC�5�_��Ig���c�b�ĉ�0����7[�z�������h�
��O�.�=b�|c%�^B	����Y'.-��h���IU��q�ܒ��ӵ�TӴ���q�X/1�����vII^�C�-+%�z��vq�����I۝5 ���S�w�l��1��'��t�M8�s�������BjJ.�B�{���<��G��C:��In��%g��i(�)-)��sO�D��?�� ������g%$H�).Jn9"�a�'��V������~�V��~�5�{�����ב�Ԏ�;��Ը�^l�݈���NMk��2v7��s��F�
ۇ����4�v"Ӭ۰�=}I����Y��g쥦�,Q�1q�P����X�oj"���}���
� �ǲI��ljGyy�22���4�ﰘspWM�\q����k�����(�0�J��t�u�V�́S��}��A�ePe��P>nl-J"�(�oX��1�{o��?�[7o���L���^/MUF�]mm-�?E�%(++Eqi	v�ك�w���Ad����֖Vl�h�p�z�j~��3fL����3�e1ƲRݨ���(rf�Ż�k��Z��x�h<��D8 �� bTU��[R�  ���������;1�'!���
��*�|i�Je� y2��뮻���!��ߋ�/Cu�`!�4�{3���bL1������0X��U)+Kg˵�� �R����S{
۵Bx��g�@��m���-n�r�ܟѣ/a��g4ή�>�~wM1J��8Cg�7CSW�{P������1���Zמ��>455Zo*3q6�^؍>s|g�p�ԩ�>a2��ˬ����	{,������$�x��h�&/C���'^�r���浜WݵB�81N�FP���.	�}�؅��]�c��C�]�_#��=Z��\ot�ڄ�q�F�n��E�H {Y��o���~�A����G}4�̙S���t7V�.���i��<���,������Bf?����Á�#��j�"
&r���/��7?f��3̵������G��Os�;���چm8�w��_�W�̄�l�5y�_�/������A��}Ҙ�_���-��sw�y��wq�ooÍ?�rܗ#x�k"˰���<�����s�}X���~��y������Ww>ܞ?�&����c1��"�~��Q<��C�=F��Fgq��_�3�E�Zc��"!�˹�S��Y�yI:�~�N���l�&Sv:���k�J�p1r�h�_L#�D�6d(��2U���vv�hjl¶�[��Hw� �Pl�ƍ�dî�#G�Ĥ����}c�Z�[��Mhj�kAd������V���"<���c�ڵ8��s���8�g���3�3�]��>C&rgϙ�VaL�ޗ�1����Hmj@�� ������E��p�1��#���m��D�]i�R���L&����/�믿�r$���E1z��{V]�!��|k��Țk��'���=��)nW�ԉ]ˉΕ��X{%��1��!|��Tˉ�P\�v��ԕkz���q��C��������׵(--��1��)����ض�?��ըB䆶�6���[��`�x���iӬ�{J����Չ�;w����m��!n���1�.)�v���y�vM��(i9G�-	��k���ō���~��m��s���|S����jjj𭳾�?]xzzz@����^\q����+���vTHG#S���l������9��Sq���}V�V��s,���s�Qь�1𜙈�s4��iGb��1��GWw~��Q3��r�������ܖy�e"w<��&|�¿���91����-�A���3.�+6�ʯ�m�v&�N���ڄ��z�?ϼ�N��Z���S0�&�5���&��g\t���I���(-)��g���}Ƅ�x���y��ͱ�?{	��_;_��´�w�O��{�A�c��R�67����w�g/c,�+�|'��U�v�ȝ�?�bpS���&����^x>� �pQ=��,_f��A��oj�hL�0e�l��$����FKK����ߏݻw[����1y�d̛5Ǻ\���Y.�o�lj�����F{[�p��m�1�QG�y����a{`c,+I���Wߡ�gȄ{��X-��8p������� 	��ˋ���qtH�X�0a{��Jpp/vE���:��l����y!�e����۸뮻@��}���}fNw���x�ε]�_�!�+������8Y���S{
۵Bx�7���e�v7NW'���{�֥rM9ΐϴ��a�9��Hi�zj7CSW�# �kl���L7�G�B_o:�;��G���^!W�<�5f�رÚl�{��30a�8k��֎��pi�n|�@<��<m>�qK3�)O:��'N�nJi^������	�|�4��:�v�|I�Htn�I��M���N��EȞ	�v�t��c�&�פy��}�õ]}1�Ą��_����Dxx饗��C�3��LV��3�rRuq���ƪ�.{��#{��s\����ݘ1b:6��� :�z�����d��i�����X��ﭼ�7�B>p؁���~�F��媿=��y�����?��5JA<�;���[��<��L�����TL��s;��+�zDƺ�q�O����=�G?�w�ll�݈���/d�[�������}�r\}������uaoS�;����k�=s��MK~l�o{Ad��Euh�̰����,��H0ƒ'�(�C��-ˉ�4�ϣ�ϩ���2�gfzp��W�H0d���a�G���A�FyY9Ə�q��X�X����K���Kd���
�z�}�f��"�ע�Y#�E�%v����M��L�"%**+#����?AOw7�p�4�~����Bii�����v�vq���=�7S7ƚY�D�X!����'����q��*n�AQ@`;0�N
����J��bv��Jm��O�2����]Ԙ�#=���1�j1g�\�sb��O�l'��.d����ѵ=eq�R�]ۥ��]�iyC�fo61�D�\�c���乢h�Ȣk��um�����q�P=�
��ￏu/�L����w�^k�1bWѵ�4e2�뱧�N:5qCݿqm7�Ӈ�>8���Svm�-'��n9G�-	����n��g'm{�ܥMJ N���S�.��
��X_a;(nc�v�������?��c�{����,]�C�Q��KcU���2^�U�}��X�!r��w��y�b�^ϲΰ���}��6l��Nf"�����m�<�f�OK~��3�\�M��ȫ�XpOcn�}fM����G43�����Ǳ��W@>���>�q�]��/���D��E��y ��6#W0�/;�G�N)&�߲;�\��[��3�]�;��+�Ĥс�;�K�����	���ܻz���ǡ�8ywW����?=r�g��W�ӛ$+����,�+�Ғ��v� "��7�Mu�{��G�na�X^�v�y/]��:�Я�h���_�5�p���Ň/�F=%"q�14q�L�0��?lokǦ�>�3o�"�a�[�l�&���;̜���
�E�m�lh�T�M��!X��<��S��/���5"ӱ��p]���5Ʋ�⻸g�K�3l�ߍ�#��:z�8�!�� �,�+�l�K7R9U����w`��ۡi��5P�d۽=[Bwy�?��<�<9�����j�lIT��%��ϵ]C���r�JYYZ�Rng�>ub�1�%5�q��qm�S{
�5�
�vSZg'.K����)���Ҝ����Ԥi�G��Ѳ���j�?`��i۰����
���A.uuuسg�Ր���oc���<~J�ˬ�hˎ����Cs>���J�	%��D������g3n �<�+�N���qm�+��<h�z�ӥ��{�&TV]o݅@sΆk{B"�hj�8�4q��ݵ/
8�4qb�џ��oێ�^&_Xغu+n��f�y晁�����;'j�n��4X��Ѿ~ΑA�Pe5RI�ڍV-u;0a�4lm��*"�hh��q?�}��8�Ғgq��ӎY�/-? 7?�*n{t�۲���(���[��_��B,�*|NA	��o�'�>��I�Ł�C/�����]���D��>}����E\�����ډl�d����/[��T`�m��ч���-8��kq�/O����/���-{���3/����7��э�?:�e�w�����N�4���!���p���3����/�80my��Χ�[A�gVu3�{K���8}�n�a���^\�������ޮ#��0#�5k֐x)d�p>Fצgd�(0S���Lǐ��V���m���O�� ���A�{ ��a��sQSS���^��4����t���c������A���l�2:4+}��#l����z"]�aƍ��>C��ԥ����$p ,�T���nk(���TE������X��ޮ{�P����L�	���l�իW�%�%8��PZV�-��E�"���p]��r���)nWꔠk�RM�� ���[e)"xC��w��\��;+~�;�[w�K��}���DEy��3�e������o��Gz��(l��w�yǚ#G�Ĭٳ1�f0����������)�!��rm��Q�Ը|sm��\SVPq�sz��54�X?ز �I	�)�u�|�(n����15�X�%lW��ow3�v�D���W�c�v�ܾD8`�O}�S�g�}�.8�T#S���j�\ܹgC��J��VVC�Ƒ!޳�3���ЋEû����B�����߹�oX��6��kG�ƣ���{�51:#尉��Ճ��^'�	-m<sn�XSU���g�r���(�����Ҵ�[���߾�xr�F&6>��wc5sr�v̈́�?8q���!xw��k��G�𷮹�z��-��7�w�%2�E�wv����>��Ӄ"ϸL�<xP����1�>�R��a��J��ĄQCQ;���ʻ�w�'�>"y�y�?�7��D,�;-�2��U?<��l�m؎L�^���ooÚ�|9e7�Ic����)kjl���V4D�6F�����ȹ����{{���Սp����~��+�JQ��F��aՕ�>>"���Ze��n}�����>S����n��+<D����N_�6V�+�g��l_%�̪U���2��g�>S1���� 
v=_;�m�X��Ptuv������������Gcc#���K��Cuu5�O��A3�QVV�{va���8� ����~hjh��M�A���;w��o����='-_D���+�c�ֺ�W3ۛ{A�/ԫ[�������� �V�T\CbPq` <��*�l9&�;�D�a������0��=G��e�v��>�?.��>��Ғ��ݬ3��~Y��0R�z�<9�����}/!I=���ڮ[1�����-�.���cWX+l�f����Ų]]]�uo�"L�.)����::�#S��eu56Li�����푸��N456i�}ut���<�{��(U���*tF���Ǟ@kk�5��y�Ɖ\��;;ߖ���|&�@+����C���lڴ������g���Q��"`��=���҈�5�� ^ �9��ݳW���uo*)a�s��C\���aod}�[N��rP�4U�h؝v��:�w��W��kU��8I��mؽs�&;CyK�v�ruҍݡƱ���n�����P��f��u�׋���m�mعc��=M��Rj�m|����>r~�weu��=�ݩ���|�����.�����D�r_���*���K�.:2���~ˑ�s���o�'����n�VLEc'u���u��7^�`�%�7�&��W��X#"�l��{[q��wa{�zd|�]|뢻��G'�3�0��i���;{,A?{	�H�-O����_�q���;G���/���^�����o|��~��6�^�HC�+�)_�9"�,ށ���`~��;����8�vow>C��gR��t���O:�y�7p���C���C� =�2s�t�5��}���&lۼO<�8���+\�n����#L�<�Z���blߵ������%���Ԍ��F����oǧ?�i̜93�D��,vc,��3�Z<�m��Ld�8�+E{�����q���oq�F � @����l"�b�E�U�9�����ɓ<�嵝�Mlǉ�7��:�dK��%Q�����;)�"	6�$z�������������������������~�6dddH�SsaP��7��i�T���`soקUTT��w�U�m�Ѧ��7��|u�+`@�O�<	#G�BwWW��R��
ٰ���� `�b��=��x���4�V?�/>A��S}J��BX�ݝ�����ZZ)�[,Z�����L�m�p{�����޿9\�
=�g�G<����\�Mk���;��==��W�<��qIȘ�='���cİ������hn;وȮ��M|`e�]�]e�]>xv{��J�ng�,6b���Ŧ��kܩ��۞�F�b��{�{�Ɖ��یx)�bf���]�����{ݷ�C�
�Ƶ]H2VI���++�p�����F(_�@",�fnhi�����D�R����V߀"�HQ���c�
kwI�K�{�����X=.�\�v�l�`Sȭ�|��ʵ�|;�/e���G8t�V�^=�U<��U��*++�i��?���'�^�ąAKcϧ�E��2�ca�������?�<Z:C�}~�1��ŝ��<Al>|	��d�;B�{��?߄+����G��M���#K-mS������K��;�Ǜ�ת��_��7��5L.���������@�=��B뽛HMM�O!���)��1�"�/�:�C�7��#��D�Ň��ۣ���z&�c�>3��D���23��6�U>�K���@���i��1{&j+>�Kks3��o�X�3j�KDj�3�8Ю�;�:���@բ%��^���\�f�ύS�����!���TU��$�lև`�1v�u��Zo��7�`�6��	��:xP�������c�NKG���5wj�>O�`�5��,�N���v`�������v��Y���E��#v�c�FD}��u�~��������(d_�2Ɗ�1�1ݍκ
d�OBsW��">��}�S�ڈ. ��_��" M�.ua���}P�V�op�Hs�Н=��Q���v
.�,_�;0�d$��8K��|8k��� �=}��|����+n��r��,�0�Jd/�c���ra�I}t��i,U��)TT���1y���P6�ӡ����!��'�onh���_��s�ȏG8vE�&�I=��'o��n�l~aa M�/�&�_��%/nnΝ���5�Ǎ+�+%CV�~_����!5Սi�� {D�::p��yܺqӿ.�G������FӨQ�t�y�v��eÆ������?[�6�/¨�\�{�U��bbm� ����{ܭ���S����X"R7
�=a�h����{ow�:cŔ�ӂ����kZ&��pߵ�$Bt�;��\�'O��aÇ��	۵�Iru�i>��>}��qص]Q�G�Y>�[__�LfΞ�_����d��g6�>`~>k��e{"9�!��Z}g��^W������ݮw,vͳc��+V8���M)^RR���Na{<�U���U�"Xe%`�ڧ}.�C_�8 � |g�_}Ъ�
���	�`����~��h)�����b^��]����]A��4�E�/l=����[�c�_�|3�k���|��6����������)�q����������?�����ę��z�𱲰=u)��=Ԭ�����+�s�L���|��-b�S�9�ivo�s�N9r$&"�HaO��*�����Y�U��+V�%�J�7&/��1Ҙ���v�S�\��o�3:��m+����P�����f�x�{v-M_����p��p��ܺuK]�b�c�L�Z����Փ�]���<vv�c���gBܼ�<KF5M~M~~>�-Y���L�ܩ���e�pP���<+���卵���}�����x��H������fw�������~�����ٳ�ڵkcއ����c�}��5�ZSl�¡��}3%׍��{HOO�,P�.\�ʢs{�E�����x�����?u�v��"9����V��KD�$x�߾�,�N.�@'��ۥ��F��¥�yė	���/'���g"��'Bw@�:ydR?S!�XM����ן�r����̵�@\9j},�ݟO1�i�v~/�Ǹ�QܮK����׎�<�|���aʄI��6�Ο;�{�� �E[[~�sj�����%KT�{cK��b!� ]K�?�e�t���	��l_��<|5��>!]��b�(���ZYKE��mR������ }� ��R�:�|���˷�5��'{5���p���9y��p�6mڄ'�|�A�x�xB��߷D�.wrOᖠ��������
���V,��j���nBvÞ�m<�se����z
����I4�?��?��wPy�	!�������o�u�D"w&����D���w���������r�����o<���n$���|�����~�|���1�8r����p��A�G�n�2um9�f�e0ƒ��M�!͇�[|$ʽ=V��v�&��/�& bu���[��U>+W["aQ�2�u��zI��#$���~��.�ʷ����gW�Lp��x��<�S'MƤ�	�xO׮����#�uf.�j�69��so�Lv;�=��*_+;��X�����'�ϓ&M§�[�=�
�ߺ�[��b�y����z{]��[;�L�[�qE�1g�|��gh�;���cg�v�mV>��i�ʕ�0��6�pqW{%}�2c,S�{�����p)c��	/$	�1Kr;�Q�2��F��U����(^\�}�,X��`0�������_���)av]�X���=^�.��+d�v�ې-��D�.#�w��K%(l��[�����w�K2�ORw%�h�C����=$u�	���g��X<N�d����  27v�P�_�Ż�K�򐺶����4����V�o.�d��۝����dg�NMvl�F�."�0���W?��՜y��FyU��t�����=�h�!F�Ǘ'�hݲ >xK0䉗k�T�-y��򅯿���Y ��(�"��v�9QM����#����$Ͳ���|B|��}��O�j�-/E�W��uTWV�����a��^x=��:��l}"�L��Od�I�U�����?�`pq��|n���.�����_�-y$"8z��������Q|~�\V��������v����Dh��?���Ϟ�>���	���o���Q�P�W�����?���4�w�Z�[5xy�)$�^���o~�׫��g3��Z?xq'��	��7����1V3,��3�
�o(�;D�������m�x����a�\�~Dr0y�4L�91Ta��.�3i�Qv{w&f@(1�a3���+L�6�^���N��p� ���̹�hlh@��� ��ŋ�q�F<��S�	��K�/d�;;��jB*��1�!�� eTf
��k�#n��� �G̘�ۍ��@�&���c鼠O۱c�?��T�>��(AΨQ&k���˅����ɒ�z�]�}�v�>��Y*l7��Lx-�����˅�<֮����ȵ]��c�n���o�h�PE�������yy(�/ �B=}�::� ���b���ôIS�k���rQ��	>��	��[��\L��[1���<���ۏU�v-�����i�x���.�g�K��&�NH�,l����k;���w� ?���S�Φ��o�����`���&�K�����U|�*(r7��vj_�ߍ�O�
�����[��1o�h|\K�*"9hn��w~��N^ŏ��2��s������?{{O�<��u�����`"�dvr�����]TЬ	c���hn��s�K����g���'��6��k�jr���tu��/�{3��sA8���;�0�sHc,S�w�s;����Pt��xϭ�%��QWW��^{Dr02'�K�� �"ƍ��������chooA$�<�VvM]2331���\^U�+���>�	b�����u�hnj�l�����ǃ>��}K����l����ylJ���1�n�A�A�����y��v��/H�O/�2P�|�*�ta�qB�)�y����n��W����$aڬ�4m�����v�0�DH.1�5�]ShJdA��
�QP䬭��(_"0����v�A�:*�D]:'l��R���k�"pmαx�=�}��v]�>�6T���O��|*b�ظ�+���q�����=}���ܼv���{�X����`KAA,Z���lܮ�@k[�(v�a>{|y���a�(�H.O<]������D߶�1Z�vA�Ο-Ͳk;�|jJT�L�,����	�%?#�N�Y>+�v����B|�k_�+/�����7��g?�Y�?~H����b���`PJ�˝�mOc�*���

�-�����#��qm:"�xs�9��^�_���1k�v��?��P�L�D�|p������X�����a��2�e牫���_������7��BZ*�JI���q��m<�?�_��Ӹo�$7�����ĥ[w@�3XR�Fks�32C
�������f��r��;L1��}�@P�.�/.�i�!t�v?�楗^B}}=�ÌWV�_����P!;+��C�;W>��}��� �BGG�9�~�0q"�_�=}�8s�<ZZ[ACw��k�`����%C�SSS��_�>�lT}x���hc,���P�7�"�9�A��A�;p�Vy�#��]��)e*>0%����E�8/�$K��~�|�M\�v��ۓ���QX�l�dM���r���AA��7�k���}��� '�����k	um��G�W�O(���µ]���=��A\����K��z������)���҂㇏����L�F`Ͷ�sa鲥�5u:�5֋�6?X�D�)
�%e� ި��%̵]"��$�GV鶰,ngI����xq{��5b�<�|��Ua���*�KKp����!gÞ�/������>�6�]��*5Ű^�T�)X��S�ۺno����}�����Mk��Fa�4T�� Z,��6��)�5Y{/n�H�ؑ�Ă��s��o=�ov9RB\�N�9!��˻��&�C����/����O��>��z`<~��G	-���ǎ2OwOZm��%& ��^�o����礶�u���K���������z|���Iq��t����>H���`�N�uQN#�05��ݩ����b&x7�����'�'����vh1c��dro�~nܸ�6�H��Z���`�ݧgϘ�����؈c�F~�dn���Kzz:.^�ޯ+k�q��U2u#=#G�`��R=p��y��W�裏���hH���TQ���fc,���e�X�d��@H�>Y=х��.�[��s�\���b0E�/�k�!����8-��}3����_~�^�� &�\�~�:�'z�vN�n��X������]�k�v��vH*܁�8\����ܲ�]1�ת�=P'����!�G�O�D��mM>�յ]~q{aA�

��vl݆��~D2�\ݏ>�~�>cF���Ģ	�]Yaȗ�v��[�{ty�u��k;�ñt��pm���F1:�SX��)䋽�]�ϣ������k��n]�n�����O����(���|��x�'0o�<
V!x�V���ԃb�UZ�S���Yrd`"�^%�c{�^�Y��Ld���u�[4�4��C�wb(���oC��w���M�Z��l?	;�����=�o�;����()��d�����:�����@����ϣ������=�4"���:��O�E�c�����?|���ͦ������C��d����_���S
s��l@�W��5[��濼���^����O�pt��م�7��K1�-'0"3]�j��kUu��ߢ�N�R4�����:��D�.��ٞ�����`<Ÿ(��+O2��t?���/U�ٴ�4�f��b���<�.���|��6?��ΜA$]]]W��EEx`�Z4�����b03a�$ܭ���+4K��ь����!�F�X�c�rm����1��d��$H�>��C��< ҉A7͠��H�Sf�*��bD�-�>�c���o~�ܽ{��)�o���K�޵][��+� �tm�nle�vU�l&����	�?.�G�.
�9=#45�Dr'�v1ݪ�=&��|�$_�\۹�R_S0}�4�de���r�ܶ1)�z7o���#ǰd�Rd������T��C��M���=.��ϣ�)��x��C�fq[X�C�̊�k{0yyѹ/M<��	�}k�x4���{��v]u�y��R������_~���N΅M�����?��e�y������PdmH^�\R�a���`�*��B��j�F�{:i�NU<�������KX�`�asm��;�۽g��p������b�K���{�ǌ4�?r����7��i�t�Ld��߼�GJf�ϾxM��D�|t���>U�K����. #͍����w���k����u[�����g����ϞT���0����Vձ|(Q^ۨ�K����0oJA ���_�����8���o��?�����gJg�I\.��>7�_wƹ,�g����{N��G�Y,�UdX��<���l����p6%���'o'�֋���jz�i���M�o�m;}_a�vk"����ɓ'�k�.�'wL�.^���>�������p��1455� �꒕��qc�b��8y�4��i�#bp��d��Յp6�1����#�#c��c�u3?��?�(XQЇ�i��� �� c��T�46 #C��.�XCM3ȋ� �T�.� ,z�*j�e`���
o��&�3�x6
��Ңwm7���K��ǵ]"U���%K�Q��x~d�҂Չwm���XL���r�JrC>�$� ��1�k��p�`u<�܆Ӯ݃}�X�~��b�������xu5b(��mߺM\���"gTʫ*����� ���O�	�=b��\m���u�z���D�����DD��n.l7�v��HωGH�.�I�eq�\@�������/�$�uq����qEޘ<|�_���
��9p� �9��+W�&H�?Xe���`���tc�
)\�t�f"w5�D����������`��/��U|���X<�	�\�U�7v��E�����N^��k�{��xd�����������32b����j�$A���{����U�a� ��o��U�e�{�syy�)ܪm��|6#GY�=|��E�9u�m���E��\��
s���^��}�0f$��:�ܦc�r�Y�%u����}S�/�5N���/n;��^z��l������X�h�.����3Pq�I���(�<��+�j�T�Z5�2�ۃ}�b�a�i[NH�ԉtmV�dro��_�}��/~��>�w:���\w���&��F��ј;c6z��������AFZZZPq�G��E��3z�^��w� �}�t��޴�g�F8�x�����rc��˥cU!�=]�C��)	 �� c����Xwo7��SR$��������|K����N4YM�~^z�%��(PǓ�;
�hѹ����6�]���N�-����u���ks�vQ�������-���H�G�W�Z��0ߨ�ET���C�1�c�iV]ۇefbެb4����ӧ��:��B��v�ڥN�[��ESǣ�n-Ztׄx?���C�֍�v�N���˵]�BrѺUq;$�,�k���|J�]�%�: a�o��ඞOvB��E����a�iy.^�Uk����πp.����_�%%%��@KJ�*�o�d"r7wc3ݠ_�n�B(`ev�x������o��T�GwO^�}F]�Ρ�ԅ �2�_R"4�n���^�"��O/%���֣��1t`��{O_S�������GjF�Խ=lߡˬ�P��l�2/P�C�W�fǾw�ޭ:��g٪Rd�A&F��C��Gc}�ۏ��~�P���8zT}�3w�ŵ[7p��M�`aD����
� ��9x� >�U�V���7T��y9��[3ƚ���7h0�S �� b�pZ�j���jY��r��Tza��yAV�[ě��D��֡����>g�DF+֮Q��d$�k�o��k;?�D�{�]�a.��"�%q�dP�~[E��>M,'�$7��H�I]��O����q�u������?{�[۰w�nܼy'NAu��ȁ��#˖-��)�PU[���V㵪��nE�܊ܵ]E7Ї�[��ĵ]��>�F�4I.�̵���c|\�u}Zt�L�,���z�ָ��|��y�~�ш��|�I\�Z�� ��޻w/z�!�Jv��I\��X����*ƀ�&r�̑������T59�AA1xpy�Ri�����.��=Tߡ�oȷ����<�����;���/�v�~f�-f}&�d��o�͞������7�Į�4ؕ��g���/�˴�����5�t����&`ʌi�WC�8��������$�˴}��G�ͮ�� �	���}�S"
R�������W��漠wn������[|8!��H��鼜ϒ%���������ȥ��rm���B�(c����9ѵ"��SXBx� �Ӌ�����C����E�\^�0^�gb\�e�T���GH��ڞ���y3g�|�w�:�� ��>~�8N�8��K�B���*�wt��:�^)T����1�Qt1�E�0qm�vF!n��%sm%nx>���vs�QU^��[#6�����G!X7�g��r��`>�ݽ���^��^����տ#��x�;t����0�3M\����*N9�k��{۵��SY�Ϯ~�������a-8�AAA��w�������0�?��v��0�k;'n7.|�=H���E��-[���ŋ �ͨѹ��x!b00s�L�8	�=��'O���999 �VV�.��������nC>����D�d>ܾ���ΩS����I��`c,���ڌ�8[C�XN�����n��~����.h�(.� Y�
�EA$8A�m�>��c��A�����)��%!����/�Doѵ]-�#�{���n���ź+�W�*�	�e�p�w]��z��IZl]ە@5![ˉ�e�7�l<}-��RQ<s6��{���>BGG�{V�:y
gϜ����0{��WU���w)�\�RخO�u�zL\۹�,l�p���񣜴��]����g�fY�.�g"���w���[�G/��1|8��������\.]���[����=��}�i�! lS��I���c�����t������g6ژ�Sp���d&� � bp0!�m.�i��l0�6�8`��O���Y"n7������4M����/��2g�Nu��U�o� ����&cƔi�x�cl;�A�S]U�.�&M§�[����q��5D����'���}}} ��/�K�[�iii�w2Ʋn�%ӷFl�%���c�ц�Ha?$p$����܉�����9q�4��P������'	�����_��4Έ�l,)-7�W���3qQ���xѷB���e�vY�|Zl�b{M�m�k@$��ω��t��Z�;׵]�}b\�� w'T���O�wc��Ӯx_�\�3s�S�8|����AD�F��#Gq��	u
�YS��Bw�,�iq��h]�`-�?�"y��ۚ��%�)׻��uH�Y�vm�ϱ��{�v}]%k,�5y��XK\�z>��	Ο9¹0��~Xm�1�┐��oo�5��U27��x�_h���v�Q�J��µ�Y�mE��@AA��d���p��i>��C,�}�f��C���ͱ�&Q�Yy6l��7@8�ťˑ���HV�L���i3p���ؾe+��έ[��eʔ)����e�v���Dr�������� �KYY�j���㏇�_\}��1�2�il �X|���n5F���v2Ʋ�ƻ�aѵ]V�B	��`�4���=�/@�n�<NO�~�;�����p.�w�b�j��o�:Y�N{lUH���%����[��[�R��.VS�򺛊��:���a]Hn&n7�cE�����˄��r�JrC>�$_D��2��(Z��#�9��P��Aa���;�\ձ��#h�i�"&0���C���ѫV����B�WV��G���!^ky�|f��X����B�"�ܵ�w�t�k;�ٶ��'V��r�
�#�+}7auI����eܺq�M� �	����{�җ�dk��,-^��xQ�)>�_� sd���)��z��̉0l��.e,�<!/j� � � �S:��u)����Rhq�Q<R�-��3�Pt��d1��Eymmmx����E�2i�L�:��L�03&Oŭ7�e�f1p؀4�L�6�{ ��]Ey�mD�1m�L�Vՠ�v��y�2Ɗ�1�|�2�"i7�����6�d�C�A��l7Z�� =ݚ{�!H�2�1�"���휸ݸ���I�x��g��N8���`T��w��V�ߘ��Z�+~��k���~�:���V�����u@�/���ta�T/
�4q� WO���;�x��i�X'	sm��! nl8���S�"od:��&{����o�>�U:֭_��a����Њ@�.�!(n�%�H\�%w]i�"ӗF(n7�y��C^+�v���{����ػ���)j������Z"�2|�|�o�����p&�~U���琕�H�;X�� V����Bw�w1h%�nP��q��.��A�r�{WW'J�Rq�6��EAAD��N����:ҙ� m���L�Yt��`"�El3�8��*V�������\�g���� �d�pl��*��7�k�;�_��.�s�����ŏq��]D2�l�
��`3:�;@8���r�����l���<-^���1�g�1VjG���)�		�%��誋̹]&n7��%�Ԃ0�ۍ��z������}����	���Ɍ��Ys��u�:��ت�\�E/J���<f�v~[_�@\�%�A��ZZwSq;_��\���k}�`5ż��Q��,D�lh(�|>�x���|@��O�0����[P�����3q��y�<tAğ��.�ؾ�F�ªի��׃�u�L��V��rm�܈���vA`nL���o���G&l�t��@d�v���E���s����1pm�y0m��}`=>ܳ�3�s��z�-<��3�V�`���]��Tƴ�jS(`��x7��`� � � �����i�c��D����B���?T��!�W�XųOO��Z������p.췺|�
�SI>A$ÆÊ%��\߀��w�G.]��O.}���c���8x�:;A$l���W�Ý{@8���G%c�c����l�_��ڱt��*{@��В�TՅ�ֲ�B -���l��pn������ro�W��`�u�|�
��OO�]�%Jt��\gYl���ĵ��R"�6�K���(:M�nȫ*7��3{A�D��.w�W�k��>�O�������뵥���_\��������to!hhh��M�0s�,,^���5hmkU�yL�Ӳ����KH�k��B>�Ԕ��p�vm���Ks7vc�Y]��!B�ɵ=�5������K�����3aS��_@vv��ݩ������f"w��]�� �vPk��E�j��E���h�AAAD22Vi@��m�Kߎ��w(k�	�7�6|�a<S3�ЯhV/�oXWW¹̞7y�� �d��w�.X�w:�݇�]D"`��sgϩB�e%���=u��� ��_X��g��+ ��ݻw���o�w�w(*��XVL��n7&�5�2A�	ܓ�U��ֹ0D�&�/�J���T����*�o2�%�.Nvo߳gN�>¹L�9Y�Y�f�/4�q���\�e"k-�~[3q��]�C��T�.�I.���Wz> ��µ]Z��v1��'k��>���n���F2�����;s�eN�A�˕˗q�����b���v�8V���(<7�G#n�l+Л	֣qmW˒
�c��$�ĵ]��Do�	������=��<nw*���o�?�	X
��f��drq�E�^į'��4��V2'��������X�xi^*�@AA�tL�q���Խ�l௹1��H ��d��0��3��8�o0Z���ذa�=r$��A$3�M��	�q��a՜� ����ݍCDNN\�5U�t�DÄ�Y�t1��Ԣ��:@��믿�'�|R��0�+�1��g7c��ZfMCuc�	ܓ�|ԣ�saH1	T�#T\:q{�i��(���`Uh�����h�ÄC̅�p.�y�QP4� ����L\T%��������PBtױ:y�-e���g��.y[�K���=$�vUyi�k�c������Q$e��L]�����8���]۵X򔉓0nl�:�zru!G���G���ӧ�z�dd�����>��$6�C��s�`�_ [�=K�"��+FQ} �xێ�k;W� n��.�Lخ�9��c0�#�=A��f{��������#��,�n��)ʟz�!�
&�ި$"wM�n�������w��.���B������
�)��C�B� � �H2���A���{�m$�K�7��"w��1�P�k�����HD�T�oy��E��d���a�칸^V�m[�� �ill���;0i�$<��~��p��o�p0��d�J�ٲ���
sq�w�ˏUc,m�gK�X)�����,ۇZ@�	ܓ�i�n47�I]Rn���ǻ��+����]��!
�<g�b������̙3 �Izz:f�-&h�A3gT^T(|�BA_^��:�/kБщ۹􁺶+!�n*n��k;$�C��k����;/�O�k�$���0��Fdaa�\\�pg�� A΅ͪ�g�n���㾵kQ�Ԁ����z����v.ђh[����bw��&l����Bt�$-�7&�v]f��ٶ����ۍ�ʵ]�j1�髩ٻ���t�o<� .�?��@8�z��w�j��ؤ�׮}[3�+�̍��R���lf�~��u�>�#�q�3q�xWW'V��ay/� � � ��47��X%�q�L��3B�ۃ}����Pm2��ݸc�z��_���{��{��)�4#Ff� �Jff&�/\���&�ٹ+�ށ ��s��-���c��%X<w=�ήN�������sq��y΄���O��Xc�I]�����-���S
�K�Bl��I���Nt��S))a�U)~��@�ʕ�]����S��� ��;�`��?���Ԩt0KV� --��/�Z͊k��R����Pΰ^'l��[J�إ�v��Zs�5�K���=$�QW����!��M�����.�'=0���E�v��.��M~J`|>��9�̜�t�[u]�룩m"Y�s�6��6,X��g�V�mt�#�ik��"�<!���$ك@���|>����O�k{�"x��v��]ۣ�`]���]�r�M���vr���?�Ia�����\����[����??Do/	v�V=������V��`����Py�˰�RGp�^��9��J��>� � � �H�Lp���7`����,�Cti���>�C,I!�@�7��b.�X��D���|��7ɽ�����#���T�[���G��G���� �{�:qX�z���Å˟� ���VU���=΃c���{�ַ�R{��$W�`�4Q���1�oq���f�}!���~Cf�UZ��A2Ʋ�')�.ݍ��\D�vލA�j0d��T�P8I�� so?u�gR4y"�O�����������8�Y�v���,�Nt.�˫$<�<��O�ĵ]�ˏSVnT��]w�ssFaެb=rwjkADrr��9\�z>��:ۍ+-��KEےm�qm��Fat4�u�>�m�yC
�u����#I�ۍ�v~�yyc���㽷��<�`����o~s����Py�#MB�2�����.�v�>M�������i�i�!AAA����:t�ܦ3>��~�3>���Ӻ��j��a�C���q�0=�fXx뭷@8���T�ܷ���������ƪe%�p�<�ܦ�	"�������{0�����!:y�m� '��뗭^�]����Cy���Uw2Ɗ�K0�һ�{ۿ}C,��V�o�FaJ��>4���=IY]�BoS�%�k]���]?� ��`U�nħR��Ty<�4`�.�3IKO�⒒`�U* ���M\�Ec֠��߫�=�ϸ�����E��Z*����a�Bµݰ_]����qzd�$�#6��&�u�\π\�ŀW�+����s��m�n��G"b`ttt`�ƍ�2u*�F�Fzj:�{����8½]M�=Q�n*l�P��/D��<�1"�)n�۵=Z(�{�哽���!B�,X�@oR�uq���V�Y�sg��z�5΃�łUYY�����|N	8E�&��h�Sd�`pJ��td`���Y�J�^hlG��htn5� � � ��L�FksC���%�+��{x3,��v�;��%}����TN�ӋW����F���e���6|8	�	G���-FzJ*vl݆��~��TVT���
�J�ctv��8�pY�٘�p>Ο:�y�1V`MXc,��P6��K����#���f��-�P�5�-�~�hH����)��\t#HB�0�����]t`����k�!�����i��4zک,)]���t�Z���Ep����µݤ���U�D,:L^��\ص������j�H��:�H�ڎ`Q!��Qsc��Zrm���--�/���Sp`�~
p� ���U���by�r������ڿf��*Ҥ�	s�(���=��`ސ�v]Fö�|�\ۅ<�|\���!M��״�S:�N��t����em�/~�+�ɿ���4���`S���;�`U��ݭ��/��LD��E�� ��@�"���y<-5p)c����AAA$�Ey=�g>�W�w(k3�	d���c��oێ<ɘf����6l �L��b��� '1&w4�-\�ǎ�qB� �6H�ؑ�HOOǂ9s�����M8��s�QUQ��;��t"d���	o�e���h�H��3��O�n��?@|�~lj�`H���f�F�\$��.��L(`X�
�E�􁪡����1�vr_v&�E�1a�$�D�m��-lε:��a���Q����e4��Ʋ͎3>���9�����^ʱ���+͐&�� z�v.��v��d�"�VW���A^X�j��m�0aV�^��;5�û�ޮ&��۵�5|��\�u�yq����`����K�2�����p!%��>i^�X�\p?fL>���`��A8�z��1b���@�N���G�~!�o+�wi��_*�0����}yu3��׳�d�KŉJBAA�sq� }M5 ��@^i[�\��"�4��v�g	N��3K���o�[��׃p.�O����=�t�2�vucۖ��9 �AHCC*++�?���g��#���A�{o_��;7mE?�&��\ܿ�o$M_aB�� mT�K�Whj$�kO��ZZk�w��>��0H���,ۏ޺`'��T���2�v+.�`�4P5t\��:�cǎ�p�iiX��DP{��jɵ=�?�vA�.���9��*���@!\�����|V]�5q����$�XssFa鼅�p�>Q�JĠ���ۨz�m���~�����j�\��4�ʟf�G.X7������d�3��vq[�$-(n7B���=Ξ9�۷�A8�z����կ~5�A��m +�����q;�'
1|�b�Jtd���'N�h�	d� � � ©,����.ddd�S���?�c���!���5��,-N�k477��7��L�/Y�~L�����q(�>GFKف�`��+�>u���XW�
e�7Q^qa7Y#�Q�`.�>�y���+��;c!l�ahc,En��}���%���XT����= 	ܓw�x�iLSڈ�8�0���]�o�A#���e6,ӐpI�r~�*e��k�O�΋��ڮ+Ǫ�]�wK���vC�%�z�8]�����D&�W�k;L�)����^[<}�\���۶� ��saؽkƏ�5k�Cyu%����qmW��{9����&���u�d[k�v-_���H��d�3HO(�ľ�Ƶ�b^]��|L����~��Sg �k_|�_P�-e8�Q!�i�����~4���M9h\�-��R(k?Tz1��sk]-FeNAC]+AAA8�"w3��n���C����X��?�T��� ��&����<�DRg��ΜZ	�;&�f� A���.�3�2ұs�1t`���ڍ�`M�J:~��iۙ5�U��PG392�
|���g�e�m̷���i��pi 	ܓ�Ņ�hom�0H:��S��ȅA�Qsw��c�v��y|��G �G��BL�:9�]�K�r~tB�D��C���k�(����I^@�ڮ��k��H�ٍi�pmgI#G�`��blݲ�UU���AC6��;oo��~}#�q��^��dQܮ�	�O�����>�u+��y*l�ok͍�j��`4��������jM��ྠ� ��ضygQQQ�-�w�'�x���Ĥ��h�� �'D[5���2���I�*%��r��������~AAA�cTf
Z�� 5-U:����p����]Z�~@�﫾������+���6l �<�o�d�J�~�����\̘0�.\Tg$bhr��9dee�����3�[wa���ؽi�p l ��6�R��=c,��=�1���0\���;lk����h�r΀���1'lH{�K:B$N�\��`�n��M���qo'��������R�tWn�@2����9 ��ӄ�~Kq�_�pI|9F��_"l*�/W�2Z�v�X_f�8=jrt���O�|�E�R�����wmg�3�NG����y�F5�M������͛1w�<u�YQX��"O�˺G�g&l��k���$Ͳ�]k������Ͽ7�y��}0����{�~�>y�5� ��k����{,���@R����wQ�z1�PfV�vw׋܍�7��2גAAA8����z��Zǻ�)��1�����=�)����x�l����x�}���s��1g�|���A���������<r�H1tiii���[Q��S&NƱ�'@v12'�����s�p�o��V����<�۷g�1�L��c��f��z�;?���=V�K��} 	ܓ��i
�j�v>H%��i�1`&8�waЂUZ$J��ȅ!NRݸq����)������;UF��/W�{5������ⶮ�N���:���!h�f=�bf!U�s����y��+G�)���Z���e����._ՕI����ȮI�n�z�xKs�wi���2nb{}}����㧡�W/^
d�����K6f`B�����~q�:����W}�ioo��z���]S�655��͛����ݭ7���soױ3�<�������.v`米�\kk�z���k�NL�6]��o�D��5hjl�_T|X����D�ht޾U����o��ʵ} u��>盽Ϛ���ЋDD��[����}�;���7�:Uܾ�=�F���9s��Ҋha���h�5?��o�����~<��pjp)�4� ~Ќ�;��.f�
R����Li-��5&����	� � � � ��.�Y�!o�e���o��4��v�_����x��> row&#G�`Ɯ� �����}�+��s����+#bh��GAaa!Y� =����/����媶�p���:}�Q2Ɗ��0��d�g�Qf>����gZ��(H��D�,r��ރ�4y�{��z��=���sa��D��7��8L��a㋩ݎ��*?'w�.���M�\�����ѣ%��&��H\ۅ-}�n^)Ô�Ӎ�T�b�������#pm�'2q��Y3��HC'|}$N�fy�\�YBխ��?��c��L��zB�O�||�Z�¥���'_��9s��]���s�k{Ѹ��_�}{� 77W]L��Į�������rL�8v����'O�����F�ߜ{\W�<v�˿{�.�6��`���c���SũEEEa�vz�V�Z���
p��RM�ֵ���S�9{&��Ͻ��EwwF���L�~��uƆgĮ��Me�~Y��	�++*1�!_"\ۙ�}��حmm��;p���{�y��ڈ�����:~�(���۲����q`��߾�꫸���uלSI�[��K�78����N����b"��E�����Ơ�j�������t���AAA8���n��4###Cp�sE�w��l��uq{����B�	��X�m߾������v'ۇ]��4��Gf��0q"ʯݐ�okiEKSܩ��&��1�5[�fq����4��<�D�?zT.��x���͵��K�m644��4��|�g�4v�i��~����3�rV�]�;���ifx��Xݎ;�>��[[P����P������T�]���R~2��	�'��{S$��;����<�8��6�����
8p �ׯ����d�e����3���&�Ҳ�Қ�1-w4�Փ1V" �{1������;1��L��N����O��6m�,�osɊU�.<��d���L@&s{���ԯ3���	*�%�Ac<�t+��>5�Dh*$�i"n7��s� :���Mq���Vw�7a��?��瓈��`1�1��Iqa��E�}�&v��$��{�9t�*�_}�ܮ�R�\$�,EģO3�{�/���Wo1M,#�1��ݷƚ�=�|V�޺�<o��V�������{���p��y�f!�9sFh���:&�{�4�����KQ�>h%�vP��nɍA��94�4V#5e<z��AAA���Dg�[�p��
S�s��� �1�T������3;�Jc��z�~�8C�8��n��=^�O�5��3]_[Y������D�Dg�gL��l6�5����h�-��y�(��{W.]��ڻ�t�����3���ȑ�8es&�����V�ف������9ոq�l)����.��ܳ���3fL���w��K�b��I�{��*���~�3�d�!6��$�g3?�߸U��>�w���<���~��P��c����+�`ݺ�ɜ��
�j��ۧ����PhCs�� ���ݸVO�X���I¤Qn�6�#==���nű�X�F�D&n�[=��������r�3y�<Nx���)�=q�\�9�z��X�D`�龅]*�D���bLԥs�v��㔉����cހ�\vi��ۅ㑉�}*���2M�|�Q�"x��S�-��m.�8x@��G�K�9�,���{<�Au�����~m]hni�-���
u��N���h]ۥi����NQ}�U�j�/��v �jM�n�������ǟ~o����~+l�(&pק%C�i�if��N���v~@w�@�U7���N����AAA�M�KAwc�|��žC3w�8@�_���~5�L�-���E��δ������� �EFf&�-Y�H4cF�a���8��C�g�$"����eTUV����ȩhhjA$��%KQ[U��8B8�ӧO�ĉX�|�c��`�e6[Y8��@{��kzݾ�Z���y�?10H��$,݋�:]P*Dp�J��̉!.�$D�JcS'���{ �R�_��Dܮ`K~�qrm��A|-�[��Na-���]����]�%�Y^��H�k�pm�y�ߍ�vݱI��Ӯ��� �ǍǖM�b2z� ��s������j�j�E��Z�z���%I���桄�j�GL���2���ֈ�h���Cɵ=��k�(/]��G��ڕ� �Ç~��/bΜ9Ip�E�Q�΋��-fA*��g�C��f�AAA�ݬ.b3M��΀�����͍���ji�~B
d��x���~Cso'����K���
�H$�3faTV6�o��=� B�钶mي+W���W��� Ezz�:H���c ��f������������\�.���ٞ��nf��|\*�T�7K�P��IBJ�]�&��Q�n����T���
��B�mذ ����epkA*7s���#{ ��vA���Z�ih����vIݣum���`]�ײ�}���@�>_p���>\�(�7�$����\80q�@(�v�iάY�i�P�A������<y2V�Y�k�7}�$��u���|r�k����5�_�/_�I>������i�{?�;O�?~�o4h�Ah�����4������~��+�w��]����	�].�Ck}-r2������ � � �%/��n����)�����b}���/�HD�]�ģNgΜ��#G@8���0y"Q��a�e��s��AD����Çav�l�[�9Dg��1e�tܾqwjjA8��{��ҥK(..4"v�iF�����Bd�������R��f�I_H����FG{+�32MU�L5ȏH��Z1Tm���n��� �E^~>�&M�}�\�}zf�]�_�lTm��
�u�"qm7���#K�ב������-��k����r�:Q���������]۽N�%K���Ө��AD<�y�&������|w��3�.(n�!�4E�����O�f���{�m�H�v}M���g��ĵ=q{l�o-���Xǌ�Ǻ�Ǟ��@8�;v�;������ޗ�(�N?�����V)-����]?���G��B��� � � �6Fe����RS�B��[�7�������/�^�$ 2� ����/uz���Il�0�oq�rD��H���Ukp����׃ "�|r�����u`����>C��'�J�aצ�����4c�������#b��1���=E���$��@ߡ?�����&���ڃ��I���.t�����*E�2so���߅�N�����q��m΁����,��ٿpm�8���wm���q���Ţc�ڮ�3J�����9��#�Ӎ	�m���\�M>	'^	Vǣ�m8�
Ffgc��b�ٵ��� ��'l��o���yX�n���	��Y�^]#����,�ڵ=�zE ��k�l��z '�CsS3g��Յw�y���w#N�`L~�`A*�~��D�M?�;����r�6��`����ټ�@AAa%����+!�ۭ�bE��]��=\o^_����fR�\	g1k�1���Â�s�k�N��� "444`��]Xw�z\��	�6�sFb�외z�΁c=��(,,�z_N�So��~
c̱,c�wpWB��9w�Ѕ}�zA��;����m���B�a��~$�o��26��Ȳ�i��{��Y�(���#�ߴ���xKP]C&lק�E��nاt�M�k;/$GB]�E�;`��n̄�\ۃ�����w#C�+�<a�rr�y�&rc!"a��۶nò��1y�ܮ�����z�x�
��|��O�f��鶃׵]��t���f��|rzz}��x�A8����<���|�j'�dt��"bB�4q�<X�;1(�*]��d�\�Y9�n�AAA�d�5�C20W�X5��-���u}���ZbE�8��/Vi6l@o/��İ��1kn1",�7nO
�n�� �xÄ�l0Ͳeː7:�/] Aě9���-t�w�p���x��w�G�G��+LL��Q���3�c��!ۺ��o�+��{^
3�"~����,�Fwk���	"�
A��봗�D1���U��
�$`�C(�-�ĉ8s�琑��}����.�A�@[�݊�vٶ����������Q_m(�/DV)-��k�I^K��(]�ż&�<�|�pm�pi��d���}�i��-�� ��U�}|'� ����㨮����vu%����tc���$-J�vY��|�qm7����<a���&N���!�-X�G�Ƶ�2΀Mm�e�|�_t\*�ei�Q�7-`�}6����~]�"P�:1D�.,��AAA	�0+-�u� u���P�wy�v����B��=`��`\G�o(�?tj�_,Қ���y�f�bQ�R��$� ��G�)Y�[�n�֭[ �H$L�4e�<�v=�<��>2c!�Gjj*�.Z����pl��o~�៵h����iA�?}�>����2w��tHM.7����FeNECG?��@�;�31��.�(�S/H+����a��d	DE[>sM$�fg�`�b�ݩ��o���BP5�/kU����ص]1�D���z�u ]^�ŵ]�7�`�����vC>Swx;\۵<BZ8�vv�,]�gN�DMM� 줲��>؈G{Uwj���T֠SG*s�0+���۵=�ےk{D"z]��������/<����O�Yg���o�駟���������ZV��$�̂mU�J��n^��$.�������_�{꽥� � � "�,ۏ�:]Ǻـݐ}��6��s� r�(��͈W���B��7����s�/,��	E �x2|�0�[����C[[� ��ƍ������PE�]� �x1y�T�,��{w�p��߾};�z�)�	���W)1���C���������ٟ��]���Bۯ��$pw0�n��� �`�5q�1 ֽ="�&Ó,��pTTT`׮] �Cn�hL�2% (7���=��Y'h6�KU<bz(�v�X^�.��È��b��.�ˋ�aP�&l7n�H�D�Ll� �v���ŐU_���4�,Z��{����,:	�p,`�����㏣������
��v+�vc>���\ۍ�����s)��[���[�ApA������;v,V޷� ������GaݺuI+b�4���B� ��o����e��pmg��-l��؀)��p����'� � "��uԡ�dj����B{�Z�ڦB��P3��	
���x�/��������ouq�2D<�;K�������1� �inn��m���C���3�oh AċE%K�{�v2�u6l�O<�����Kop�����Xs,����9��)���K�AM���.����7D| ���)�B_s��P��.sq{�O��nezAх!<��
�ƂT��� ��=.YQ���=2I��k���a�w��b�mF�/QShG�ڮ�7�B�(]�un�>�˫ ����+�ε]_a�����o��������9رu]�A8���wՀ���l457��Z���t� n��]ۣ���A�e�Ć�Y]"��E��ȇ�k�,�C?�S�O����3x�{�3����b�2���*+K�`�b�2L9�sF�?�7��� � � �2-׍֖fddd����/������Z?���e��ϲ��ݫ:��az�,d�$Q	?&M���c�c׎�$�#�1�>Ý�w`՚�(����JD<���Ŕ�p�Jgp��%>|�W�vP�^|�7��ͱB���K��6��̌��Q42Md�H��`ƺZ��rK;�C_\���Aޱ/����H�D�CɅ���]�f�p��OC����tm��D���)��R�9/�W�A����!/X7�S&�WT��KC\�=��uTI1$j��g�1�T0[6m� A��ݟv�܅+W �`,���	n��5sa�>M��]�%"x�h���/76��Q;�'�k��,9�6���g��[@8����˘5kV������1���Bwq�A޽P	��9#���zK� � � �D1?�]u.i�z$�X�@`����~	�dcoE����>�1�8���L/����f��I��?A��`�$|�%˖"k�\�r�.^��7��C&���w�Q�N��ބKb����+ |7�*��B���ںE�}�hH��P��S��xGuo�M�n�� t҇R�tr��t�v��_��i�&ܻw�3`��y狢,�k��z���#����k�V�G�B����J@6nH7��<"���n���W.�W,����%"x�x��E��n؋�OwP��L�2q�S\عc� ��#���x�̙7�5�j�(E�&n'l��(6@��؍��sm�ZD��H��$�v>���R50z����h�K��_�����B�߯�@k}�5L�J�&6�.�ܬj�m���_�wȍ� � � ���(��ܕ�b�3P	��|��8ت��8(Y���<'^��.��ѣ �ü����
��%�����]�]%�Z� �ͩ'1s�L��u��ID�IOOǜ�p��)΀c���a����ǲ|�1���o �X�L�MM�t�r--���[r.��Cw��b�OL]�M7�@�Tq�J�q� =�/��F;��s�=.2�3&F��.�������#qm�jl\%����k�>���ntO룉�c��.�'�{N�bH�;s6���� �H&.]���&ܷn-�S�tm����ѻ�G�w�G&X��W�/ŕ��>�(^��@86 ���1j�(�{����W~�aA*�t�)r�>ՠ,`%k��\n�ٍwR@AAo�MCg{��Tm�K��z p(3�@���=�dxe�o�������IӦ� b�w�_u.�;�ښA$W._���qx`�Z�=x��ND̙6{&�]��֖���۫c������.��vc�V���X6Ɗ��P�����{��8�3��IV� ���pW�"EQe[�eK��ܖ����ǎ��wt�an��|�ϳ����;�s��ZIJ�7p�DQ�DQ�	� �}���UY����D-�
x~VU'��s������y��@?��7��i��B�{�R�>���0�,_2��=� UR��,'��|�g��ӧO�ƍ �Ał
�۴�,��n��$~�r���VXk����v�~��'�>�l��;���?ˈk��,)�t�x�ܶ�?����!�"<��={�֏���A���z��L&X�������N�S=�k�;*{��N֯_����p㫯A�3<<������ T07��L���|����=]�%+�M<��9~L!�B!Yd��Q�N�FX�ܡ�jT�A��/�c	�9��Y��fk��ʺ���o�>��a�s�CM�'$e�exu�wp��qR�G)0>x��a����q��Q�ID_b��m8u�8H~����#jjj����K�M�c��{cY�"w���xl���7��d
��ڊ"�<Ei��TЅA3��I4�A*/��$R[Q(
ͅ��M�pFc����m(.N\��"k�k��Ĺ��w-�v�X�v��=^h�3Z*qI�5{�Ե]��.wmr���<��%΃];v���sx��B)d������g��ס��$�����v[��vؚ�ڇ�4O]�����+6ۮ���'�����?����>~��_'�w*l��OM��:1X_�'��I�w�[&"��ť��9	B!�B��X_fb�I�O�N��.�nu������������e�C�y�l�W�}���Z�-ES�b�I�V�坻pp�LLL�B
���~>p���uܺq�d������Ԅ�O���GL�۳g~��_�+�1��ϸʴdް(�7�\-M"rǰН5�d
��-�/J��l�%�T��|V�T��*�� ��H~d�彳�G����b�Xb0-�v�l��N�X>�퉢�]�����rm�	��2��n����Ů�xa���8~B�B�\`||W._���;046���Iq{�\۝������]۽�0�]۝hiY��/<�s�ς���͛�jS�w�V*b�����qA?%����čA��En�Bcx�%%"�H�k��j�ΒB!�B��֖bL������8�Cw��ļ5Q?�|��4�>���<`��;==�c��@���=��LR]U��݁O�����!��9Cq=k[����?0 B2Ŷ�w����h�'������/�"k䣁Uf�+��*�5�r���4k�9`�����#�ho,�W]S ���<dQ�����9H%��bj�'*���� f7�����[wn���E�u@�v�ص��ێ�%��$��rc��n��m��䳬���bb��w���Z`G�2�ɶ���կ�=Ч`������l�\�ni�k�Ҡ"r��,����D�
�vg��o���/c��Ey�����
'�L��M��C�����P9�!t�D�U��=:�$�����PB!�B�m�c+N�I�}�T�C�1���s)vY�I�:�X��m�l^�����q����`պ5�^TB2E]m�oڂ��|J�!d� r��~�-��?��^Fo?��HfXTW��m��{�6�z���K�={/��6�2���Xz�=(�1���.���ҕ���X���5S��$�P��gT�i��BII�+q�=@��`�A*�c�ʌI�nՃS�n���>��#��`��%hji������ۨ����w�M�vc�A\ۍMA\�ѹ���y<�c��y��%�w��5����Zk��D��a�vC/���w���O?���!d."�e���?�'o���؅|tl̼�ˊk��|�\�>w]���e޵=���=�������k����O@�s��A��?��.]��σP�߯�QC`'�>�L����>:2������$!�B!$�hZ�]Rw8,w�l��_Ja��r>�J0H]�m�1E�yBII	6<��d���&<Ӿ�����2��5q}{�W��W����B2������}LOѭ:ػw�.p7���XF�0�1�S�n7��qsw��c�Ǟ�Z� �9(p�3�o)�4���P�z}ø��h�G��2��L���ѣ�{�.H~�L��-����P�����̵=)7�#ub�	�-�s׮�qzRk��K�f����vS�n�gݵ=/�2  ��IDAT---��gw`Wh ����������?}[�L���H���_Uۏ��>L�%l7��&=�so�u����h��M/�et?���a�LLL�U��[��PA�<]�
��]wX�d����*M��v�2����XW=�/��B!�B2��R������B�']�J�$�5������=_h�/y�l��?x� ǎ��mڀ�
�	Z���m�n�E!sq�s��a�������o��q'I����}-��vD=���׍����=ch��'tw���9El����A��[��=���)(p�3�!�H\�|�}�f?H�ωA�C{�\�{;gg���VbQm��$=�v�Kz�]�e��x�Tl�oʞk�T(���P��rѺ}q���-vm�|q�Z�⎝طg/���A!�q?��{�����? RY�!�(���^��Y�g��=��h�c�/-+�k?�>>z���������~�;�	
*5��Tc�*j�ud0���_���%nw82�Vڈp�i!�B!�d�5U���H�^}�1�f3ƒ���r��	B���y@?��/~�ᇘ���]�@Yy�lh!�`Ų�h]�G!��u�=͡����zN��}�~��ٰenݸ�ɉ	���={�����=����D�n�c�'��$b�'�����X��uS���!(p�#*J�0�߅�H�+a�-lפ_*���U�@�C��08eE8��<yD=�ܸuK�U�_���m{�)nw�G]�n �k�mC q��Mqx]۝��Ko����Ч��n;�D�s�\���w���p��45c�Gs�2��>}�!^}�UT-����`V\�eq�˹��&��]۝�عk�9���~��'N��W^)�A�p���V�_��A�V��g�'�˖tNH����{�B!��QF��+�%� �C�Y�f�%��r�����wOI��g��S���A��lIN�'$U�`I}#�suB�<���I�|~�~_x���%��X�q=�]�D=��~��ߢ�8.	Η�_:�M�3\�/��0��rs���M�D߼t�7ւZ��@�{���с��gwxT�]��.)��v�`$�UKi&��P�� �>��LMq��|`պ5���,��I��-�"l���K���\ۓU�Ɋk�Dt�ˢk�=�������nۃ-N���sm7��[7nƉ�G���B��>|���z\�><�ؚ�k���eB"V�HGܮֵ=��`=�>�܋$��o����
���"�ֲB�
��Ml��<��]�O6����-�XE��Gk��M7!�B!$c�o,���0���m�mgc����4��rq�b�s��B[���}<x>Qς�J=wHH��_��zp��iB�|���s�ȽdU	����k7��ͯ�����Z��oGG����#c,�5��Yc�'�k�m����K���C���1V&��=�h*�H�ؖ,���v�s�ҥ��b�l�w�C���a�����G��G����v��z(�vȄ�]�!�D2O\�M�e�RѺE��Ի���q9\��KK�u��۳'�u�B�"�[o���bhH��WSq��h�8?q{�D�����`�v���׵m�v=tO��@�"��ݻ�+Vx�� T�A6s�f~�����1X����1�	u{=!�B!$S�/���ӈ�D�$ͽ�vc,-i��7��O��웙�.w?�I�s���#L~Q��_�6nۢ�߄�C���(ӊ���#cB�5B���Xݶ7o�!�E���߲	��^ Qχ~���1���c� @9!l׵��9Ck���_�\7�;} ��<�4�/1���5He=�]�T.�T�]9�dKt��:��C8�vQ���%l**�ύ�&���E�����um�}�o�og���]�>�vm���\��m�曻�ř��D�L,���q�2�vY�]����f����`����d�^LOsV!��]���[XPQ��1�L�L���q����44���{���gB�t���G�"�����?�D-b��}����ì��E��=�~Խ]��`sd�LO%rO�1`e]3n�p50B!�BHf(��������B#?(q�2Ɗ�t��š=S.�n�3g@�#V|^��������*���s�A!�x�v����Q|{�6�-�֭�7׿����Z�;�G�����3f.�N��F�c,�O6����&�֮������D�[6�k�"����=O��R��i���H�4�#��Y\,N�A�t$U&q!��l�<8e��O?�C ��6mt���X��r������>����ԉ=L,�Y�vY=��>�"Ϋ��W��h"NK�h���g~��6{��G��%��-).Ƌ�=�=}���@!�ξ����O��/ޣ��zY:��a��abú��#nόk{��l��{�fGp�q�&,^҂G;A�"���o�F����B����hbl�N���ܯ�l,3�pc�<#�n��q��B!��6+�1<4�����vc��e�9��W��&��`���՞�e{�졁N��y�V����Xֲ͵8}�!���9}/��&�&q��2�}��-�q��4�Z&&&t�;�7,dw�p�����x-�/Ku�!W��EKU:g@҃�<aI�F�	���%x��̹�)�U�]�.�n�C�_Ygg'�?���½��L����yn-2��<�mv#^�(� �(ϴk�m��`�q�qm��M���.�w�m�pmכ)qm\e��8��ك��"�b�ھ{?ޣ߸Bq#���}���w03����������26[�����;c�9�7�������Z<x�;��޽� �f�s���;:����67-�CR�n�2���u{-!�B!$]��Mc�ے7tN��zXr����9�@&l��������K+�}��' ꩭ����A�lYҼ+Z����	Bqs��i|��W099�GO���кz%����@�"&���w�����|vgϥ1���]�W�����a��#�� t��	�y@$�����r��E����C��.�Q܁���/*�r�̰o�>:=��%�X�a}�\�MSp�!��#^����G%���}Kc��v��ZM��]�ĵ]K~�
r�ڞ�b��]�vK�%�6Y}��Y� n*^��8��5	!�x#�����?�+���X��q���.ͥk��~YdỶ;i�ݷ	� ��X�J܃�矻B�:mw��*xRe̍�)2�=��RՀ�A��B!�Bңd�ӎɵ�>�<�|�g���*�M���0�r�'N�����AԳq�2[�zy+���!��q����꫘��BwO7	��;lxf3�� Q�͛7q��y<���y)JOEƌ����c��E�r��Wfh�`�/րj����=�����8��+�K��]���\�Y%.��@�I\��R����s�0��6l@Y½=�E؞�v�����#�����k�`]�k�{��$�qn��S�!�k{B�8�t]�ݓ����]/���C!�������������������Wn/�����\���2lW|z��0��vmڀl	����o�����<x��O���ڸ�x!�+������ʍ��/�����F�1B!�B�cqUC��(++��z���'��V}����̱�h�G�y�l��d��� �YTW��eKA�l�]��׮�Ⴧ@!$5G���?�.|~=�� $,��Z��g�cr|D-�?#�A���X�|�o_ؑ+4��F�:���e�gC���ۍE��762{(p�V.���x$� U½]���s`���w��"��M�th�C�_�x7n� QKqqܽ��"nw���\�m�rm���]��h��k����|a�S��vmw�W=�x�-��v�:a{�˙^3���o��-��k��j�x�{��8q���!��azz�������:�cj:�<�k�v��P���ꚳ����� �{��^__���u���������^��
�vc��RirQ�ǀU$��Ë���P�/ !�B!�̖����POQ����?��#j�ի�} �����3�Y�~��B�%Z���ѣGAԳi���쨩���m;���} �q?t���x�7�q�,��B�a��v�"�Z����ӟP]w�1�\�n��W�,y���q٪k[k8z$(p��F{��x������q~�|E�H|�-���6k.	a�9�%�,ȝ�*�PAii���%%%���&<�wI��TP�%u�6�
m)�c�����zLQ�Ġ=4N�xow/����T���񑆛��+~@�O���_&�����>�"�(��2��m������K��S���e�[��������./���q��m�`rrR��/�ѿ���e����X�;��ק�~�Ǯ�~q���K�7G*�]|߆��155�����!���a�O��B��v�j����]>p!o�$���gltT?��]O=#�n��0����8~��_d�}�W%��ݻ8qԲ�n�z�4��`4�����A��2�os�!p7�WQz���0�֍�.�X��VC�OQV܊��|�!�B!s��� FB���XEvc,�������6�!��Bth��Ǿ}�011��o�1�'��U}N����n�8�d�W�T���ÃCY�{|l%#��Ψ�ǋ�Q6�Ϸ��9>1>���,�����,�_�۟=��;>�hEh���:�s���+\[e�����8�t��'ר<�D�Je��n��R5���;/�=U���;���^x�E\������W�[#�.^o�@��|]C��[��F���!�Vy-מC�����y./�ȶ1�������n��}�g���9A]��"B'�&>W��]1-UE�/3½�>;$�R��A*����pHN}�g?R�C�D���\���1!��'U������t�/>�m;w���~��n�� ���t��(�m�W����_c��u�*�@MZ��vm7�o|�%�n\����-ǝ2�2Q �޻u���(���tm��/�V���K���M�b����X���[�n���*�!�ljjRR�ݻw�b�
�B��U}�B�.�����J�Wy������;�⚯��.+?~�e˖)������G����w���\\��:�=t�}��@�ziڮ�w��t>|�M[6��cϳum+�����r=7��ux7˄����}''���؇��Q��{��T ���O��;w_}�����X���:g��`���1h�����ݱܠ�������~�f�!�B!��)/������D��J�;��~�v��A�-V�<��5,�6a��KA�!pW��?@+�Z1����q��+�
���*���~����ֱ�s�}�j:p333�qB�j<Oh�k�
��]|�)���B�y'�s*E�Fݪ�*?{q�&p� [�y��E����l�T8�j41�B����c��PW]c}rB�
T��}4�w�0�w�|sg����ጱ�&��D�F�:����?6Ѕ�e���etޣ��4��ڄ�2��e
">_������.���> �@�ҽ�(4�z�xq1W��KL�nܠ��uٵD`����v�J�����qM��܆���&M+5Z���g)lO��%���q21z��v�g� q��l��D;����L^p��W���T:dB�\B��p(vo$Dڏ��$��A�".Ll�B��;̽�l�~�*D�A�J]^o��y�N�m;��'�Q��^|��'��]�-�P�^fPF7���=a�pn7��81H��,��6n!�B!���ٖ�D��Y��4�r&�5ۄ��#E��#Ih��kN�B.�/���+W|����XS�˪@���Ps�8�d�/����M�^���4��`�"�!:k\ܬ�n���Z��?�.Χ7^����h}}����ʌ��6A����FI�Kձ�C�.��T��؅�Y�Ω����1��ÙB�g/�7�~q�*H��{{z�׿�5>=zh֓��d��%���������v���U�����\��.�+�㩼�����re�[9u����[�Z�������{c�İ�ޚZ�)�1i���=���cc��\�K�j&���qU�A�El�o���e��Vw���$�A���`�Buf���O?Q�����L<&s�tm��{	���b��y�<�k{ a��<}�voa�۝��{q�g�f�u�y�����I�v���764�~�4|~�*!�d�����K���ft��J"��{��ҵ�u�y� ���f��v[Que��˗�@cS��<Q�޽{�����U
�]!l��:��Ӊ�շN
݋��UIa��/?=$V�R�&�B!�6K�F0	�7�c��v3�n��Y��*v�2�rR(����b��\�ۉ��۶���|�;����S2!����s���/����N�����+׮��s@�!�5B�w�w�m��?̶1���՟5ӈ���]��(k���%���
�RQR���2�^��R7� �u�t���]�m_z��P봐�%;;;q��Y��n_���2Gi�\�=��β<um��~Y=q��+.*�ˑk����5�,��;
��.X�`!�5/֗�"��y���+�TWc���l	�d86#����9֜��=�^p�#�(�|�U�����@�����>}/��r^*eӍ������4.�w�va0����`]C1�~:B!�B	��E19�n�g�t�sf5�r����Y�B7�J/�e��hD-�eu��e $/>�<���s��N!�������?�g/Q�L��x�,��+��cϞ=����\A#�g�����c,��"3��9C��>&��@f�
��R��Xf0���I.��� �]�F�p��}�߿SS�D��½�JP��x,���p��ZC&\��(�ڎD�!������k���\��C7����f�����,�i��̵]<+-)��͛���BH�8w�ެ�ח���J�޵ݽ�t�Ac�µ=��ƥ�y�3ؿ���2��
�]9t�.p�m�ww�ٴѹI܃�rN�^9ͳ�.l}��M�� �B!����o(���(�+*��&��Z;S^	��&w?��\�%?~O��3���MAH6�mG��.}uRB!����{���ĺ�k���o@HD?E��.�9���y�]�vt>0��X����ٵ�=�%:ࡁA�.jƝ�i��Pஐť�-�va0g�_"����V�T�`mV��6>� ׁtVM��UX�pa╗k{\�l=Où���]�����;��C�ni�G=2���k�����<]��u��k�f��n-a�Kvn{��������c�����&'019�,O[��]�%�ȵk{Z��4�P�Ov����@�q��A��?�3����ׅ�0�x� �n��rR%WK�V���K�M�I5 �B!�������d����qc9�8V����X��Su�
E�tG�	��Y**`Y�
�K�cay�]�
B!����_⹝;�t�<x�	E$+׬��Ϯ�y�D�F�s��]�m^c!�9��h���֒���+?���ƺ(��nVP������S��s��t`p|Y���2w�A*#�Z���f���_�ڵk jY�q���ߵ]s��;���;c��칶�c5�vm���]�ʹk{"�ϵ�-�w���m~�s8r�0&&&@!$����{�����/���}rQ�"�,��{�!㱅��&v�Ǻ}��� Fu�����!�u�ʫA��1x\/��E��;����Ace����@!�B	F�D��\�<��˾J���;�I~Y�P0�L��e�/}��Q��vq���:�-]�cG��%��\p��9����12:��~*5IjDf��u�v�
�:��?��?���B=o����X��Bg�ڜL���=$��3�Z���wEll,��ؘ{�A�A����t���ͅ�21s����Q�4^RхA-KW,â�Z_�v�.�*���)�����-�gߵ�v<2��,=��(2��E��f��C�[\�5��C���m�l۴ϝ��� !����i|��x���
�:H"�k{�D��(�WZV�_~I�5�����{�x�B��ۼ���s#R��܍�4�
j^KFl�֋��	8t�B!������zQ^^.u}�2�*J���X���·�ub�Y>1Z��A�xя"w��Ҳ2��YB�P�^�|f>��	!�䎃���;�ctl��bM�Z|}�:&id����nttt��^��|`&���]��c�&���]���7������nT�Uax�ZհPஈ��S����`r ��E�����Rŷy�[�(g������C�@�Ҿy�[ܞ����8��947]�e_o�{S��[l��"H��u�A��pme�˗���C<~��Br���0؏��*:�'JC܋e���c��X��gBp,������8~��r��1������N]��
�ۼ�L��Í�ZH䞘\��
����U�@!�B!����o�_5ʚ\�c��� �v/�, ��ݗ|�E��Fc,��Y��Ŕ/�Ԉ��+/}��}��-!��q�=��~|���c�ჼ�����b������uu9rD�!�=��X�P�1��c���c꠫?M�d�����;�Q:9`.3t��s����U��KǺ%N!@�&�ҥK�w��:����d/̩k�=6�k�D�n��<��қE�b��2�hx��)��k��m�]�5��XX^�Kg΃B�:?z������U�����ڞ��wx�y���4ڔ�Xk[+T`���q�����t��������2��׍!�|���KZ����*�{��c��m)�9�O!�BIA-�0�BT0c�p�v�>�$���ܝ*�e����ٳ �����ׁ� q�w���@�BT011��'O���_��3 $k7�Ǎ/����4�>��XUUU���v~/�>f�=q�縴�2�;�*r7&�['�k�O��џ��R����a�'���RC}=�%�	�\�ܽt��=.{����P�'���h��`�̳a�f�E�\��%9��v[,��z�f���p�>$��QH�y�㊛�k����0>W��Ƀ���������lZ��!�����+XҲ�e�7����ӵ]��`��ڕ���v���';033�C�n��B�t�e�T5��A]�+�I=�*mcc�X���.&[	!�B!�Db}�сni<�1��oc�1�2����Jn�/~������Q�ʵkPV�U�Hj6�߀�7�E?!��C� ���lX��o|B�(�����m���M5����y����yot�~�Q�>4��Ț�-[�����[����Oc�/	�
x�9���vG|��3@2�̠U��{?���L������-˗�_�Ե�^&��pmw��5i��k��===�v-�k�~8~���2�k���W��$â�k���۞�����!������/~�K<z����场��>�>s-"�G�}�X���E���a�F\��9�.^��G�����3�0���m��'OZ:��Wߺȱܠu����{����)\�!�B!�x����c(/����c���T^��u�w�0W��lݝc,���� 456�<R��oRG!���7����P_���� ďu�S��?:v�.p���*l�s�3��˱��]���l%hy�ݥ�D02<���b��1V(pW@K�(Ɔ�]\IrKR}��:g��禘� �l�O�>��<*++A�P�ؠ�ӆ��tޔU���k��c�ص]���U�+.�k��=�gQ��|����[����ܵ��n�v�ٖq������BH� ��}�!���?��G�΍.iN]���fKD8��]ۃ��˻)pW�p�?p� ~����B�}Iz�A*�>���]��`W�����ޫ@!�B!^�����D�՟c�e&��}'�ܡC�n�c!۹���=��ܿ�.]�{�B�j���j!�C|G�m،O�}B!�C�ɓx�7q��1LpE�C��4/i�㇝ j����n444����dB�1b��4�C����G��n]�9�)�E��������N/H(pW�h_ a������J��
�}���/���l
��l$��Hq����>�ʵ��!���v���õ]"D����\̵ۡ��䱻]���/�P� >|B!����0:N���v��ӄ5q���{�ҵ=xl����+�t�2<�wDN��_�>�x۽���`��Z��>w_[�ܠ�@�1X5�׃���Nz�xA!�B���M`&�Z?c,�jSAͱle-�3r�~�����W��]�� �q�z���qh?Wi'��|C�O>x�|�U|z��c��v
�bc�򗿜�X�9VPc,_m�Ĩ:̣ñ�+@�C�{�i��`hp@_fй�� ����b�nq��!vW׌���Ln��3�P�� �ѣGAԱz�Z]���Kݿ��黶;��Brdյ������kΥU4���ˆk�����ϊ��c.�DS]=��B!��ݻw��e1�����u\ܞ�k��a>���Up,6�}�5���/��������>�<��e�<c�I��N����^6� �נU�������>���B!�⦢�C��()-�:�K��i�e:��_��+Ih��v^�sn04�Rˢ�Z,��$�w�¹�g111B!����8._���}g/�!^�,[��j��������=����O���g���K��}w��l��OQ\�SL����1v�ȗ�%œ_���{�A+.�v� U|[�6�%g��g���ӧ ���>~�?ϕk{�ܚ:6���{���µ]3�����0˲��.��uo�������A!$�9{�,����(-)��d<���{�{�l���!n/t��0�Yrmw�nܼ�,܃��!��3==�O�����uW�M�u !��l�)t*n7K��j-!�B!�8��T��B8�iǸ�+<sp�jݥZnЯ�Ν;�v��:�lh!~�]�O=Aww7!��/O?Fcc#V�\���n�/V�_�Kg8B�ΝÓ'O��ܬ�V�Ξ�Xn�e_1ͽ�Zʼ�E�.&lnj*ƕGS ���=�,҆0������E�*�[\7� �񭵖ƙ���P�:::B�d�e�+P]S��s��.���n��=���"K���z��K��N�x@�v�_nѺ,\ۍ?a]�m���69�q�3�pp�~]�E!�0������/~�{��k�G�<.����\���⋋#x��p`ߧ j8q�.p7(�z����������?@�\%���d�z�1�k@=!�B!�ɒ��ޑ 9C�r��֜��,K�3�kn0SBw�^(V&j(+/����.�QW[��E��8q�B�k��W_{O�{�?�Bd��^�k��bb|$�LNN���w�y�`��Y1�
l�%�oK܃�#����)\	
�9DӢ��1O� K&� EfR=���R��z�,No�ʏ|qf0��:�nhϝk�ԉ�ܷT��ڵc�Q��Fyn\۽�SV����ڪص�_ ,_��n���� !�"	x��|��W���q�<}��0�9�ӵ]���۟{Gb�X�ϟǣG�����3W��M��3He�c;����=���@��&<�$NB!�B���w"�#ghwp���}����G��DC����|�;�����k�~4!2�ul׶طg/!�G��o��}GҀ�H��m�*|}�:�N�<�܃�_B�pu���ːǵ��7���&�Nw��jAVf+��j@�A�{io(���8��+R8�[Ov#����z�⽐j��B��2��T�/^�ÇA�P]S���by���ڦ	�ø���oE����rm�8�;�i���k�Ȳ?� =�����)��ĕ���aQ-��2D�R��e�:�?@u}��z>���E��*���=h\��JlںW.\�=bb�Hڿ��#T�Lݚ~�'�t�}�[�0�,+�M<O��`�R���A��!B!�BH�����QVVp�gs�&]�ٹU�U��]�]1�|������K�P�8wW�[B���/���GBH�133�S';����p��9"c��u��ŗ��W��ӧ��ۋ��:�u&rx*�~8M��ew���}hw?�����j�&YC���.[��q��A��=�����Lw$� ��%.�R�V��ևI��T93ttt��Q!k6��N�"�B\@�n�C���":w�:�k��#9$qR�vg=鸶'�е��[k+��eµ�-�w�E۷o�BB)p�����ܣC�;�vyd���g�����+6���θ�v��]!'N���A(�A+w�#����C���=�du�r����X�e �B!��-���I_Мab��)Μ|kN�5^��P���C;s!7�W��cǸҜB��.GyE9����]��100 B!�G__�c��K����� �ɂ�J,^�D7P#�gllL7���O~�W9����]F���Ksk�s�&X����tpO�7L����M��7	�
�sH�t?F-.n���.^KZ$���vr��`&�4^<?z�(����u�J���� �+�vHE���.�;�|��]o�!��ˤk�S�n��̵]r�b���M��q��ELN�B
���AUe��$Ǯ�i�3�ڞ��|D��k�]۝��[W���	]����3g�d܍�U�V2'���@U��O�.{]�����{����c�Z��B!�B�QW<���9CS�n:�Y'�5��rp�c��O!�S!&�u�n�{;�SQ^��e+ph�B)\�~v?|��<~������C��	�{
��ܖ�1�s�碤s�!rO��S�bELc얲QP�~J9����Eq�8��e�*Ѐ����r&�-��Q9`�ξ�^��;w�u�*��%�
�k{n���횵6��Y��[ږ����k;q�����`z|
���!���gddCCCh���Ӟ����rmϥ�<h�k�W쮗^�G��H��'����?�K�z&�vbݬE����N���{����B�>:�����; !�B!$���S߾�s2m2i�tp/
էI�$��jnЯ����ϟQCuM5��@��ﾰ�!������#X�d)�!�+�bxp$�����WUU��=�7�}e���p�����eyC�?o����� �
�s�Ʀb̌Π��18�y/Q`�������Dŷks>,3��}	��c$s�.6ѵq����:��}HE��x���6y��]���tc���5�µ�8f� �&n�����n;N�k�f��~F��C\�6�]��� �B�O�>���8JKKuA�A�\ۥ��tmV��}�XU��N�l݂O�����8H��UB��d�Z��`5��TԼ���`��U���A��bU������B!�B�ʺb������ܞ�Ni���ܽ]�:��E�2
-7���۸�-��ׁ[6l��W>���B�����ʲ�_�.���+�d��5�z�2H��uBO��of5痩��i��m�wHc,i[��Z����� W5���4�?����1=.wr�<�mU^.>�p�X���� ���u��15,��E}�1��*�������d��0��y��n��S��)"O�3+�vs_.Q|"*�<.�k;$e���'j����[���|B!s�O?����]��|�s����У�tE����#nψk{��\��[��l}vΝ>�{:::R�1�Q(�V�y�T�8�/7C��+s����]]U��Jm$��2B!�B�� [�#7��7�2�$a�mX�D���`.���E���������@��ښE�,-��@!d���ߏ��ZTWUc`p �Xi[��.�����#�����I�c��.��Ԙ�m�7�c�9B��7�)�9�=���AR@�{����d��r�0��b|1S�.h	;+se����۷q��5�oڐxfum���S0���2d�v�ݽO?�[���C��9��"xM�ڮ7��ڞ����d��ɏ�T�k�H�qI��n�}<,�k���˖,��{���!������4<����u=ql.X.�ϥ�����
�}�
�1::�S�N�?�AN��a�3Y���A��uҨ�=���D/q�&���ղ�B!�R��`4	�3�����Ͻ�.2dY��PyC��3���g�p\B+V�����Xמ�?�}{��B����x�7���A �ki�rܻu$��`�҂XYLP8+8�ۗ��6�[֟���l��L�|]�#ԗ�������-���}�̅A���pg�8ù��E�:�/���{|���=I��r�d�pa��J�J���-����]��h�9�'��b�]����Ԯ��mq]ۭm���g��n���n������ڞ���w�]�%m/))AK}#��� !��e�<y���Ge���$J�����YsmO������_�k�3nqK�._��������w'��
ZO<D3�UK�X�p���)n���	�Ep���B!�2ߙ�N���c9Bc�碐��3yo4w�$�s�~�¥p$9VErͪuk@����z	�;N1�O!s��}���z�9��x�XY�n-��E�p���91�R�t*c,3.x?;��u�߃���1��E�?����%��Fyy�t�JvBk���e������_ZǈT|����R̞�z�ЅA+V�BIi	��v���H{��C&X���!n��_�OO�6�B�`��k9pm7��rm7���gp��AB���8~����1<2,�N���vmO'��];)pW�����/��/(.���@Sf���[���T�����ܽ�����X@$A�"��@!�B�ǈ��b�p��3�c%�&�W{v��*�xy�6Zn�/� j�k�Ǣ:
8��%--���Eoo/!��]����r|M�x��467�zQ��Ar��3wٶ�d���򑜈�9�~�S7<<8�������Z=�h�D��7k�"dO&ӋBX���`b��O�X�����9��S��u�������ȵ�C�̵]V��8�vmw��)���,�����cȺk�}kC]�߹��B���ߎÇ�ŗw�Q�cK�4�c�H�wV���;VO����k���6���155�[?~��W�b۶m3�4�}şG��W��#��WK�#nQ��2������.!�B!d��^��:D�~Y�m�e`�Zͳd9�B��m����܉�֬!Vĵh��t�>B��\8?|�M|z�W� 6ZW��Ջ�Arϱc��?�)�G��z&����XN�v-�O��׋\ۼ������K������!�XE��*���<�U����Uk�)��~�j6��:u
��� �G̮Nq,bl�k���{yP�v#6��=jJ���ܸ��"x�{=�eڵ�������5mi�btp�B��=�`� ������y���.���-��xY�oYy6=�W.^�-��ELwٶ�hJ���V6P%��8��_7��[��2p5=,�Ț@!�B�����c���_��fX����/J�nM
��;9�V����v��e}������� �ʋ�=���N�B��@w�>s;�ن�W�"&��W����03C�o��}�6nܸ�u��e,��9�P�X��C����Z��L�n�6�	]k�7�gM�bt���}A>c#!b��C�-�cWI�u�j6��g��am{{�Ea�ʵ=�I���x�>�wm��%q�rm��އ�]���{���z�ҥ8�!d^r��A������%_E��(�^���;��m�N��"�[������|h�|=�{_�r����T�"��D���[c�V#��h���sp�B!�����H�+��3�:¹����=˰�]I�Թ�B��m;�<�X�b9JJ��1������8���@!d���ݍ�PS]���~"(�(G�t� �[D��̙3��]�mn�M�Mf����n�O�7L�����T����qq���,����(/��]n��k.3h[rPsX��pc�q��Q=���z�2�B�.�Be{n�6¥@<T՟�c�[Uu�>yj�O222���N��s�%n�z�L�n)��NNOIE�1��6!�k/��^624��;��l�v�L.��3<8��%mu�[�ڃ~L��va�B<�|�z������1���(�[8��ttT�(����$*�]\o�o�����cW]�������������=�8�T�?�֊��|�޾����m�J�x�9M��� z�{PV�>'��<�]$cn}�m����*�^������r��鍝�S!������p�z�.*���~/��%��c]KK��{�a�)�z\�[�U����U������c����� �B!��C�F�~�5o�y�ܭ��d�<�Ù3ķ��W��T��
��h[��XY������B�#';�Ə���C�A�AۚU�+B�����-��?�k�2�rN47��~�`K����C�}XTр�QcyA�{�YU3�'bqy3OV�lk�������ݍ�ĺ�d�X�m�}�?~��K��U���'�u7-nƂ��1V\�]\��{;��Qص]v������������!�����.DF���f=�����r�����>���Y%�~� Y��&����U�m_���_�^����*e�Kq�UU���MNN*=���Re"o�B[Q�8n����[u��^���.�s��{�$���_v�b���M1�N��.¸�K�SS�(-+Eł
�}z�7���Op켏{y�wVK�k����Ů���y�]f�����$�������o��u�x�<2��eg�t�DY�DYGG~�����@S��1�J�C��#����S������'�p!�B!����B��_�sr��d;ۜ��o���(�ܠ_�Çq��]=O!C����VF��&�g�Y]�dp��&�|���U6�2<8������q������7��=59��ё�c,�u/nlҍ:��ef���~ܾ}[I��H�����J�Wy���D��7*�]\g��OLL(�0v�u�2dS�ً���
�*��w�?�_����x�+ku�����]���*��W�;/Py�1:<���^�����5���Q&Ӯ_�cT!�s��W��������?׍�jk�N�\\�����ͱfk�e����iIM�|���=���Р��=�Q�2U��8��35\�Q�e�
ݓX��HY�K!X	N�>��$za�D�@t�Ŀ����V6�^վN��01��ş�']��]�8��K�l]��5�ㄫ��F�Q6��Bq��\��.u9�J��g]�aQ]]��Q�8��sm7%�	�{R]g6�ɣN��׹c�a�}[�dmw���m�ܾ׮|��VVV*�����j%u��1h��~q#�5h�����c����PU��cW]��]�`���W��c����^U�b�l�ʖ����q?��_�����2�ۼ�"tKaoy�~�ײdI8��4���?�޼��-�������o��������Bs�~/�!l7b��\͋'�<�m�v��"Μ<�tQyo��{��.�� �N�a�)��r��������;���N�n�JtT,�� B!�B��CLx�&��	r�6I�<p�0Er0��-^�"�s�~�'N��E�^�qLU�3Ch�Jt��c߸u����ݛ��b�J��񃇨ZT��Ʊ��L�����z���x�Ҝ�+ηm�7�??�D[[T!Ė��y;qݭ��QR��cW]��'O����_�@屋q⮮.,�<x� �/VfΤ���B/��ب��|�ο��k8s�FFG�Rw_w�~��'������z���z�0�=��_��ŗi��{{чƧ�{���>q_"V���<�r�nc���n6�X���9C����yC���e"��"�
ܳ��`�Խ�s	s�����BPQ�\�:u*}�	���^��:�I����wmפ��Q�X-h=n7v��^����z��}?�D�.�vg�E�u�%�bN���N��\��|_ض/�\���	��L!��$��_ÊUm��띕�<e��� 6��ݷ� qY�ͦ`=�8y�<VL�\�f5n}���b�"&��H��B�8Д�z�ĸT4�@���Ⱦܠ��]��><4��M��O�B!�BH�����܋�},Μ����;,�ܠ_��s�@� �	1���.�t?!��Ǐ�{���Ǐ�A��U����>��/	��l[>�g�����:������qq���JͰ$⢉�Xj&��g�5�%������C�e}q�J����Q=���z������ ��u�J��m
��o�3x����2C�n)����p��sm�Ǝ�8M��!Z���[��ʵ�^��,�|n�}�ڮ�o�����Ï@!��%�֮[��/D�vqgnE�qmOI�]�5!M�z�XQT�n�{f�3�+@�4q��E���y*F�]=n��M�9K��ܓ+���|���o(�ɻ�B!�2��[P����x�P�<s�.c��
R�՞���,S����2E�� �o1ћ���&,T��,�/6�[�_~�\q�B��F�,p��-�[�_�n���u����-�=Zqq\N��9�L�!�R3����shC�+?'�;����Pʋal
D�Ydբ�I�/wl�T9��!�L>�vb�#�g2�Μ9Î�"V�l�!w��hy�LH���n��B��[�?�]�݂}{���n�h]�ׯ}��
w!��9�?~�֛���P��v��s��&�����u���˒��=���K�.�wٶB���4�%�V�GX���:�K�� !�B!�����nmZ�|��_�|�9C��$�z���_.�Ο?�����C�vbPZR���&��!��o��?xㇸy��DDg��6
���ݭ�mݺu����+���Y�cYs������ ���b\��]�Y��dc�6o����J]�Iz�,��P��\��{�CCS��8���^�v[��k����r���K�s��no�۵�k�(?�Mu�p�!�'������Eii)�'��Y�g޵=�"�|um��՝��7��W�����J�/)t��x,�U��y��k�s��r�ց*�C��Pl�t�#�B!d>�T>��ሴ� �����v+�����&��B��m�3i�E�!��+���K;w�tG!�'�;N��gw���� dy[+�^��{�1����]��Ps�nc������Jهv��f{��;��2�H�KL��
ܳH�Đԩ�ӅAs;1���\N��`���2`%ܢϞ�M�
Z׬��k�'S�n-s�г���ƻ��̵]Ҿl����ݽ��q��ז��8s�!�/�>�����yx߾a.��k�<�����^�鸶;c7?��
N]]]hjj�_���l��S�b�A�q�=&0<Ћ������B!�B�ҩAL}�ܡf�1�ΤyC,g�О�O�;�d�/��iC�	�$s,^��ee dQMF���!�)�+������@�9��T,�@��f<�|�[.\�������b3Ghbl2Ӆ�P9C�������E��h��r7�g���';��봗z�/�fhXN����^N�r��5W�u?�Ն�������=m�e}\�!�K�M.q:��\�]ù.x.\ۭ�5�E��fM�%������j���q���ѩi��p� B!ވe��q-��Ȉ�y:�����gA�J��`�����d՚�(+/����џd���)�;w?�я�&e��!yg%���x�V`���pf���������r��B!���9��@_�?q���cY��󆎜a�r#�|���c����|�� �g��V"xa�N|�w!�/Nu�����*�8B��;�G�ń���j����zߵ��1V���]9D��}r�7Vy�
ܳD{c	�#Q�I�� y��~�ۉ��%;�ˀ�ŋ�L��բfѢ�+�v] n/�J��p�>$�A]ۍz\��ʵ=�xoB nۋ-�.lw��;�O��R��������8�̆Mؿ�B!��t���Ż��pm+8�� q!bϵ}��vQOqq16lބ��/��+W��w'�ࠐo���l�xͶ
��@Ź��ʚ(nt�B!�2XU_���)����'����2ł{2��4P�s������½]L�&����K�-!+W����o�U�	!�/�1�4/_����t���m.�9���366��.�����Dp�6hW:���������`[���߱�Q�TE�98b��,��2v��Ig\H�\�8������Iy��|��ԀեK�@rOۚU0��LK�ε]*��	̽�c�,=�v�@�g��]e鸶Ǐ=*�<0���)i����zt>x���	B!A8u�$v<���v%����е]�����U���k�m~f�
8u�m@'_2�c��r���@�UE.w���dc��b5��B!�2�YU5�����_�����p�~���}$���!���l�|�2H�Y�b"Ŕ"�w�5fM�*����X�BR�����7ߠ���%/]���x.��w'����˷����2ǒ<���]���kk4t�8`�2KTFG0*I`���w�v��yXќ�����$se�J�jϝ;�{ZW�
��.uI7�,����0^'y�%�V���no��Y(��d�A�C /ڑ�v�h�C ��>��F�ڕ+����B	�Ç�\��$�'����H΄�<G��h����cκ���,VVϊ�V,�����0H�x��n޼��k�zƨv`�4�];�۵�����AE��1�zE=!�B!s���8�Nm��;��^1*�Ê�@+{yðd;?)��={$�,ok!�m}�/�ЂBHp�^��-6���/@�7�W�R� g���A�[��⢽�%Ϋ��1	]�
[S,�(��2a&[b��,19�﹤�|v��������(��.^drPʏlX	��������܄+%�s�v�gܵ]&��/��������m��ݝm7۰�u%>�u6ru!�2w8|�~�֛���1HA�v���ѵ�3>����Ѧg6�ܩ3 �C�{\�pk֬	5��O��t��V9�����f�8��P]ր�q�?B!�2��w%�}��\��R��&��K��-&t߿OQL�)+/CSK3������e���!��G�aӖ�().�����e��e�����$H��ꫯ��ى%K�x�D$G��Ѩ��;�<ٯw�}L�l������P��j;�g���FGFP^^�q!�;Nr���\7��\�_0Gi�ǕO�R\f0�X��*����Q�`�.�v��#����)�w����
o�h����*,w9�[��µ=�'x�]����{e�8}�6!������)*�+0:6RD�I<[��;;�]۝�o�@����������<�
���s�sP֗��rls8*9\ܭ�T�ފ��P�s88K!�B�\��T����.�t�<��\}�"W�$P��P�k�|��}���������cff$�,Y�\?g������ �B�r�dv�܁�s��g"������� �C��Ν;����'s&G�M�?5��)������?/��&�;���PRT�IvamP�����N�Ay�k6�yr�N�K�n�,����By�����%Δ�t���3SHn"sI769bø�����%����_�m�;��um�	ĳ��G�� �umO)6�o��S �Bf��c��w���{�\�º�;��vm[���rii�8��`�Z޺��I����)�	C��K
�d�A��h{$6�'��.�^��ec��B!�2�i�� �n�&Ib{cy=��/I;`� ��s�o�����I�Yֺd~S_W�������B	���f&�P]U�����˲+(pW�0w'��#̬1���,s>��ۖ��L��\��=��=> &�k(Ƶ'\��
�Y��l�E�U�GQ�/DJ���,��]'��چ��a\�z$���ա�:�<��k��L��̸�����k����n�k_Q�W\\������B�l�����;����C��:��rm��l9�#Lh�\ۣ��p�*�E�7n���@rG__�_��-[�d\؞��Z�*�se�U��i��KZ�b��i1�c!�B!s�%�Ә�;����˛����K�74���>N��a.ȶ�^�5�+���󍋛A�7�nڂ���!�2[Ν=�W���8
2iY���źI�b%,k.���A1�pu1�NsJc,٣Ȧ�i��V~��U3����Y�dz�K	x;1���6H���ra�Ǩ�R� /\���@rK�6��":w�!� 1��Z��5�2����"/���M׵QwY�\�]mפm����v��'=�c�mj_�3'��N!$}Μ9�w���.p���*�k{�����7�r9�|_pI&sߗʬ����Z�ny�d�J�H�{�Όg������qΝ��z�c[[�e��k�U][֒�U������ 	 � ��׍" &H"���'�tm�~��5�#���l�0���.)-���/���rJ2���4 �
Ύ�	w      ����1���5��V��M�:h��U�1w��Y��1�{�.�����s�[�1H/K��fk+2�<   �	�x��O�ss��{�Ԓ��h��*m>A :677icc��\����냜#���[}m]w���ۨ��ܡ�C�1�sQc����@������U�Q���l	�v�>f�>�A)պ������KmW�ڵ]��*;�ѹ���&��� ]����+*�v[K��;��j;K�>��S�Z��CL  �ش[Ϟn���4�W&յ�G�(�^���l�.]�L����1w�ܑ�G��FpA+G�C�������fpS��˥�Nfi�N      ��||�pm7�*c,�����Gq���+�'(�$�8���m��_�@ �|��w���v   ��՗_ҟ����/��������G�Gݼy�._�I�0�w����Cr�j��q#���ꬹk�ża����X@�0��Y�T�T,[�R;���g8�B�H��I��=(nܸA Z�f�i�����ۅ�B�p�!����vm']R�g8��k�u�<)�y)��y�qm�{um��W�;�$kV���H���   ��y���&p�,�n��X�k����۱}J]��=f�Yz���t�k��G	�n�M�Ȧg$#�,�)/ Q\��@��O/�d��'�2���      ����,��J4:Zt$�U}��M����e��Z�k�E�9�۷o��\>GK�+����2m�x��%   �c�m����"���&�NV��Z��FFAQ���_���<�y@�(��4�9����{۴��:��쏢������tR����si�y��GX�.Z�"f��w�Q�JA����7�|C Z.u�"	Ƶ]":���ڮS��=��i�]��:yI[����yj\�9�]j�ݶo�?�+P��L���   ��{��1�./���������P(������U�wo�����>��=b޽{G�=�k׮%F�V�L��*��W^|"�ZP�����2?R#      �p��\��(��ɸ�5r�FR�0���24�A��$c��^�ӗ_~I ZV��Q6�%�^>��1����/   ��믿�?��O�ۿ$�N�1���
m��$�?���t}�s��:1_��yV�vŜ�)v��3y��7���W�tc�C�f~�JՌ<P�tbp�0xsb0�ZeE�>+6-D�ѳva݇k�f^�6�v���*yK/�!���]��W���A�]�ڮwD�_�N����&    hX�����v�U���	�}?J���z���{<�k�ȅK)�˵�A4��ͭ[�Z���*��~�ٮ���pI�J�+�7� �����B���W�       ��b�F��1�,�����U��|��ܡ>@�A7>|Ho߾%-k�H/���i��S��  �����--/-ӛ�o�����!p������ܤ��{�Ǐ[��uC���=����}za�L;�g[Z���56p��H�jB�Ze�}qI���*I�J��GPJ�ݻw�Y�����.�;�����E��e�Q2\�e��"u��c?y���:ϐ\���s�����@Ф0Z���	�J%   ���~{�-�����~�LRO%BA���p�U~(�FFF�ҕ���ۇ��M����׎�8�I�c��Z*!X%�J!&(�A�����j� p     `8m���HfK��Rc,�C�z��Y�ۇ	��d�[���]������������-   As��M��_�������3Y_������7n���z�s}��ݍ~ukQ*'���w� v��]�f~.j����@�0�#����R�2�/r�p�NE��̆��B��F�i���ٵ�YF���\�me�g=;�S��pm���2�M�m�=���F��?�F���N   @X�������;ؗ�O�k;��cG>q�ޗ�ݷk��Vytm���!p��/��"�v��U��_��{�s�i�fF3��       �p���f}V.ҙ��ܡڵ���\�3L��U���D�����a���.ғ��   vϷ����VVi����Q���y��~G :�ܹC?����>�9B�u6%��KiPM.}|!_��)
����qs��@� sc:+��h��ف!�u��]�.e?��>�A)q]�Z�o���@�8���]\�5aC�p�������*�����$�#���|�rm7�U�ݵ���k� ʷ�ۤvm7ʊ�︣�C*��   ������\�cgo�,É�O��wmo��X7Z�v��W�#-�_���O��{�E��G��`�)���U2�H�@����$���{��rw      ����zB�¨ÙM9Vҷ�'o��k�Н=���	D��:�����KW����   �oݦ����{�a.��G�W_}e{�=�u�:�*a}k]w���-������?g�e�h�R>;G�:f,`@� Wg��9�8�nIm� �07��'�qu�Ş�$`Ÿ{�.��l6KK++�
a�Ñ�t����\��V��n�������by]&�'��ڮ�+]۹6���ѹ����k�y>
Q����ý  @$0���_3�tm�P��ޠ���u���iii�޾}K ����͛t�ʕH�I����x��,Xe����Un�*����^/!n     `�x>Kک&up�������=��:.yC~�0���A/_�$-��k���WޣG�%    l^>{N�����&������5���M�������n�k�>W���i�
v�/	�y>7���b��N������*�e�X�Fə�vso�.NE��!z�P�0xN��$v����s$�ϭ��T���2޵ݢ}�J���µ](s��5ތ���9���e}��;�Ѝ6��ٗk��}��]!�'�����n�`���U*   ��i��<5?G�GF�v����x��k�X��G� p��H��wPo+�]��N��_�q�nY �E��pp/��
      ��u�7�Upp���(� ��"�ża��C�0IW��c��7����)���$�N.�������   6L����'�����Y�ӓ�P���o��������煵�!
��~6׷�b���g�����l}�A�1aA�dT?��$Q-
�m�3� T�d�QO�r����u���'-�/�/��\�;bj��;�vN�m�͵]s��ޮ \��gb�Z}~�^]ۭ���O����   D�7_C�����]���%X�k�����{٣���W�_��	Dǭ[�(�z$�>v���Ry]d+1f�(�      �tF%n�qޙ���[����Y�Bخ@���u�~'�Y=�N ��.����  D���-��ӻ��ce�=y�@4�>3�bwٺ�ԃ�a�!t7���n�<��<�`�=�eƳY�J�t$�f�pJ�R�Y�r�n���V���۷	D��yn�A_���69�����K��5-b�v�y���.�]��&n玧rm7^��ۚu]    D�m�~C���+�P�pm��\��W�x�v��s�T���)�h`B���=���k����P���s�5��K��:	�UN��`389:�b~�J�      ��r$��w5����pM��T���FEzn'���s���^�{;  �H�q���c��_�+�����{԰��gnQP?}k�i���.�k���xs�
��`� �11��ӓc*FM�����S��r���wb�+j���y��-={��@tL�����D[�ΐ���l[�]�ퟑN�(]��N�s��vᵣ��;�g�n��F���W蛯�&    j~����O���>n+��*vI\�{�M�������X����W�֍���M7x�����X���un�8.K!X%۷l`����F��,k>gw���e���     FrDǇGT(ly@/b�L��rڵ��'�u=�upp�����/.H�SS����V   @�`�X��3��#�����f��\���7oR�T���g���i~嶎=o���2M�}lo�ϼ�d����!e�i��^��xo.KT��=N-(���e|��QGZ�	}�V̽?ZѲva�ŵ].��<#�3Q�-sm�
�%��g��zv%�Y�k��L�^(�.o=������vvsm��>96Ao޼!    j*�
��:y��E���6�*��v�{����@�!�o���Ö�}���y��b�ʪ�ra0�WR���%n���x�0?      ���y�3�&�e}ǒQ�=�tI��7�8�l�6�#��X^]i]� }��w?���&    j������1�귿!�.X�xay�޼�"����Ağ~�ib�a�i.�w������7�H���x��7�ժ�>��g{5J;���X�2�tDE7�v?Ir��~�,1�������V��ѣG�eem͗��.��	މ����J�tm��9�w����@�z+]ۅ���ڮ��a�����.�ӟk�f+�����[�tne��}��   ���կ~E�ӟ��W/�|ֽօk��vY�J��W��%�r��}iy�
a�k�3�|�{\���qc(f��=g	      0���5(Sq�ޔ�����_��;��<�@�0z��&H###T=�P�Z%    j؀ƑL��Uk�v�	�{t�>߃Z���h�Xe�v��\��]�k<�a�ͱZK�.N=ۣ��{@Ld*t&qa�%��1�~8$+Is]�e���w��&�XZ^�ܿ�?
�t�Y�k���BpI� \��7W`�uum'�c�ǵ���� ^�v�h��v���)v7��|X[^����s   �����z�)BUjأqm�R�&�v�drj�5����;�p�֭�4��	��z8p���-�l��A+bv٣����t��      |&�:�2Μ!g�e�7��)�~��.�c�^��"���U�T�Ax@��N~��ߡ����   �����/���|����5�t���J����=J(Q��?2�����_��g|�b���23�<�"[?��
����H%���
�8V�Z���0>>N��F���bb�������'&'���'����J��tG%�{�C��s:����U\��muy[�˩T*�
w����r@��c��
��޿}۶�׶��)_q鈴�fѻ�o���[.�9-�كG����ȓ���b�����666b96��b.l�8`�ξ?�r�988��/��f� �s����z���%�<w�Y;>>n}�����,Bq��0������WZ];GG'���k�}描�iow������n�����׿QU��Wi�����?��g�������I�c��7[��ޱl���y:;-)����>	�W�k�؀��ϟ��˗)i�j�i���d�'���O_���)�n��     �a [/9��]��r�^ך9C����X$�u�Dސ=�m˿����������*d�   ,9;5Cc,0�L��Pq�H%��!f�œ��q�W������wM�y�.�XBܠ�3�S����Ѳ�MuQ��xa�]��p\�$O��q
�ezA&nBp�\�%�k��㡗s��;��kJt�V/w���V��ާ>�f�S��˅��3݋�{�N�޶��KK�!� ��`~�\\��2����ߺM׿�qOm'�L�vѵ�lS�՝�7��O?q�ǥ��ɧ���?�ҥK��_����Y*���}��i���+L���K캋&P�p���������~�صq�{����ަ������K�����y����c9>�?ZXX�mpA����~�3z��R�noo�^o��k]�
CpmW����~M���O?��������G]��i�W�v&l�V*�~�|׺�{��i���}{��wR�$�I�^�u�Ν�g9)
a˸X�|�K�"v�"���׬83����      ���5�����`�s�B�6!��H�~��I���/_����݁4�byC�������Y�}��㾎ͮՃݽ�qB��������&���~{�^��%�Jg��[YZ�������cai6bF-����ۋ��)7gb�`�{7�<w�=�οR��r|f�=��L�0����!�g���o��Fǋ���#]_f�`���	g���;ψ�>�trJ#{�{�p�og��}�}��8������O�Ȼ����X_������ܢ���JX�[��i�`s�7$י�������ww�`���~�����$�[��Ī�lSߑI
t�u���#-���)��v��&�G-q��K���n����le�<�.�_gs�vv�8'ׅ�:�t��T}������u+����O�5�+��A�N����v�$/�s�0BǇG�   ������u�۷�*��Wq{�"�~�*E�rex_u�ܫ+{��Q0/����Y`X�D÷�~�P"2h���d�2����.V���7�%x��_�����     d&F2tvvJ�¨ҽ��b�7��V%һ%=T	�8�l�v����%<3�&q����'�&1;����O��{�)�l��əi�˨��c���{��\:���ZY_�ݿ�����������l�̙�w���t,�O�{���[���h4�A��L̜��|����&����6�{��=��e�(�~o�ʰ����~�/�$]���ۺg&Jq��|���~������D8�X�����k����Y�gtt��IX�����7oҏ���ԃF���tx.��_�_��N�(���Z�ӆ����,ig�R�pbp��_�H7q|p������K�?�o�[aB���y���S�����z|G���ќ\�����\ŵ��;��~��׵����l�̶K���������+   ���{�飏�c
�u��]R�k{�����O��݇`ݯk;O~$Ok����]F������_�����+c`hkQ��O����sA�\Ly�
     �!��l���j�;���`$���E�~���$�(o���>|H :ص���L ]\X[��O7   H
L伲�L�߾!��ϭ���{��QK����:��|?�S(7�r���>�[�0c�
�FC��39z�[�4�{ ,�5/����&f'م�t��	����v'ɑ�<x@ :V��Z�uQ4�ݵ�+ٵ�*K�k;;�����ǵ��.��C|O���v�l����	   H
�w��`���lkZGgYQ�\�Uu�ڮ��ӕ�߃�=B���9�
�� B
�q�;��K+X�}��՟��� ��]��ևP      ���8Q�"IP�^�}M����n%)��Z�@m����<�;�� =\����?��   ��p��]�џ��)c�Xl9�����N3IWA�=���m����1@��K<7I�x�R��0��RY��V&�� �p!���F�I}A���?B����g]�\��=b�W��7K�lI�V�ڶ�%�Bpm�I�F.1D���;��Ѻ]D�>��@�o��smw�ݕ�S�ŅEz��	   I㷟��~��?��/�BkĚ����zw�v���k����k�6��ɓ't���X�M`�.�.x������28��\�����Ϛ��       ��2��PYq��g��D�����[�H� ��	·�~K :�ޞ:
#*��7{  �t�~��F��Uk�v9N�~��`���Z6�m�N���������};�ny���"���s�|�l�Ni� ��N�#)$�v��])d�vl�[�j����8������trrB :�W�h�Kx̮���	bpI��W��ծ�z]ۮq��}����v�\Ϗ�~���/��   ��qxxh��k{�mRW���G����γ���
�����G��0���k�"�{[4�0n�>ޏ��[_����      6�z��.�X�����FWlyC�[�3�<�<{��vvvD����t��w>��7n   �4n~s�>����~���}t�Q���+z��5������仺�v�A�.�Zy?�_�_�=.3�*P���= �g�����<\�F��{8J�`�8�c�A&�����)���ܜ]��~D�my�].��zе]V�һ;����.�D)��e�trt��  ���f�_^���ǺH]���'\ۻ�����rt��:��xF X�KF\�a��bǥ�!`%�M���1 	T�J%�-fh��       �`R-[����ۭ���!u��G�7t#���G�D��-.H�ctttD   @���ۣߙ�&�.0�2RX���Çt�ܹ�ЃA<.{.�{�}n���=oH�~~/9�F�� p}1Y�P�D�¨�sV��y��6�뼻�>ѮX�"��
~����A :Vέ��iF��R��,P��N;,wQ��vm�� �k��
ܵ��&��^x����+��W�}N   @R�}�����M�K������z���um燐W�vq�/]��=Bz$�]�?�н�W���u��ޏ7�I�������Y�     P&FX��7s�lI�]s�N����`�����SD�0Zf��(��H�VWi��   �ʻ�oiq~��w�H�B��f��p��@4����&�ܢ����j��7���F<���r�y��8m�{�\���r�(!9-wR�3�C�ca�1_G0�%)�~���cyu���S୓�ƞl�vN
�ѵ��_O��ƶѹ��$>�4� ���x�
����'    ��{ȓ�c�f�T��S�ڮ��k;+����.k�������ݻ�h4Z�3F�"t���e����b]Y�ݳ�]�b��X��T      8g2De�֌���<�=oh�5��$�y���pp��e��kWާ��/   H*�oݦ��G�����})�����ci���_u۷���~�V|Q=@]�74���z��w�昵��L����(�@��'�E�2g��v���.X�*X%�u��v'9����9+t;.��	��ݻG :�W�5�F�\�ۓP�k��пk�D��E��j�Y�h�M��l�_�v���ֱ����E��    ������O~����զ�<M��A�߫�=.�v�peu���g�k>;;;���I.\�k?�����[�N�ʵo�$-��/V	q�n4Si�3K      ��ce�(S�8���.$�ct�
K�,¼ar��9��cai�@z`n��r9��;   ��7�4c,������A�k���
^�.�{;�{�*�L&#5��d4Z� z�K��>��T�"��������*��#2%����W^�xA��)��FL.��مYA�ݫk�U.�׵�o[��X i{�v*]ۉ���v��wm7�.�[�����A   @���ۣ������ۄk���ǣ��������iu�m�xI |�ߍ͞u�����н�M�ݶU��ߺ؏Q#���מ�,��=�(7�5F      ��c*[��b@�J�Nʁ�Z��!��G��k{_�~�Z@4�����ӏ>��7n   �tn5�>��ݺw�@:�}i�lll���>���v�;�W���uD��(u���r}xO�wS�������3 p�|�LUc$���5�\�|��;N��8�$�.�Ӧ`�x�,�,S6c�j�rmw:����g쇀<:���.i�]��k�M��9�n�;��rm'��]�vM5�|�u���c�Ѭ��\Q  /�=�əI:<:�L��R[���z~�&յ�������\�t�y��i(�MJ��ؕ�R5{�]��|^pue�/��)A�     �`�m�)���Ͱ��9��P���t�vٺ���#o!ӳ3-Go��'�����   ���f�����.��P+�����Z��2���?��XD�n�[��c��˻�;�󆤈���eTg3?�PZ���OՒ}zq�E�-P�p�a߾{8*�	�?N :VVW�c�M�]ۉT"x�_�f:�;���.m�\��ݵ�lm��K�v�#��dmĵ]����6���:��_�[7n   0(ܼy����˖��Q��֕{�]a��˵�����[�[[#�=��'E��q�q)#`��������������ͥtrBYm��z�@      @4*%3O�O+޵O��d}�ֳ.yCUB�%��W�� ��d����Ez��   {;;4=5M�������G3�b�^��"{.�j�E�ۋ}z����z�+��~F���9+��ܭ�M3h\��Hp;.lV%?�Z�낌�����E��ڮ~�t-b�vG[a{H��r��؆(\�ݏe������m   6R�Z�t��k�TD�"�v��vym��v~�������ȎW�ʀױ���µ(���7���q�%.� yv��S9zyP'      �`qvzB�\�S�Ж7�&�53?��uI��7L�@y�hYX\$��]��~��&   `P�}�6��������������x�@4<y"��"P�|�P�R�W���k�@6`�R:i�a��
�}�8��Z�J�Q��*Ub[��e!��[$!������-�bj��D���QF�z�M��Y*Z���{pm��%�]�]�n����9�˵]R��&����G������  O����"���I�õ]Z�����˵��M585=E����ٳgtxxH��ӭ׃���q���f�4e}�â]��݉�-���     0Zy�Z����G�vU�[���@uސl���&!o�P�<�ava�@z�6�H�u�'   �J�
�<��0��@ :�`���"C���l�?+���\�^��۫��,�X*�hb$CǕ�����d�����R�0��2:"�.�p���u���Ar]�� �gfh�P��ӵ�#��T��=��i�߮�܏k�ޏk������pm���{-m�b�3��-sls��y�s�6   �ƽ���?~�!m<۰�G���,�O�]���jT��Ы��v����t�&�[���3�������	��lɷ7��;/5s����jv
���zݝ2�e���       ���T�޾d�����������$�����ڦ��c��� ��Q�'������-   ���=������]����4�G�T�T	��Ç�I:z�$
ԃ6�jI���˩���5s��$[a���hm:C�ә;�������T2��u���]b�cX�)�gA�j?HQ���Lm15	�i"C���:��pkm�Yd���(k�`�����W�����g�͵����\�e?{��G�i{{�   �A��՚i�0��pm�ϵ]��z�����˖�]�p��ۅ�f��gQ6���B*T�eX�7C      ��a���k�9��'�ż�8x�y�a��&�7,���a~�i����_��   w�ܡ?����	f�I�4;?Oo�^6��W�����}�g�r�����������zM��*N�q�2�4F��	�}0��SU�𸋋�T�t������#`�6>D͠9�3��".��4����ݵ]�Փ��w�	e��U�����f\!���m�S .�Ώk�c_Q��P{Y��]�$�A�|�N��   T?~BS�S�z�u߂u�u�9���ۧ��c�umW�Ӈ��Gq���*����܌��Q��)�\X��b���su:Z�K��E      �\��}�gQ�������C�P�7�Ǡ�ٺ/^ o!s��҃��l1c   `�`���,$�ibn��0�/]�40�ޏk7�2��BT�o����>�y��\z���m�#T����5P%�P�\�m���"�@,Kb����D��Ғ��[��nWP��|n�K�ڮs۵7�����,>���\��O�ц~]�e�v�����t�"���   ��������O<�ǵ�O��]��{�7"<�v���>���K��f�d���O�J��]��x����_��/��Te2��^)�      #�2�$��]�>�<�yC��}��q�N3s������s��%>_   ��w�hzj�a��
0�P���KNnQ�S''���I5��ݖ;���k��_
��9�R�t�uPT����`�i���%�ݮ�pe���3<H�l��l.G3�ӝWy����������ؕ�f=��Ei��Vc���)����k��NB�*v��� �:�NSܮ�������drtu�e��f�+����   �J�ѠZ�ҵ^8��5�µ=�=�W]ZY�-$�#�ɓ'�׃��}{��]Ӭ��B=Мwb 3P%� �.g����Y��       H<z��I��o�ж�|��yP��ٳg��]s������G���?   0�ܻ{�Ο;Gw�}@`�a� :�LZ2�#P�︖�O��X���m�~��]>P��.[;k�e���}P*7/$�*2.T�]��}v�@)�Q�6KZ��WDa�ťE�d�d(�"o�;��������!��J�v�#ng�I����v�\�.��mm��i����k�}��Nz��3v*w���I���#tt�Q�   ��_����r}8������ܫ+{��k�������k�G��ũ���u����2T�:�A��]�H� d{6;��D�^a�      6P��U"�9C�AL�LS~$O %4���   0�T�U�e!�L��Q�����cᣚ��W��[�4Iʚ�+���)� x7����R9;!܁/f�Y��+T,���[�@V��^7�sJ�#���	�#d~a��$0�v��,�ε�cۉ�#k;�//��f�mD�fەu�cyqm�vJ���x�\�H_}�9   �Kj����r��+w�nR\�E��	D�`�'�|K)L�v�:1.Վ5��!�Px!�!T1�+|}���d��dw      ��b�*�*�9�#:���i��
�ffn�@:8���2   ���=����:�w�
��m�hx��!�j5���`�(P���jQ�7S,��-. ۟�C,�JT�iT�����Y�ʐv�=0e<��0
C6bC�����0	�^a�v&� �0�0'\_N9Q���Q �	�Cqm��k;/.w�������~;E�����   0�{�Z��(󺭼\Z걞�nH���� ����b3��x��yK�"����1�gF�����oT��,b@,����     ���>�E��Ǿ�8.�m�\.���y����K�闿�G   ��Ϟ�'��)mla6�4037K/6����C��ڢ.���A�-�D�$�[u�}{��\�E�.�X���n���=2W�)S񗜶9�u�#��1/R늷���oP(��,P�񁝹���3��g�v�5qs�L�-���xsm'y�I��h�F1��s;��ڮُ���d2tV:%   `X��ݥ+^��f��+pm�����%n�Qp???O�l��u8\G��f8�d97؅�f_��������pE�C��H�       ���(�f���#o��q�@l���	�@:�kj40�  ���~ϲZ�@:��jt���Y����!Pb߬���4��A隽o���d2�L=ޥ��{�L�4;u�G�g���Q�ū�h8V�� ��#��ׯ	D=O�L�J�ݛk���[7kr"m�����zDζk��л�m����7A�v���u��A�_�?���
=z��   �a�իW��s��C�����[�
���˫�>������}��@���a�+D���L��bԕ��{�X�ZG�"��:��l�       �g"_��Ϝ!����˗�czf���3?7G��m   0,���hrb����7�GK?�X��[��c�}p�/���u��@w2��~̱24�O� T�{�@U�h������ �vq�#5��L�;6p��
F��o6��6�`&��z�2�s�3��,�L� ����ڮn�L��ŵ�!n��.���bqm����߾�7   ��Z�Fz���jx����um�S7�v�zn���������{D-H�s�$����|��׉{.]2����+�;      ������n}�v!�}웙�h�����H���������g�   0,<�ؠ��O�_n
��4Z,�Y�D |T:�$��z۷ l�N�]��K��{��O��N�7��V'�p�?�@��#9�JU��$�@[�����~����i��aN+�����K��Ե]!�����Z��&'�õ��v��v�ޝoCԮ���=Q����Q�Z��   ���c�f�T���ٵ]�PO��@\�����[,���-�A |666�ڼwi��]���R����vW��U������~�/0��V=k�N       �d����GbyC op�L����e   ��R�D�㈳����Y�z	�{�2�8.�{/������~"��u��]�.�sČ�
�6 p��vfKB��u��dImQȫ�0�D��}��������?N ��;�:Rn�k�W�s�ۮ�s/�k�ŵ�&��ӵ�s��bq�2�v"i�bwj��]������ŵ]<�񾍏��λ   ��{w��ǿ�)m�~m+ϵ]R
�vO�Tu��KK��������imm����s��$,�H�Vq��`�����rvz�|��f�      $�z��U��=oh�)�7�o6�ߋ/D������T+   ��ѠL&C��#nff��3=E�q�y�$�_�z\�X��5�����(h7�|���Yy�D��x�rVrMD3D76���l�N<�2!`�g�F]���-1��v�*`�vC�M�2޵�] ޏk�&�N�v��P~��]۹#+�Wtm�&n�ʺ����[�_�˿   0l�)��h����~]��ԍڵ�K=U]u[=��#���-�3A0w�s��%^�ľm"waq��U��X�ʥ���h_X�}����S�     H:,o�D3*�5����߼yC ����^�B�>"   `�x�t�ί�ӳ0Vvf0032؀㓓����Z7I��^���%�vu��9K�)tw���K��f~����{����T�tq���m\r^�<bB��gs���g_�̍D���\(��ium7��RGP�+�k�̧k�Cl���L�f   F*g�t�um�ֶ�\�=�S���v�C=U�z0R(����ku����n�0���7+s\���<���o܌��z� >C+�     �t�G4�T*T,�[�7v�,o��ؙ���=�..Ӄ�w   6�={F?�� pO�s3��Z�ҫW��>��_/�64�|ܾ����f=���%�����N)��TO�������d���P]`D$<�A*�%�y��2IN����ׄ0�̈́A����&�㻝���8e�j�"!���7�v���7�"uQ��pm�0���ŵ�^o��j��m_���|t��S��"u[�I��aS��5�p���"��õ��@V���4O����~D'k�ݛǋ���{��繳ABq}���޳c�}�����ٱ�����7��\�� ���8���Ϩ01FG��B�d[*�E}����תUr#�v�_s�۷k����F�}��Jɵ]dna�޽y�}�2�nWX�x�sn�"͊^�ZdbT�D)�h�[��x>;
�      I�L���{��yC!�����}�~��@4
-�H4  `Ha��ls8 x�'&(��6
X�mss�%pw����_��҄��κ�Z���-oHB<������4����t���Kc�N��g��"�E<��'��������靤����[�A���ߧW��,���&�q;���)�x��V&
��m�ʚ�b޵�x���KOُ!ݝD�-)pEl��Q[�vx�O�9��q<�Q�|!�M�T��٥G�;���qzF�ǖH�0M�λzx�MNNѷ7����E�������v3y||�=L�W.�[#��������M��={�Y�5��
�<�����󑑑�oN�y��c�yq�γc��I��e�io߾�>��v�w�+}|�~J����1o߼�k�~���������޾�K0���.��P�^�}vo�g����U�0R��ޞ��U�.��}xTΎ��'����bF?߶�>�.��[&�po      �����'ޝ��{�yCqP,�ۭ�c���E���J\1T�s�������Ўͮ���i��p����;0f�����Yl�^�T�����O�OЍ������Ȏ��QO��,�:�qǔ%��]��}��g�+���B�y�,R*�b;�ql����8�{v���q�ާ�3��޹}�ʧ���#*���g���]L�g�,�7����ǚ���z�;/�{{C�������e�2x�E�9��p�����{i+�Ms,� yQ�̖���;Ӆi�.��´��N��ET�*��
�`#~NOO)H�{�>��~0��k�7N<n�~僫�އ��]������j�k�y����������ݵ�VOӅO��l������7��+�폓ҵ�ٮ^]��:�&����9��e?���w����d��O>��^�����������`�*���-��8`�����c96�������R,�g����u���{�:���gc�B5�s����3366F���?�sg�Y�4�����-,,�(��g�VL�o|�����������D쾕����~�S��]۝��r���;��t|՞�U��o��X��_[_�p�n��W/��������3��[�t��4�~�kj�^P��5aiו��+�kj�I�3u��      �b���c��x]��&R���8o��_AC��@�"��{lb��Lx�R�2-P��p=����1;�i����_:�=�6R���!?~�����q��yO�{o�"�y�����q�Ń����W��t��z��atǏ�w>����x��&��p� �{k�1I��Pͬf�/�ܢ�ҳ�4iRѩ�������|�;_G�O�I�u6���D�Au��nIj#H�����N*����X���^����K�0;;�zE�2���f�Qfsm7�qmS�-�1���gB"�fu5�Q&k��Z���m��u"idBr��$�Y?r�:��M���&n����6�T�Vy3   I�%��N,<
��"x?������'"�z����ա���Odn~�@40�;�b�ȓdw�^�W���uDq�:X�P�{�ә�T<D      ��ԩ&����H�'����F$�y��ϟ>c*s2�kV�o����}va��C6�9���*�NK4>5Ic1��ۍ��˥��߽�:���ޣ�Ϟ���hd�g�LOOOS\�y|#n�����3'if ��� �sg��l悸���দ�bsp��g�t&r�g>z����׮���w�?������L�����D��X3�s�s����pp���n���E�9X�E�Π�_�؇mˆ�~��O1���_�s�rog@��y�R���X�$`e<e�"w�rIoQ���[T���LZ0�m_/^� 3�3�6��mN���B�Q�M �ߵݱ/�k���l(߆ \�u������k;9��Vh�����)��@�N�=    ��g�ra�vv����wmW�k���Q�����������{�U vvvZ����Ůu��+E�
GgN��)��Ur���(����A�     @�ayC�K��Wn�ٶ��^��8 ֶV� (&cāh`�-�L�   ?�z���3=3C �6,NZn�-%���mP;_�ꟛ��5C�u����R�� �tI��u��mT�#%��f	Te�vˉ���`]�n��Nr0�딅'''�)-@�L�~�;�o-@�v~?*�� Ж���rm7��6D�ڮ�ֱ�o��������'   ;t���t�>\ˣ��k{߂����Gh�Ph�@�4z��-,,�*0�mZI��c��y��S���.�Z�	�!&       �d�e���q��.T�۝yC�����2��г��B[�^   0����������^p�lf-6;�1�[�.�����w�+G����r�bސ�+����y�d�4�\�����2Ή�(�/ޮ(V!}nM�0e�۷o9m�02>1N��QS	޹Z�x�[_��ߵ��Cǵ]"ZW�Br�%&��m7?NѸ�������sg�ѵ�:?vv����,}��o   ;�����U�ݟ�]V?R�v����}
��
A�.��=ө�������AP�0�V�l]s����ɬmV�b���x����D��c=D
      �?j���^�\��'�|����v黤8o�^�j5��F��������W���   �a���'t��З��^�&�)���R����o�O�C�s���]b��=�\K�to��g��3?)M@����Y�Q�R%��N�=�2����R%!��7oބz`137�k;9�um�H�.�!:�v~ �p�����	�H�o_���{�	��k���&   ��Պ�u�]ەM0�v���1Ѱ��@} ��blJ&t��Z�{�ʸ�w��f��K�0�]�E�vO�'      �T�ʔ�f��Xƣ����;�ud3@�����O���D���/�@!7�r�   �6�Dq��p��Hl�&�?��ڢ���ĘW���/�$�vY���
�X��!�4~`>
��r����'���:x##���,H�)pqb\�T*n���IF����G ���;�'w���~]��u����~��{um'�ߢ�]-R�	�[?|����nP�P��]�   3o߼���q:>9	ŵ]I�޿�<�v���꺝�1��w�ޅ�_=���΍��ҊHkk�6|__��2��]Öٱ,�b�*      I���Z3�es9ǀU�Y��A�D|��ڷל��_� o�095E �h  @���^*)���n�XI�����m"w5�Fg�n�%�%�W�~�r�[f�Ŗ�1%@�Ѭyqے������X�2هA���`�;;;�����	�Crm��J���۵��J��N!��q^-�]�Y����+�H�]?��d��G����   i��Ç��?�1�H�µ�뱒��η`��`S�� U��S+�]�Rv����A�|�S��;1�g
�     �T�3ds]ScY�B�@�7�	�S�7k�5p295I`�-����   i�tF��Q*���9M��A$�9�s��r�gc;�L�k��8Ck��B����c���O�Ƴ�ո�3ɓ�ݝ:��qg��F|�(C�*:����t��Џk{�����n����$
�em̵�l�µ]*��m��������O	   HGGG��e�R��{��_]?݁ \�yFG���7o���f�T���:}s׬];���*��C���w"�;      Ief�y�^�;�1�I�N��3���ʺ8����Z�5o�T����F�����fq~��>yB   @Z`�{�_���%0�����=*T������Ͼ�9D��z���ܡ3o���"�͏e pj���j���]l*�6��V�2+JV��ۭ���{P�ޘ���
ăpm�]��P�յ��/��֕�v��i��������.��rm��'������4�R�D   @���+�+��{=�/�}߂u�u�ۏ�(��P����|\lmm�?IP��Jˮ�x��0Es��֮',/)�B�     @R�.4��+vc,�l�g���]���l�לagI0Ȋ#o���[�0��������O   @Z`��^��;�9#ܣ����`�-e��&M*�f~��yC�v6S,��,���j@��ɑ��̛��rY���27epJ���3X��=h p���q�Eꌨ\�u����T�n4�^f\ޢ�]���\����|��J�е��#�Q��  @�`.��|��ժc]�N�pm����{=���~���4����ׯ_������u�w����U"ws��H�&FL�z��`U;� �!��n�#Z��CU      I����IgA�.KP��^������ڍ1s��5q���;�~)���q8�?��    a��v��I�u&u���kn����|��*����iw����ĳč����mIl�A*պ������-�@>c��Ϗ�ir��rm�������2lr���vq_����gLW��]�p���n�K����N�յݠX��Y�F�  �.=|H}ﻴ�%@Csm��=���	˵]�:;7�{�����ŋcmG��y�S"?�]��q����(s}�iu��     �dR�4�ݱ�bsI�� ��;�<�ob�l��fz��$����o[�RA�0"F�E��!%f�߷V�   �6�:fr����y���?c��l6�z��U��Vi�5��7�����yC��\�n7��Z��4�^�O
Z���+tuq�'�5�zc���8��b���u���c���!>3�3���k��˵ݱ/_��6xi�b_��b{Tۅ��n�Y^\���}ZZZ"    M���4�}2ҟC�ڮ�
�l�nR\��z3�D�	D �L]�pa�T"Ҁ�!l������j����}68n]�%��      Hy�F�1���>��K�����.��+�����Ak�319I`�Y?�FO�?���Q   ���˗���J/67	/�0Ɗ �3<99�����u�,~w�[j���f~V�myCu��܂���V��� p�I��wS�ncOb��m�|e�m�R��~�{{�f����𙞙�<��~\�u�k;_��=7����Ե�YG(s��7��A4�}�]���Um�~�&�ƨT*   �6�=J�Vϵ]V�g]��{?W��lzz�@������n�:����$�+Y�S:�T�-��J��H      ��mԬ{x�'��O��i��yC��;�K_�[7J��!����	����<}s��   Rǋ/�~���9�S�G�u2����q��m�*rW���{���e��|�8���[�ȥG���3�L���w�ywpo?'�l2+I�4԰/��G��sb��q����� �m�k;2��3O��d���N⾽����	ǳ�K�-��V�'z�Q    LjoS��k{?�p�v]�g�aӏ[^�T"FL��C��enD���w+>``�͛�h��2      ��Vo���!���6��u�o���sW�O�,7��C0�:�����a&�e�y  �J��*�s�L;��(���w���ի�0������7�q�g+o(����F9�`q��|���L�9�yubhc�L5�B�j�7G��i_���m���#���a7��2�v���pm���\�M�w���2�z˵]�_IYK�b���"rm7D�e�j�   ��rvV�\6G����P�S��^(��Q���'n����31g������TB��:i�]��k�d�pbw.PU)�       �Ԫe�}�Ù]��n�l��=j�~�chk��i���7��h��'0�@�   ��gp���lTt��m~6-�µݹ�\+l���3?ט�==3?C��Z��z4�N.�v�4��Yg�����~?�I���@Ut�@�Z�.X�tm'��Q�v[|��K��:���n	Qt�v$�G�MR�z�v/m�(��R��   ��勗t��y�~�α��A�۽���\u�;>�{d�)�t�;@V�Kf��:�*Peݫk�x���ئSΦw/htRF�     ��Q��)#1�j?�r�\��&n�d��F��a�0Ɗ�����%�ɴ�   @Z��|f3^p?���_�����>le�6U�L�7Eiw��@s~�"n�<��Vr�O�*����񉎮H�S"�ٵ]D�"tm'��D$�۵]�˶�ͭ�"/��q{�6q��F���9���$    ��|������]A��k{�'��f��RE]YMi�Iq�H�\��5�Z6������V�n��[E�蕲/	TA*2��f]{�J6c{�0���2�m      �D.CT���PuTU��I�X�^��=g����-b�^���7�cp�f�����6   ie�y_9;3C�
C0����=2���"������� ��Frl���s��kYB�x4���"$R����ו�-�@UX�#P�v�@|8\۹�+�X�
޵��Nׄ2_��n�v��r�=�n�o~�   i�\.S&c����ڮn� ���+��ӵ]R455�
J�p�KM��6ʴ�RפS:gg��a�1�%,�p�1@��S`��#      H��l�Q�p6����mV*\ڇ���=Y&a����	��^�� ^έ��7���   ���js��]\��}����=*T���ͯ�B�*T�5g��ߙ�k�:��htRI�������Ӆ�=���`�9�ɦp��T%�m����86F�\�+q
����D�2�k;WOx���zw[���+�N�筝���nַ]���n�x�~\��c����k    R��ݏ�յ�_q� ���u�g�!p� 6�*��
~{~�h�D��b2��!l�����=p�\�x      ���"�p��y�}�tJq3�o����	Ⱥ6��v��ä�_�c�h-�R&�!0�������   ����+���'��|>O��<U+U႙���g~��ڟ�f~feS��T� p��T�y�4�y�t�:�)��T���QQ<r4�����!>����gN�z(��2q{d��rq�%V���+qmo�R&@?�����;�C}���u��   i���=���õ=q{���:Wsbj�@�looS�R���QFTZv�=q�8���8����o��o�:      ��D�y�^�f^����,��|���O�$��V*r����������#�    ݴĭ�v_[�����A��R�&{��Y��r����#�����c��Q�'��`�#A�]��
D��TVY��d���'�h�� �������=��KD�Ra;_dkC8���l������zsm'�����)\�%mj��1j   p�9{��tZ*�^�k��v�k;�����9::���cO��u`P�]�ޮ�8�,�z�`�,�0�m       Y������Q�ԃZ;6m�}�#�y��8��35}����̸`�H(�C�>�@�   �$
��0ּ�=܇�=l���R7��-��ʌ����KA���^�5�@�x��J@��u�A[�N��O��:ʰ���#�۷o	����d��h�qg������/�v�p}�]���"���   �v^�xA}�ݖ��_��JDޏ��o�vV��0���`�� |�����#� W������*:U�p���`�Hw      ��h��4�o����f�0�U��6� ��Y�)c��W������16>N`xay�ӓS   �N�Z�|.G�Z��pR�}m0}g�f~v�˶w��1 �-�`�5h��iw�欋̼H�ܕm��t�J������+ ��	É!��ο�z���+µ���ί'nwݦ�v���PG��nqqv���{�   ���:�86ޟ�9\��u��tmW�B)�o.�p�
э��pW�N�n��+��m�K�U�s.֐3�J      ��P�ڍ�x��^����/h�P'���+��!�� >�&��˹�U�z��   ���zk������M��f&�6����i*g~�*t��r]�|68Q�\�@�$ZS�{wpo��4��*[R��s��~��wmפ�r��y!���Nr'ٵݾ�ו����Nܱ'���ݻw   ��F��ZlD*"���o���������"������!P)]ܻٻ�����\p�Mܮpp�Q��      Y�5���;?PULL�5;�~K�P� ZM�7�q�����7b?�;�1�W���E��G   ����-��{߅�}�-��xa�m���Ѱ�w�g�Z�Ϯ�tup��XȦ�o��F2�K���GY��ic3�kk�H^�0������TED�8&��ڮqE6�v�흝��u܅��xum��-��k;�_�T�U    Q�w��k{���u#vm(���!*،[i��� n競�VĪ�`=��� f��@�     @��i������J�sי���FS$�%�H�	�888 5�l�!    M����(�{���(�Q��kI��9��I�X��ֿ���0�$17���=�?� ;�߁*S|��bN�U����T*�6b�6tC"v�����yumׅ��(�䡻��N'���tmw�����n߮3�E�7G��
b{r�Q*��|�4�u   @�z���\!y��KǊԉ�O�x\��6a
��`��^�=��+q���BA�.	�����      $��^wܿ��V���0�}�[ZPQ)�.R̯��
�Q(��	   ����h*��=:�`��:�b�(rW�����G��{�X�0Ki wd�nsTk?���@����TE�hK�����.��kB-R�	�ܵ����ڮ�_���   ��ĝ(�vy��tm��"*�v~E6����U��2ȁ*�y#&e���U��*���+b	�:n����      H�������A�>�~)5�B�0:�1b0�:    R�����8n��̳|�����f��-o��4��l}&E�s p�T1����c�M�#
�)`�v��]������]�S/��O�MH�y�;���(t�H���7I��]�5�u�9�   ��κؼ�)��;��ȣsm�'��n���"��T)����ciybL�j�s��vmK���&�Y�������      HZ�2���߭�b�Ј�;M�4IA܏t���ӏy�I
� ��F��>�@�   X�wq�����HKͦg�,nw��+o(�se|��=6X�0��t�ePp�ii	T����{40��\>'�����*n�^�Jq���.n���������}��!�wm7���l�Qr   @�x��]�z�N�$��pm�Y7^�vU���c���{�Q	K`/ƨ�AT���
w��=�`�����
�      $�F�b&�����;$�:�DY�Q�c��ݹ�7���h!��A�
*��	    m�ad&��FƑ�H.�k-�f��~�kq�g���l٬���5����{,�����sMC���^��"e���&�m��|>�������l6� ��b��>|Dַ� �v<S`)Ĺ}��v�wg�=xh+SȦ��o��f/h�tpЪw����M%��\��vک���C��3�m�tyc\\�e������Sz��M��9m�z������*�J��1�<�j�J�r9��f&@���q��� ��z�y�q���e��q�;���8�o��z+I����١��#�q����U��w��t��ݞ�W�%O0a���;�>õ�g��tg���q�k���ޛ�I��g�/�̳���>���[rK�|���w����iw�[�ǲ{,�#�j��ե�+���Ȍ�8�	F�@�#H�A>_);3 @F1"��}����,�fξ̺�C6���?��;��q�˹Ee��p8����7���_���!d<�"      @��N;?��Hu��zᬼ�3���W%Ņ��6�.�9����}�\֙۷>�Ã   ���#���G�׿A=a.�,�	�E��s�M��r��`]U;4���y�:oȷ�O�� p��lqc��tO������lR��	2�M0��+Q뛉M\��oa�7n�ѣ?�@)$+�=I���I)��W,l��Z<���ӧ	Gt��\�SOc���x�v?(�{�����,�'T�	�}���z����Ŷu���O?�E_�{������Y td0���۷�L�y��M��zN�g�~��'}����z���յ��	}ٽ�w=)ux��wg�|ϳq[D�~\��ڙ�����}��[6�p�������w~�w���p%�����OON��gOu���]W��>�}r|LO�>�4VwxW�����^��w���������>|�������M\�-�(�Y���s�A>eL�=E�p��x���q����!�j�!      �g:+���aX/��In9g��t6�ڥ�,�-6���ަ�p��`0c ��������ܟ������~rx��5����N΂ݮ]prtl���8:��� ����췫��-=��\��7c���#1e�_�И����kg�yv�̐�,���}W�L._{��3�&W��������>o߿O������q������a�����X�~������k���%ɇˇ�﫸+R�s���z�͎���%�������������9�2A����$vpWݘ��hɁ*�q2i7?�_�@[�Sf0���*X���us�?�����7�)Ru�//)���_L�B<�/�:m���H�õ����:e{f/��P�u/��긄�]!$_���r��m�;�Qt�{A�׈kG�K�/=�����ݻ���AD8Ha"'���� �\����U�L��^{W������\�&\����fT�=����>o\�ۇ}�
к|����H���q������g[�� ������L������h{G���3f7��y��������8H4����:�n�z��Hro]����.�i�y^�v�p�Fܾj�e���i����;�]���6]M���      @�_σ�\<L2�b~���9!d7�&ʪ��(&L*[�Jx��]��p�.=���V�~��7��ӏ�o_��ݛ{Q\�6Lxe����?�3����qGe�����ٳg�
�����̙��������Ύ��8]^;X�{��=z���/_�7,����}���ݻw��������l�����~�?����|���W��{�����1��o����}k}3����F�"e�y��d��]ܣ2}���q�_�/�^�+����)@���ٌ%��7�|S����nX��+8A�l�%q�Gf��B=^����~�X/\��~j�X�n���ɣ����~��Jr�K�Ƶ��P�N*�����}e������"   �'ؙiIyZm���
���3�V�r�pm��s���I�@g�E5�
���E�"w�=�y^��k.D/��      P������O�$s��NɹAZ:\�$t7�ra����\����Ϯ�a   �,��>�?�yC;,3_�onQDm�ū�9=�p��7 �'cw��m��h&,yߞ�db�Y�̎��*��-*U�����ȹ@*/ZH��tmO
Г�<��~FQ���Ke)���9������]��O�S^����F�ΘM�   d����x����YaѮ�i��ڞU�l�v�n�7Uv`w��
�]SN�L�?�i�A�n0���ۅ����vgM      4��`�<?1v�I��_��>g('���椬ݙ�yC;�;!�����}   �t��Xk:=7��7�u����[��u�U��0�=e�7d����kN52�k �!��)u;�L7~�E,�M:1��?
vbX�@���9��	@���.�M�;b�Q�k� $�����.���J��Q����e��     �o���U]۵*v��+������ʇ�ט����&Փd`�K�'��xu�8fO�x^<A��;pp     �:lt��x^��3�5�k/>�����DE��?ߟL&��:]�    �0�PS��Ev`�X�`|]�՗Co��7Ê��۹8���6o�S��Ѱ�@�G�[$�c��7eRԮz.�L	N� �b[�_\\(�n�oϵ�Br&�D
A�\پ�k��<Ȟk{$�����?�6�   @����;� 9*�v�k�%X/ŵ]����H�ڀ�3����e֭���g����v��EU�굪�       �K�෗H2�P�?V/xU�N������bwg,�srrB�|  �9�   I<���L�V`�ټ���Dus�zq�X��;�tbɰ'��{�+z��m�pR] �lrND��v"��H\�V��H�^d��	�///	�O�� ��I��um���]���Ūk���^)R/��]#�O�rm��-|�gT   2�g��ߠ�I�cP1���������um��E�[P&��`8�:�L+ͬ=�<17��uΎ^\!��P���=      Ua�s=J�qIgE�O���H=P��0w��H��vC�� �w    	�kM���6`F���6fչE3q{��n�z��>�ƹ�TS,.o����,W p7d�+�����I�%��X
TUiBw{���e���D�Zq�,l�D�NH.���ޑ���vŻE8G���z=�um��^��t�   ����)���s�;\��ߵ����5F�Q���mbr���R�*���)�G���     @e�D�U�<�y݋�s������3�VӘ ���!(��k���/�ì    ���z��n�1ެ)�>Ʒ6`:O��s}�'n�ŪDQ/�����yCw �n��n��	Qn-�V)+,<$�e��n�^#sGB��/O+�V��5BvI�>���ubm{�풐��wm[ԞS���b�D	q���f�O���     28?�~�W�k�����!nw�ڮ�[����E"�E8�7C ���"����>/�;��,J     �����bWpE̞C��x����ԨJ3([�Y벃X@\��lmmqQ    �紵�Ig���%�ځi=�1���nf�Us�U�-�z��Q��;G�!��\��7�8Yn���W���� �i;t��V�� ;͵�����'���'�*A|)��A=Q��[v$�]ң�u���5��	�u��^'�7tm�w/
�766���   @�- S�Q��ڮm���i3�C>�����m�)3�e��ֽ칽b�<��'��ږv��x��      @�t[�|	{ ��Lɼ�j��dy6i՗�Uiw�4 p��*�eg{�X   �������{M���ln����2�E]�д��a��X<F�7\����^��i.p/̉�<�T�[�V�+����\����RYȭwmOuW'o!���u��1���K��<��|��E�9Iu���K*���    l��^��/���Zy\�]����"Z�����x<��#��x I���"��%��bt!p     �2������S������ �����t!�+ۛ��pL    �h{o�@=�$r ,��䪸��$�T���H��z�"q����3���k/V?�&N)��e���U�`_� ��E�E���Y$��k;�k.�v�pޞk�X�ͯ��������+L  ��ٌ�er2���4'q��pm״��k͒���O��{�X!Y��E�	���q��      *���RZΐ�G���&S�u�]��d��%ǹ�;���Lc,    	�~���>�z��4D\��yk]s�&g�(D���ý�v3�Ș�����
O�
Ik� ��{���:mYQ�L%�����.<��vw��i��������ڞ&��w�T   �@�n�ڮy��9�!n׾�>u:]�e�%p_�����\��
��EnR��b�ߦ      �A��Gۂ�����k�������zTU��=�1lW<PO666
   u��j���ԓv�X[TA��2�-c��?�_����o?tz�T8�Z$x�խ��ڎ\s���!L���	�x�v����r������4��I�{��|)�v�r��/?�������e�vA_   @���]du�v��]ە��uqm����VSq;N]l�m���5�b)4��H3 �a4c�����g[��6�      T��������T�+}�b*nϢ
�U�B��
,�T��`%��e>   ��a�u;]��wk�aޖ�[̓3̚Wy�~�/���e܁��݆�����|ERz�w�V��/O,�0>�E�����]�)w�um���ʶ]۽�v�sZ��]�P�k{t��%�)   >'po�k���������"�^�@�4z�f�J���C$�)�W?�      @shyB�c����K����z�1�
�%+�p���:po�7�%    @u��dmas�V��4?ły[Z.��M�5=e� y���t�f�������)�X��� [ʧ91Į��{i�v�q�F�v�@�N����v�S7wm׋�m�e
���/����u���ή0�v�3   @�l6�^ݵݼ��uӺ�]ۍ�I�f���<�]�@� P���y~R���!�     @eh]�ϧ�'t;?{&s�7�C�    4��:�ƹ3�J'k�V��˕G09Ts��ɝ�cu�TCZ|rY�h���Q�د��.Uv�;[.��j��\���R#���+�����q��k��J��TG8�?!\OI�b/��׵=!�   ��l%q;\�+�ڮ?�N[I�`�y�Z���A8?@�0�+��Қ      �CN<��{��9A��Oe�#�����    @��\�sǘR�N��u�-Ff׺���_�V�924�?�Ғo�7KB�jt�z���\;���c��ڵ]U��k{F�+��/Z�����t�,���ڮoW>&�k{���3    �!}O�ھ����v3q{���Δ��qm���nl�hNr�Aq���K�{�'     P!�8��:�񥌄�v�d}�����`�e�N�Z�#�    h��d�ic�k��tJu'�+� ��(M�/ĩF�D���]x�d��E�J�g,� )`�f+M�!+P��z�^t����5b�Rn��*��+�W���/�s"�\�iQ0_�k;�<a�   ���k�ڮ��޵}!!��Rq�cVp���� ģr��k��{y�      �J8���a����~�7���>w    -�'�ƹv���ݕ�ܧ���7��e ��	X���w����j�Jsm�R\�%��R��j���T�k;Ie�Ӣ�w����    J��ܕ��S�6=CL��󺪚帶�z�E���u=�E�|0o�F��NiE�Ųi�      nH찔7�'��6�n��ua��3    @�x��`�g;4:ohl�%�I�F�����.6�s�^C��D[GJ<����5H�H�A(a���=�H]S��?���I�r������uumW֡�\���|�#   @�j���k{ �^cq{^�vS������|����y�V�K��-6ҭ��U�     P�Ni��ZVN�@f���ÝYoW      �y[:iW�Д���⑿|��3.�nv xv`�Y���]��e��(��M]ۓ���,�v/���sm׉�^x�b_�k{R�ηS�k{�>bT   @*�Ʉ:�6M[�5Ƶ]�ĺ���k�O�>��Eշ�>��f'�dm�     �
��3P3V1�B����f     P?`�e�ۊE4�V����Z��!ѭ�%�j���s��}��m��l^�k;�(-�۹���%%w(l�_µ�����>�ye;庶׎�   �e6��_%��!�^]����B��d�qx�\�yZm�l�T��^-�[�r��     P��s���OJ'���m��Z<X`m�C<     �c�a�{�r��"h�!p<e"�zcV]@�@���\�M��Q�%�v�NX�.��-3���   �c:����pm�q^���pmO�� �0o��JK�1�     �2���sO)c���1p      ,&_Vh�-���I�����E�B+͸�!p7f�L2�U��C�k�v�-:��ھ����	�b�L�v�ڎoE�B����*��2���c?�b���+�����Q[r!    x�[p���k�Yai���4oXQw5�v�Nvhb���;˰!���      T�<��RWc6�����    @�h�0#��m��l/�O�F��8�t>�X�t�h��]�c��\�.�U�k{|J
���?}��k]�=�A!��T�k{,n'",   ��0���祮盾�e���`Km+ PU,�;`|     @u�R�˴c���6S�.ͩ0��vī9�+    z�=Yk<���y�Er�Ư/���]��g�V�]�k�T��ڞ��k{xNĻ�S�Kqm�����pm�1�   ��f>��#Sq{u]��륹��XP�k;_	Y;`a2      ��x� �M0���)��2    |O�*���F�O����!p7��Ce���̵Ԛk�,Ҷ���I='*��]�vV�+޵=)�O;'    Ȱ	���1Wwm/���L�^�v����R����VN6@�*/�     P��(�>Vh�ٲ��Z-�M�   �`�Yg�X����H���Mi��P��b���^�k{R�mѵ]�/�'i���Zյ]QV�k;��   ����攛d�µ}q{����r\�źH�١�n�      ��G$�&JX�uma�3    ��xX�l���Ҕ�� p7��Cu����ϾX��V�n��NI�5'$W���"ɑ<�k{xNJ�}R .��+�'յ],Ksm_�it�j���<n	�v��    5��۟LVvm�S��庶���w      @S�@?(�?� �����F��G   ��k��v���.M��A�n��1��}�@�n���ݡE��=N���k{�%=͵=)�����	ι:B_�t�'�NQ��r����.~�,��>_}�8   ��m�<�%��k�ھB�"\�5��>�"��g>U6���X2ߓ�     P0>�
柖@
��9a��    =��,��m���M wc��!$�*>/��v����[z�>X������y��>�L�g?���I-����5(R�ˇzRm���{�O��O?=�w��,J�K.8?;~�y�J(O��g��� ]כWo���cv[�z�L��.���c�bg��?.<}rr�(��`0���sg���驳k�����Ņ��ٵO�Sg�.����ap��\���]���w�}�~\�����}�M&'����{�._{�Y7��>oٿ�p|Eak�<��d���7�����r͕��s���o���n��n����k�����zZ�Z����ѿ��E��NNi{{�l������}^U��2)lJoؐX��*      ��vI�ņ�V`�&W���*;���wO_[���f`�ߘ��8�w'z���b�;��*�\����.�	�]���!� ���3����.m�m��!e}�5u�b��B�\L���.`_&����t�x�[;������k�S���#��k��~���;�ߨ��r����K\��/����E�U�um��?|N�'̟�b逮��}����}��	����+Ta��gϞ�޼yC�nݢ~���o���ٵ3�%�޻w�I�/^���O��+\�w����{��{.py����mmmY��v����۷���'��~���ܹ�lq��מ��������������Q��U�k;����~F��\�Y���wS����~�&�	=x�P8'�V����?��E��g����Ee����`n|��A�     ��0�rɘK�Źʎ3�\��n���C��l<�_��j���prt��%np>�������k��}����q` 2?.`F),�
f���5wi���w�?�ײ�+C6�A,�r�WWWN�g�;뻉�L���\��l��L��=wtt�Y��+�~��B�gc��_~M�p�����NzG�q6��ݟά��=�Ɩ^M�=�p����$�?9�Cl�fC򆸫�ܝ�d::M�R�Tܦ�+<�o@��7���䲰]/$_Ԏ=�>��ۓ�m�2~�\�u(QG8'��Rl??���^)$׉֥2_ѷ����e\;-\�)�^���	ۅ��#   @K��"6+L�nV�L����fuu��!n״iz^�^�vq���-(�C�ơ��K��f��      Tѥ'��;C��ĥ1V(4q%:�}��}��O�����o���޾|\��+��/�������S��_�u����������&v�裏��s�U�̜�����������w����>���M.pm�Ča=z���/_�7�.۸|��w,[\p��]'�7ِ-���_������������3c�*����[�f��;��X����湵�>˝mll�8v5?��9�HB�n�J+|�B����S�����^3um7�k\�=R	瓎��]�9��\'l���B�%��'������r���:    H��ti<��]]���*X7����Nʺ�\�՗5/�A%`WɈ��X��0P��0�     �:,3>��0]]
�m�     ��Hl�U�mkm�U���6���5�	��7�p3�Q��(�P)����lʜ-�tmWG��k�(�(ߵ]<�pݒk�J�_�k{�1    ��Zfߓ�\����uum'��*˵�o����n�u���?V��xF�#� ��=      �A;3Α�NoI����V�-b��f���Y     ����Z�{�'�b���!z�����ԃ<;�/pY���k�(ZW���K��S�Ϊ���1wm�w�+���'������4�   � �{����f�;��\ۥ�q0ٲ�m�ķ�/�J������       G�q\C���������   �L���09�D
0�>�#T���		��e�q~Z-����7R�l�0�*;��W���wm���C�rٍ0�I~i�vE^Y��+]�5.��)��
��
���9)�Ay    (��E�smW>������0\Wעk���ނk;_w2(��*gcނ���Z���      �Qχ����G�ik[A��0�aG�Z��!    ��q�=o3��/gl������k�,g��Sz|K'�?Y�B�k��xBŹ�3�O��.	�=OZ@dٵ]hWю�k��^�k;	�H|���Ν7�G   �������3���ZŻ�ӏ����ڮ(]O�q.(���������ߓ�Bz��     ����}2�:$���`�,�;�0�N	Ԙ&�   �e�x��L1εB��������7v����=��C�n�LvL�U�N���:eͳ���@��%P>㫫x�fŵ}Ѩ�	[��Ȯ�|��]�e�k{� >Y�_.��k{Z���Z�y    Ĵ��I��++j���}�z��tuM��Tw2�������z��{�틇p�^��Gm�k��     P3���9���s��C�R��"����?5a    4���\T]�^Dnr�i�<���9uÜa�c������!�@���UR&7xx��Y�ދ� p�T�>۟�e&$_ŵ=<�+[Ƶ�?Gc�v��X�k�HP��vR|�*�a�V�   Z<o�=��k��0���"\�M��Uwm���ʧ��0'{�/�3$����     �����)Ɣc)51X��!yC;La      j�t�q�ʞ�U�<+3�g�?�:������	���{���ү��Upi�P��Ɍ:�Va����K~�z��3]�I�Zn���yU_tK����*�rmO�7���۵�{�Ն�   ��j��yWum��4���k�I��u�]۵���w+4z�f���ew�<�YE}�<      T6>���YJ,�������ք�s�=��0��e��W    ��k�������%�̮3��ɔbv~q�"���!��;bSQ��Lb�&���mHuh=)"����	�a2�P�;�((׵=n[)nW�ծ�|l�ڞ!Z��ڞ���������2S����Uuf3?<\]]    DB�,�ھ>��|]l�m������`� ��ח��!�     @e�r��,S,��s����S�r�=%� gK     PG�7�Cּ������+�Қ�)v���x=	wc���@�N,��Z'���[�*r_�a���A������.ѵ]�6/���ڞ}>*��T���]ۃ�|^�"]ۥ@��j|E����   
�&�pm/I�_�k��x����T>Х�p��ȡ*��|��=!�0gF       �L���m� �fMZ�	�?&��f���Q�V�`�-   �D�Ŗ��l6~@��a޶jn2���Y9q�� g(�9n�m��!WS?vXX������aC�[���L&I!����	q���8��F���ڮ�K���Ο�ޑ��v��j<���:::"    ĴZ���Utmן�y�����L��A�|�U���H�[^�M�     `���@�sR��!���3����s��L�v�?Y�3��LgSj��p0   $677�rxI��`�c�*����M���l.��F>s�gn�;�5#��!���P�xnm���U
9�
�1�{n� ��ڞ&n�]ۥ::���̢Cu������w�X�F���FW#���%    ��NF��'pm_7�v�Jv��E��=D��{{҉!vl�)�=��=0�     ����z��H��}��C�_U��a�i��dB-�޵d0q���S   @�~\\�'l|�P��q3̳�x@"�(�T��L��UC���2��D�>����fl�q@h!6*�2�A0��t:4��b�LBqWp;%]�����e�UD6]��c�'�'�q�Lҵ]��ʮ���O��pD�;;    ����`!O1��\�>�$�v�C����9i��k{�Z]��ءW'���M��u�D)�Nʭ����X�     @e�L�s	>o�\�k�+ա�dU�<;�����d2����>(����   ����w+�y[hh�DLf�������������b��UC<� p7d8���Z܍��N��B���(����`aۣ�-` p/���0����>W���ι��r�G���um�(ص]����S�^�k��T�p�΍[    �����Ǧ�v���~�e�����0��E�:��߯+:1,2:      �>��z��������e�;�u��JN�����mnm�L��c,    ���6�9> PO`�e�:/LNK杧���9�d�����\2���~E�jՄ:q�6��&ĕ��P(S���-C���9kby����
pm'��[tm����v��{��=lgI��4q�*��]sN�y�um����]��C���y   @f�����^�k��/ee�s�4P�k���e\�yF�!;��!�N�N��      ������g��紂v�LSt�j�xeU)7�F8�\�s]w��ԓ����=�1    ���_� PO0������e��������]�Hx�=5j��P>r9aw����/�7��h�Mi(n�E�������0��KKvm����vmO��tm�}�:��=�k�\��j    Dvv����}�3��l�p�jӵ]Ӭ��}Eq���[�k����n5�,�*ωA�$��|��C��       4���F�.!�_�|��w�� U#Sh�|9C{\A T[���&    ��\�@�;?ۡ��Q��5����Y�A��H?��c�*�3F�������o���r����3(Q���R��5��bw�B��8 ����]�CL]�}Eٲ��$ճ����.ӵ]��Z    �^�O�	��Y76W���z�v�����
AH;��Ǚ�s�*9)��*N������Љ�!�*      ցaV�M�ļab���d7��	�,Fа"�3����3C TW��)u��3   �;��!찵��=���F�{�a�#w�q�V�{~4�F�LڝvꪈD����SyTx`j�����%P>���$�.ϵ=��%n���D*q��k�ԗ-����)�^q����!p   ���G�q���y����z�����k��ڮ�:�����N��P_r܃�za|�k�<�-vI���       � 3��[�D��.q�{���I��-wu0q;�(�1@     �F`|k6_�Rް�-e�_ۆ<�V���/��s��|!W�r<�& �{:�*����J,����Q�*��H\(A0��0�.�j�k����ȵ=^���c   �i�ظ�\��x��u���k��
w+���o5h�����Wn����S?*W�������܉aM      4�`���	��屾8�O�V�#|͜dM�ۋ�-���7 p���     4Ƒ��v`:O�d�N�;�d��wf��^�Njr�g�.���B��&���f	7��	q�3)\�(S⪘U�����!�ˮ�ĉ����\�#B�ԎPV�k�ܽ���r]���a�"]��Sl�[�0l�A    �i����"\�M��并��˴�uvm��k4���l��o5��@ռHw�'�+r3Z��Pџh       �`0���X�+�3٢{�A��oo���E��L��g2�1^�?/   �� �^o��nf����C�q�"g��B�Pz.nO�*3<�E1p��=�N����Ѝ!���Rߐ2�_���,k����m�s9^�
J�ȵ=ֶ�����]ۓm9pm���}U�v����3��͛p5   8d'���V74�6i�,�v�x4(�f-HNT��W�$�
2�+R��=4%R     �p5Y��Iqf���u�_�,n�jn0�]cY�5w   @�Ÿ��[;���X�ӭ���A�\_�����34�<b�Ӧ� �{ڭ�i���v⢛;&]���Q��]q�u�w�T���|?(ӵ]�N+��gԉ������=�'h��ӵ=,c�?�t���  �l��x�(µ]�@��4�vCq{IךO�nVw�v�����q᜷N��8F �����zb[r��m��4      ����t���ũ��w$lOI\7E\���yC;\�  �3�ш��~`�   ������@}����{5�j���>��BS��V�9���\ix���I�, �Lp����`X�f�����<��tmg(��M]�5�\�e}��	������U��Y�{�9ђ��a���~B�߻���/�K    �N��Ksm_Aܾ�k{�y���QWI�uu"�������gaA�U:Rcܯ�@��~��'      @���:4�ƻ0��ƄI~V�Z�<R��6�Z��`���C�Uj���}�����k    ��۷����@}]b�g�uA�.�)O�Mf�fX\/	�U9C.���w�)@��ߋ_.�M-�S\�n#�5!4ugpd��r�B��0�h:�R�n]a���9��u�B�k��8U�n�ھ8s�����g;��ג��.����8{<��hk�E   ��������i���sˮ��Z��s;�//n_յ������6��|�,�wU�*��'P��A*V3      �j�j�h:��%T#�D�����)V2��k|�����w+� ՙãCzt�.�   ���wn�/���@}�0����Ύ�����v̷�Kܕs{NG̻���1��a=��Vw��o��r�9*#�&����z���cQ��H�n���-v����,ѵ}�w��]�))_ڵ]rcOз�ڮ>��\ۅ㮋�|�   !7�nқ���B\�U�õݬ#�-�������ŀ@�T5Pe�2U±r���q�U      �-{q�u���0�����'����3dl��
W���r|rB����	    s�wvhpqA���9���@�4i��oڬ[�.�����4"�pݮp�s\��vs��͹�����V�-�M���X䮉L���C�������7Vwm�K�����v]��~Q ^�k���#�jv���L��G,�;�a   ��v�[8Z�v��sm_�����D�1��A��^����!P     @=�Z�x�N�|A7֟��#�	�'U"w]�`�4a�s�ilC�n��xL���I5e6�Q+��    ˏl�:���l��g��k�"ͷ��w?�a�-��-�'c~�9��\i����U���`��������Uڭ�d��`ss����\ t�vQ5N��m_����c�d�vm��z:Az�k�t���I~-�qm�w�   "�H�,��<a0cq{��<�V��4�����&�׉�//.	ء��*mP*�,�D�*u�
�*      ֈp���?�"Uݶ�QZ�����3�r�MI'���ሶw0�-M��      ��C��MY�,�[���LO9V#��UZ�לE����`<kQ�spo.U�j.ZO&��U��ʘ\�UYg����7o��0�2�n�L�vr����EQ�����}M\ۅ��?��n�   4���F�!���k��n�v]��6��_bIk42P�,�>����f�"wYC�	T     �.L�v<~'q�*I'��|nn �S�+A��U<�c,{0!��N3��    h8X�UkF�!;d�������yp<���#H���yY�<���7��=��6��U喃~�+�g�B7fC�}�6�Z���o�����u����}���'n��C�޵]|�tm��WWWt~z�i�'RI��\�Gz$��������Xj�\�������$k��/��d�J�~B}��P������)������jъ�kg�<�q��_^^�;`K��k��9W�O&g}3\�������嵳��3�a��5p���~4����s���ί�#��Za8��6��m'�6���Lo��?8;7vw��_D��˜���Ճ��̺M�<�y�d����ɉ���s�4�<�7n�>�� P�+�T�s������b�8f�;      �c�/v~&1�����7z^h%eq�^�����v��Ԙ�X    �0�LW��h�q�-�0_K���8�ǟ1��v�����%��3���=��G[�`=��O:�II��F\��0��L�/���C�j���_����*�^�\�^&4qտ����1���h�P<(Ҹ�����΄O�oފ7/'�W6�����UH)<9>&6���U��PInvN���oG.;=9���_��ӞuX�P�s'��B�������@�w*,.�����Q`��3�/�����J�����&^����=τήv�py��]���N'�q���[�}��oo����:8:�%�6Ջ_\��{�<|E�vS�{����mj�Z�P(e�zv�{-s�|u��	�ٜ������\��]�-�(�nݺ������t��.o��
�K�7k���     �c�Ue����Ry(1�,˺�ӎ���Juqg;�r���Z</_��j��{W�����7��㓹iE��\pq>�~��9������yS+�p.����>���\���f�k�r��_{����A`�����}�̙�!���Y�.M ]�w,o���������[&���O���_��]��{���kt9��S�c���C�c|vϹ�[�Q�yݹs����*�x��������y�0��MG��ae��Ϩ	@����أ��c���7�ue90�n�Ď����	1����ࠔ����	�\�g���U��O���{�&]�tm�cA�O?��X �s>7rm��3��Vp�Oo^��W�?|R�k��v�Ne�����(�De����O��a;Ͻ[w��l�p��=r�l6�P�M�l�������%��g�����+\�w�lQ�����{.py��g�Cl������l]^;���W�����MP]��g�$���G�Gt:���[7�-���svzJ}�qf]��\'"7;/V���?���Q]�����O��{���R��kN�v�{��)���d��rn�FY�
�h���gM�#:%UIq������0�G�@�/-x      8g<��E_�E��X���(U&�u(�ں�6ff�Pw+K�biL|�0���,D�vߟэ�{V�f���'g���a׽��C�H���֯����g?��~��/��]�.}e�⸮�f0����Y\jww�I߮_{����<�[�����w�q�?��{ޕ9����]3��7���u�i���}��:|W�w��ɩ�1��8#��7��햛�����K�c|��c����Ee�yX��h���D�8@Z��i�C���)�@��8��*e��H�jP)p��P��J%��UpP(��P4���_(�r�i�	ѶFHN�]�ħ	ă�^��=����[ �Nr9a����m露���{�>�ՑNU��|���5������Lq��^����  �n  ��IDAT �mn޼E��pX7��\�j�dX��t�G����<��4&�W;������	�A��`��V�U�/��x=�����_h@�� ���     `]�<�h�������:f;?'g���K�ܽ5�-�y($2�T0������U��3���b�n�k�?�^�G�����;]��>^����G�����v߻�����g�T쳯�������"3csտ�����L����5ؕ����.���{�>Y���>��^�S�wq��v6�`�g�t��X}�c��]�����|���>���<�p��}�a�0-�m:�Ͱ�T��D�0�1��.&5^�.�{�G3�;��q$�WM�6B=u�*!tc�(���^7�2�۷o(�p��u���(�k�P�8a{�@<�k{�?��{��G|���BJ^sY����(�8r�   �D�-n��KD^��� �vMFuWum��u'�??s��aӸ{�n��+��� U2P%
�S�}��Ѥ@      ��ńh;�r�TC�y��� n1��G�r��:��l��3��K�bpA��0��v2    ǃ��v� �s��Ma��2̧�b����
G�P�.�+���1�`ܜ�.�\rp<��A�9^Ȯup���bPkފ6q���=/�!�ځa���dsy��>�L������Z ��W�k��������\ї��]U��r�*   �-����d}�.\%�_M��Sߖ�ڞ�g*n��K��v`�4~���n��'�L��a�j�w�^�xI����@      ��E����M�d�g�^\!s��� �AV�w~f�X�|��r�    ���M�\`\k��H�J��Bm��X~.�#�����1�,�o
��`<����7C�=@|c�7b�����*�;Q�T<{{{�0\��M��.˵}�c��5��'�6qmW
�C!yѮ����Bv�q)�v�8Sa��n�Iާ��A��Ǐ�/�    ��0���l�x�v�)��ȍ�jO�������*ܺu��A"��^��R�┸������`�|�A      T���O���z�O䅯IS,mB\)lg��Bg��"��� ���3#e�   ��t�]��	�6�]	��2�4�"��P��I�C��}~���G��4���z��ጚ�9���4�L�`C�;�}.0��v@ws�V� p����|!p/ɵ������\�E�wm'ѵ���s��g�۽��?E�^�k;W���>��C   �
[�up|�|�a��Y�0��v��e����^�	�S��H�����a0W峎�����(;H�����0��ے��"~�?�      �Z�\^����1}�N讛7H	l�����v���e2��x<�_���;x�pxxH   @y��!�y�O��/.i6k��%��\-��u:�0q��D}Ew�;��	�$�������/��a;D�*������U"v��� �*��A�n������>.ϵ=C ԥ�]��sҜCQ����R��B�
�zX�Ե�/�N����E   @Sy��1�x�J,,A�n*l��5�W׵�Z�{l3h��`}E���9>+� �x\����]�ڼ(��n�`dW4      ��l4��v[X��'�u;?�[��u�V��s��7o�$`�������]W^�yM�<�/���   �&���#��_�;���]���N���<o�;^��*����)9v�K����e;׏O�1@���V�+��P���C�0��Jv���ba��+r��U<����K��������$\ۥ�b]۽ص]#W�{q���N����.p]���i  @s��ؠI��]��=�r��4�v���k�����	ء��4�@�i�J�DQ�8X���ɟE��      �I�z�.��&�I�[���5g��Ur����bp�{�9=;�O=%   ���7�4	�c�c��aY�Ue!��)=g��J���ۻEe��\����S���='�V/Le���8����3X�%+ڋ�W��[����$\�Sw��tAz$���/���mõ]�w��n��v   �(Z������j��F؝K�nV����U��������*����-��MԋHĸ@|�$P��:q�P�S�׬@      �D��[i��x~>gu��ynܸA��՟r�   �3��-�vp9Os�w4���*�h�;QjA6�nw��7��='�3�iHT�spO&��*�����"\<�c�N�����\�v�޲��~���W�߃E�����L]��g/��R��M]�úY"���(p�   ��>dcJJ�W���ʊzza�Q�"��D�Zq��9��+��>���w���|�Yg�>��p/����2~�O\�ɏn�Tq������      ��x����} &�s��崉d7v~����G����)��T#�   �߃�g��5���\���;&�s_Q+�.�R��a�0���R���='�Y�Z�ʈ�{��7n|��a���ʋ� ���N�⾿�O�\޽d��P쮪C���ĵ�Vvm7�Ǯ�gu��M��SM��tm�pՕ$Z_A����"��5�N�3�H   @�w���
e����z"[[�v���	ֳ:��\�u��߿OU�Ѷ�^4V��sٹ����}�֬լ@      �=^�r�X�<o8���pʡ1�r�34���"��t�o՟�hD�.b   �s�>Ů������6`�R]̯th��F"��D���q�K���d���g굩I@����E�aZ�Jn5 mC.܌�Q���~��/�*3�S���9m�A������&�1u�=#�����a��
�v��T�k�ԡҵ�TBrJ�G�'�������+��E�����l8���V��   4��}���j�m��t�
�vsq;��o�������(�~�Ow��u}ne
�{H����~tK��'�O�      �Ʉ�9�IIg"J���ɼ��9.����Y#l7ŵ;{0�{�ӡ1��AP����+�s���5   `�O>�����@��a�������V�l~�v|�pY����DjG��:_�I�1u�c� �99�"�$�@�p�rN!��[�����E�!uP�0w@`���3���m��8�v?�k{��<�_ڵ=!ʷ�ڞ�����ƹ��N��;  �Ʊ��M�W�\c\c�v�~5�:\��]+;�3$^�������0��ڭa��>*�ىRp�
R�Q�JC�Z���,t3#      @�Qgn-l%a</���$�ک-lU����)�e��s��ǳ��|��@�@T����^`�   4��7o��/��@}as����@�<~��z����\�U�st�X\Ԯ�K�ܵ���ߗ3f�5�� �{NNFD��@U�C��=,�׉�V'ǣ'Q)V/�o]T<�����(^UU�k�ؖ"��pm������T�v�8_�Vi��}��ڞ��V+p��F   4�v��kA��\]YQO�7�[	y������h6� ��6�U&�������mpA*��e^O!nWa.��z�       1���1�"�<�3e�ga~`��sx���"��(2��j��y)��3�L���6�6	�f�תЇ   `l�Z{&W�J���f���:oXt�Qg�g�3�����:=q2w�ZH?C�R8�����U�vn�|Ω��rM�*jK+lgTk�Y���m��prtLk��N��<�o���a`9���S���O֑]��kΉ�wm��m8����_��   �&���K�+��]Ʈ���fus֋���ԝ�ھ��}y���芀�Y��^[��G�dT�U\@��(�b��{>���      �����^�+����@7wH5��Y�Y睟a�Um�g�ל����-�q  �����G�1�z3�B��l���T���G}nҜU���9���ỳ�p���v��f-ހ�='��)�6Z�d4C�&:��n\��:煺�Bn߾M��G��U�k���^�k��ܗvm+Ku����\۹��hH>}
�;  ���駟ҫ�oR����\��޵]]���C�Z/�	�l\����6�;��7���0���G��     �t�x�N8�'�b�路�ȹC��Q��2�Z���ݻw	�apvNw�������>~���[   ��G�>�_�ｺ3�B����Eb�P7�����Xa���珇��|ߣn��L>+��~x��oF_���|�g.�ͷ��:�BnݺE���2]��B���@��Ĺ��˩A��B���666   h
��ߣ�����Wwm_M��^D��8�<�}�6!p�GY;lUm��u�J�0F�J.z˓1Y��~�.���       �F0^����$���8����a����'!n/~NT��"v~�����zsxtD���w   ������7���@�����h|�0(ʘǫ4�a�P#�Wc�e��7��}	���jx�8��*.�E��ŉoy����VyE�:��
�f+}����}��k��,Ӻ�+�J���N��|�]ۣs[\e���v�   ��n+˝���[��������.�������m����$W�+�8'�H��	P-:�T쇝��%��      T���)y=/�x'���b�M.T�iq�]���;7�z<v~����ug6�R��%   �)�q(�2�g|��-��7�I�7u��:-q��_H��uixJ��%hw��_^$VG���LZu�'��P:2'r�Q���������|J���4p����#q��k{RE�8.��µ])�V�#��'˔�v�/G��.)�m���\/�ѣG��w�   Pg�R7�L��1�kf��\��ԭ�k;������1�#���-�:�G�91h�T�"���M�C�     @Ua;?��}����j��=�.�͘K�c�~�;?��v��|�;��4L9�TZ%�   �
��	��&0b�g[d-@�s�0�|r����c��9.�����K0i��N�k^��)��!�O��M�
Ri��<iO�k��n{{�<x@/^� P>G�����]��d�U�v��yF�:���ѧ���   j�G}Do��G��ڮy
�/^�^+[�Űv`� ���u
F��p^.�wb�[Q�����\ݻ�M      T���&/.�c�Drz��b� �eeR1��]G�s�,g���������@}9<>�   Pg>|H���	ԛ�xwK�y�a�n���9��4��	ۉ���ߠ���\]�l�H�����Mɉ��χ����C������z��	�8<8��ˇ/\�\����k{X������텺�S���<
���v��N��{'   �χO?����7�ߥ����k�YG���u��tz|L�,�i�W�`T����]��W���NiB�c�q�yN      �^g�z ?H��DD��ryC?�F���w*��]~*m�S���Wm�޽{���Iʅ��g紻w�@}�Ջ��O>��  @�y��3�����@�9=9!`����ޞQݦ�u��E����$f'}!�ݼ�!�K0��i#�"��=d�7e��޼�*���љ��!@������w�R���?]��d[��v�k{���]�)�Ni�틺�\�墍�M8�   �=�~?XإB���L@���q�rD人Uܓ��������nG��9��hn��()~j<@���D���G      �j3]���/VM3Ǌۜȝ���d,�5H�/3%Z��b�ߧ�O��_|A�|N�O p�9���vo�   PwX�pt5"Po���y�X�K����v"}<@#j�bW�B�ǣ�W�ىH�
�����Nت:P%���.�g�&\� �n�a��b;��]�=y/�&����������kT	�UZ��:��A �׿�5   u����ԟ%���j����4��ԣկU>W8�ۃ�U$U۲0�-�������PȞ���~q��s9c��      �ː�ۥ1}�7#9�'M�PN|��yGy������]G�r��w;0��#����#   U��GgT�xT���SvX&o���[Ǽa\7+׭��B�.�-
��5-o������=R'��d5qu�d9���!l7�� �*mC�n��7o]�%7�EY �N���E�*�yY��:Y��j�������+(�n���}��� p  P[~��ҷ�^	ej]�f���`�y>a�j��r������><��ɶx�葲|��Q�m'�!�sX������E����lܼ@      ����M�)�z"��?,�&�bY>�m��e���s����?~L�p�lo�޽{���O   @a$�{��@������W�yC�����=��b��Q��K*?5/o���=��o�R���"ǅ0�-�[��T:�*�Vi�M�����hl��л�K����.	�%q{��z���b��
�e?{�w��   ��r��=��̝���j���P�^D�rD�UܯVW�Z�ˎ��ء����tI~�yT�ށ-�&�3F��Ǫ.a��j      T���G[|Z��V����C!�-΋usa��{��v�1�c,{��!�?_��+����=�  Ԗg�|L�?��@�������~)�V>o���6��#&M�@��~X�ܽ�@����F?3@�'�śS�s�4t�*��*�ȕ�"we���h��ӧ�j�h6k�
WЃ���sm'� ]�72���M��k;���d�2]ۅ��ybM�k{r��ڵ]�<���-��ڢ��   �F�3��uպ��f�u�k�a�e������ת�{�`VW�Z/*��c�����6���Zx��ɽ����X�\]���㓿��u��uq��9�      �ڰ���f�b��o�~� �+TDnqr���y�����J�w��%`���� ?�򴠾�[h~   ԑV��Y�N&t1��P�\�|.K�ބ��J�+�O�J�|{B\���=����o��r��3D�Vn��s���L�L
\��/C�W7o��o޼!P>�����#i{Gc���3�2�1A�^�k{�i/!�^Ƶ}�z��e����^�E������}���   P'����ٙ������8�X�.U<|@�l�ɶ���kB9m�/�$���?<��DN������.��.�      T�w�3j�l��}i~@~���8�ķ2������V��*��p~ZV��0!���ݸ�G��\M'������   �:��΃�%��sr|�9�%�|�ɓ'���a�����J�I�7�ڑ��t:t6j�Bܗ��'��<�bh�U���p�E�*����Si�*�Wm��nӇ~��%޼zE��{�;P�k���òk�\Y��S�k{��]����ڞ�X8��z ���C   ��g?�����X�����nMD��WQpO��f���@�n����Lw�5t	A*�Bt9������ƽ=�$����&��v      �Δ��76h2����� �7$
S��"D7៏r9E�:��[dw�6=	�������o���}����?�9   u������/	ԟ�Cv���-dg����c伡����c��!505���L��^Ȯ
4)n�P�>��!��<J�pZ�\�tW���ӧO����4m�7/_��(ҵݳ�ڮ8�[��]��'���.���܄�	  ����dI�I\��hµ]�Mq���oVq�*���裏���m+����{�q� %��k\?��      փv���3e"��NVS4_P9�e��ù��;(H䮣
�E�������+�s|xDO?~F���{G���o@�  �v0��_��?la&���L�n7z��a�w�$fW�de�۝>5ܗd�w��U���.q]~�Bw"i������Q������vx��5Mg3�[qኮ���`^hյ=������9�F��+�v��{=.//�����   �:�v���_�Za��`=�k�\\�����{}Fm�qm�K p�I�cQi.���=��H�ߩ��ǭ      քv�z�=�'._�����OL�E�T�iO�)PO�ȶY[l�g�� '����	   �l�8#���L`��Jސ���!p98�h;����ȍAvb��A+I�k�� �*�>z􈶷��(x�A۴Z�@|�~�����ǏL�[��[%$O�������뗯�����q᭑�^1��e������~f����Ǥ�ۗ<Y�껗����D&bt�/pš/_|G��W�n������ϩl�A���}���Z�N�Ex<��Ņ��ٵk�W,prr���F�9��嵻���l�.�j�&.�������Eq������eN�p��O��`{���_���kp�x>��<������w�����r�i�S�������ſ�<o��'r}c\W^^����ø0�)$*f�����9�˱=�u�:�</�஢Lׄ4�n�O�����n��M����: -�W��=7ߡ      ��L�^jr�T�)]�Ĺ��%�*2��T-����G�7������ݻ���;   � �^{��5����'�nt!M����@�0��R�0,���z7��`H�9�e�����/����▌D�eǶ��+��~��I����t�s�vEֵ߹���o�(���Έ�M�2&n��?����a�o_�~?y���v�����П�ş�'�<S7�����㿡?�˿�ˮ�{@����Qټy�nݺ]��7�гgϜ�̈́�Lpz��='�����>}J�`BWW����q����=��v��� 8�*���iypy�lA�۷o_�l��ׯ�Ν;��|����g����*E���A]&n�!?6�V��f��/~�o���=�v���� X�q��}�s��3�������5��ؾ*��(���Q�Z[�Ґh.�A<�W��x@�����l�      �>�~�<����'�ùH,lO1ÒY��9��P�W��?�E�1����U<��ڿ����~��89<��̍�����N�N��u#�8=:��_~�of2�����0*��W�������ߖ����9����ܸ̞4ܜ����]��v�9ˮ����I�gggA�M4g
��\�N�y��8_>����Ɖ��y��_.�wt=Ʋ7�G���H�?.���s���]}ޥQ��Rւc�S�S6~qc��ܗ��O����vn5��Ɛtb��ԫ?��w�殐&�b��Ѝ���7o�7�	�"�(�D�J�׉��zi"y�P���|,Y�D}EJv�8Sq��"xR��}�ci5q;�b��9�gp�w�E7o���   �:þC[���`]W/_�UE�y�_}^��ˮk*lW�8�{��=;����,�ܪ�Ӷ4��V��XM�Ȃ�<�����?      jN�Z�g8֏P$�żaXM�FXq�]���jn��Ç�P��ss%<�&�D���k��ݦ�O�c����o���޾|E�7�h˕Q˗_ӳ�����00�x�Dt��?��?��������l�r��3noo�I�M~����igg'0hr�ks&fN�j��/_&*�v{w�ڳ�X6faN�.x����?��?��_��pK���y���{���펽1֋_=ƴ����V�666��})�ua���;_g��V��yãQ3��/����;}����pÆh�]��@��-���>�&LT��W_(�W߽�(\������T�ĵ�O���*)�[�k�'��e���da��=x����o-��������ߧ��o��   �u�g����n�� xl*B_YOe��Wܛ�S��y�~�sUUֿT�g�c{l[�����,�dߑ!yK�v�"�%��]�/�$�g����98      �xޜ�0�'ʄ�v2o��[+���|ar|e����ǇG�	�A������[!   `
ә�_^hǇ�ڂ�?�����������z��W`cs����"w~F�ffdz»�0hR������=�-������Z$�Ƴ]�)ݑ=���]�3��&��K���(����28�r��'��Z�v�̣���H   �����'�������RW0�;�WUpoxR����vm�R��o���G}D���Fu����Ϲ�����#E񀤰E��a����f�      XG�;��g7��{�>o(��!)��3��<OS���U�-2�۷o�{��f&p��g��9��G�E���H   �:�����_��6w����r|tL�O�<1މ��y��Q&yì���=�P������Bo�f��vF� ����58>=*�7h�N�+&� v`� ����{�/7�4��)�hE':�I���TKݚ�3����={�������|؝�}f����}�Lw�{Q��#)�˰��@nP	��HD"��D����f!�EFJ ���c�f]&)�k;�qU�E�x���q�e�.��zX��\�3��������"���� �B���[U�cb��ax�"��	���>�U�~��{��$&������oDG�����`i�}F�\�9 �XEgklnEr�4cqB!�BH�YM	c�f$	��ȍ<�Vdm���e�gA	�n��-���R�|�+���E�hB!q���+��h��1�$�N��Q��P�mM^uC��uк�1Qy�v�XF������ ��,�;�~dn�X�H��AٳgHx�d�Epmr�g�G��X�c;�E�յ��~.J�ڮ�[��3����B)G�;����]�zQD�A����kwC��V<_��k���#���uX2Ѹ��_I+���9q���$Uډ���B!��򢮱���ܽ�kIqU�����X���)�b�{��A|��� �gyis�shmk���-ΧW󛝝!�R�l޼3ss ����4VWVA�a����yM��q[���u��a}�Nա�= s�48�S�*�+p'��Y\I+k����W{��-�;}�8u�L�\۫�O��yl�cP�\�e}����6hӵ���X?>f\"���m�A!��+��ǧ_}�k�!X�k{��Dܮ~�Աc#���d��e�1�T��!�$�u{�j=����RH�������B!��r#UӸv??�]����(n�#��8��P�>VQ�%r/������b�g
�+��~��'�՝; �Bʑ'O��R��p��0��uCE;���qܓܕc}eݰ�
�_�®��(�u��6{�*w���L��xg&J*F|�A�N���X]嬫0��ۭ��u]�AZ.煸������͸|��fl�]�n��һ�;��_۶m�r��B��$uU���݊��][:y�zq�XC��j��=��&c#� �JT��T�W��>�Ȏ��`O\YXYщՍQ[H�tW) �B!��X2괄�m�`/p�
��
�8����z+?�cmq��� �!V��{� ��gqqͭ� �Bʕچ:$	TUW�l|&�s
aP\(�Q7tO'׭fb��z/ݰV�0U���$*
��7���:�c{�vHUr7Y"G���м�ܒW�}b)4��ųg�@J���������T4�v�Ūr���p�XTZ�퐈��v[�W�����XY�[�������3����A!�����*z�}	�K""��)lW�W��u?�y�{�)l�+�SI8�	Ư��
�%FϿ�p#n�ds�H%&������';i^�1�m��5���B!���bj��ƺÚ֊�pL���J�#f�+�_��R\k���+?����8H�03?���LOO�B)'�n݊�	޷Tc���x���e"T/��!�1V��åVˬN,��:���/�P�������WQ���ȴ��擬N~E�P�z1��СC������o�oX�k�LHO�|�؎ߊ�sm�}8c��n�K$�ر�%B!�ƞ�/㇟��u���҉�K%�74�����U��}I��0?7b�������x�у�+��j ��{=^���HD9U)��e`��vB!�Bʍ�y�)]q����,l�'��H�s�)�¸
ԃ�Ӯ]��e��Sx
���ql5�P+���<Ĺ�'p��; �Bʉ�'����wA*�Օ�Nπ�Þ={�c06JMQZ7���t��Z�G�p=��� �U�n
���Ԃ��E��*8�t��Pb)
���0�����p$�1�ߏ��epm�]��pmw��+��um7?c��˞�k{���4Rx饗02BWTB!偘%^U-�7˵ݗ�<��� �T�ך��bGy�*�.i"�JT�,[��p_�j��[|b&� ����|B��w��T�v\$�B!�����$�HL��j��U���bY�V�b��`~�ul��0Ƣ�=�+��O`��m ���e4�4�B)7j�밚H�T½=
�c���M��o��ڻ�u��6W���̵���^E��)pHuCR���v�_��q��zJ�U����[�J8��������W�\��	��q�>Bwm��*׵��66>�3g���w�!�R�8q=�}���CB{P,D�q��ũb��)XW�l�ر�Q���*Q'��ݯ�r43W�Zلu�0E��r�\̤UcS+�����"�B!��YJc�f���ܽ�XN�sl�.r�c'�63X��ݤ�̯���o��$&��(p� �fg�y�fLNN�B)�����H����Hx���+�n��<U�P>�]�9�M--HNUnݐ����޽4�����u�1��:Kc�Ų�>S&N���t�رȒn�HwW��-v���s��[{4�J�ڮ)lõ=ݳC�n�K&ؼcgzyI!�!�B��������E-"�S�T��K���>�~���P2�W�����c�A�����%9n\]�rQ�]w>��K؎�y �7��#�66�B!�R��74aq~6��i�%7xM�d��'���C�r�-�j�J�ё�@*��~ƥ�g��g��B)^;�:>��5H� �IxD1��S�0���&�K��'�L��m��U�(p�\�u��K/aeMRy�ܰ84��.�jx35�Ll�ݻ[�l�r�!�������ع#�k{���q$�k/q��k�뜊����n�K�^����{�����Y����x��!��8#܃�bk�s��5��ب�ŏ5�o��`]q���+�LT����x�ȑ؈�u�wN����Ð��q'����
a��9�M�{���B!���$U״v_?��Ȫ]34��ng�Љ5�`X7�Y�p��&PzN����0Q+���467�|�BHY jյ5H&� ���?��i���JQ7����w��p���� �a���:Wzݐ���Wc�Y��tn�ۭ�n�� .#�/��lm������]��s���I���� ���v�ڙMf����Cr��ҵ�޴����vm��Q��k�����65=�#G�P�N!$��=����wD."W��Ϋt�� �T�����bĮ5��p�������8��r���m�hD9ݰ��'�K��<��7��*^�B!��#KhP��k���-��]�XV�AI	ͱ�Xw4W~nll���H�YZ\������A*�']�i!�ӧOA!�ę׏��_�>��&&��X$��� (i��E�ZU7��)�c�������k2��M�^`)���� ���;a�tb��JD)�W�$��=J�{��tu���鿳�vG]�m��q.q{	\��q��:E���������4!��8"~����HZD."����9��+���Ǫ�U[��8�Xk���0Hx���k�	�&��֞��4�ݞ��cv�DU6��pu]�(p'�B!�,�X�A�b�&]�,U�Њm�(Zk�V����k_KK:��������Do��y��Bbώ]���Jbt�u�0����겏�#Fף����p�=��=�w�a��T���Q��ܺ!��[I�ik#�	������"����3P�h7���<��]�U�\n0\:�>KO�p9�4]ۥbw��Z*l(��\�Q�+�k����s�+�k�3nxl.^��B!$�����\�cu�)L�|�v�� �T��A�P`�?���A����Rn�n��L��}�����yU�������&+7IE!�BH��b6�v�b��G��8�ǲ���!�e�B�z��b~�ū��J�{������� ����Rz2���<!��8"���fi�Xi���IxR7�"�5E[�б���FX.���~�k��B�t��E�����I�D�ډAqa˶�8�C���d����^y����NLL`۶m���]��b���n��\��P]��m��K$ص{Od�[!��|�;����y���pa����b��Vչ��F��w�1%��T�#� ᡚX\N�
��	���cҊʅ!7�ϵio��������S3�B!�R�N�prs��@��zM�������1��@��^XN�W^�X7
�*����gN��/��:!��xr��Y|��]��b|t$<��Y2�6��ۯﺡu��mR�ӭY2C,��]�7^o��o��te�)p/ɚ��jJZ��ve�� ��92gf���� �09K<\^t��������{��[���cG���cB!q���ˉU��܏�=��\%�5�)�rL��=�`
4������b�E������'����7�VM�n�q}�	�I�M\�B!��r&�v_��ڊ����_�,׸���6/�^��V�����	�ŵ�{~n-k�:�����m�BH���55XY]�������*c,ʡ����U��UՍ��j	�%�㦶v����(p/3�z�).8�ŘW����賛K�j�������}���8v����;�p��������æl*�k�zlY��{���mF�8�b�o����|<5=��^{�wB!�����x������\O�n(��/�XC?V%"�=���O�f�y^#C� �!&>�r��$�˶�b��5�Sg�w�,5��k!�B!����o�1?o���4��Z��qG��ݺ�ڇ��Xn�W����W_EMM���^�=LF�F�r���J�yowZ����B!$N[�|�����B�"��8.&V��V7�����{��S����z��KoW:��х*�r\h�|�s��q�ex3���D��
�NzQ�.O��Y�f/ĵ] �gv��<붧�]�]}����˄�A\������
���.�3��󿅁����@!$n467cee%�8L���]u^��������X�K-Lp?��b�c}}}�q98+�"�ב���8�O:����I*�C&a��|R��dB!�R�,��6�Uo�`�p��:k�Yr��b�u8c�(�[�lI��?NaSXAсï�T�{��浛�B�{^~|�	He!&\���X��}6�
�.e�u�mF�qzn��{�d��Y����V�
����)�l�̢(`�A��]'aeub��G��E!�+1+�����"FF��c�N=�v��Ј(����ID�"xw�����*�u���ΰP\۽D��F�}å˗�ч�B�G����P�q�"r�
[�S8�����P� M�z@��y���bl���_!p/&qOtY�Rִ�r�r/�K�]KY��B!��7�+5hi���A�Vl�Κ��swPW�"\�)p���A��c%�@SSS�nL!��a�8�0RY�����Hx#ⰈCMѡgϴ��9 ��N�2c,�6�$�����.�а��^��qq�n�<�r�t�0�C
��'W�|��-� ����Jܵ]��jC"�N����8���cU�v�!�k��+�gc)]ۭm��v����k7����?��BH�>zw�>��R��"��\�b�4�)�+}�
��/5��^$�x/.G�>k2�㞠G�sr&�I�J5�<7n�'P�&�L��E��3Mq;!�B!�Nߌ�W٪My�	ʱ�z2�5ga��k5ȉr�f�P.�򗿀����"f�g���R9|��G�>s_ݹB!$�=w�>��������MJO��q�)�8��_��~��Ms�B�T��ɣ��"��܊��i�������� �*���%�u�t��y�ɑ#G�i�&LMM����'Op����c?��6��C�]��*{c&�p�vg�/�v��8#Pl�:��6C����ə�A�Yܻ{�BH��ر�33J��4۟0\����4����y�Ā��u�8_��4�7 ��88$���0W"t��6��^cxuK����؈�N� �B!���N��M59a��K�f��*�U��F?y��q2�
��Ƶ��Q���_X@k{��!�Ă���6�ayy���{{��q�X1+���a��4ho+�k��f^`�����4Ƣ��X$j��2����)(�e�W�ʌg�K�I���Z�8q��9H8�<�J;z�/�R���+sm�v{<�P=W��r4�]�ak˵�u����#�6��:|��B"���s���GW{iD��*v��^� �c���u��c}��}	�s����Ƕm۰�~đb%�̱��M�y$�;2X������B!�BH��\��onk��kb���"�е��1ctd��k�AꇢfXWWG'���W��T?���O����B���gN��H�120---���͑��P����U��f(5�b�0�Eb>U���pc(l�_��Ȋ�s1*!kT"t?�
������H"�@_��]ǵ=���܏`]*:7�򸶫����~����킢����nH�W���'O�>!����XY���K�NDn脭7_�^
�ZDP����M�󘙚	�ӧO��OL��P|,��R��>�&��ݜ"�d]3!�B!����{Ø�Nn-�f�[^3��#菵�ʤ�h�'rG�U�~	�ѡ���V�y��adl�^}�wB!��y�V|����Bh��G�@���ɓ����>�Sݰ�5E��=7��z���]O�r� Ǻa
܋��Bv���B������a&�T1��C�b�N��K!ɫC�������Y�{9���D��vm�ƹ��7�T���ؠ��p�NNO���S�B��KW.�g����������avX�u?�y��*��yP_"x�dM�� �Zf��LV��s}�=L뻵R:I*�x>Y�vd.�M!�B�F`��q�^?��઻���laݲ�c�O��O\�pq��=<Lq��/�T��}8x� ���@!�D��c<���P%bN�$�!��@duC�x;����˚+X��bR�u
܋ĳ�$v6���0���$�&IV�b2��>�quW�O|��%iV)<}�o����]�a�Q�#X����8���*�A{T��n�W�����Z �{Umv�܉��!B!a"��������j��X=�u���"�b��W���C������=T���Xf�R�%����O��'�e�J{E�u��HT��|&�!�B�L�Ԡ-eX�d���@5��.n�aH�*��A��C�-	���!
�+�g]�x��-
�	!�D�������>�<��Y
�ÇK�����[�P�����uj�NSm��.���X7���H̯h�ֆ��{� ݋TZ,���N���!d-w�'Bl+f�?�$�����,��۳me���n�q.Ѻy���smwoxt/_��?A!����K���I�D�Je��)�=X��k����Ep�X_"x���k�߇��R[[��^{-6���gMPIw�k��=�3Q�˅��3H;���B!�����I'�r+?�c��-JͲ�cG�K'7��B�	'ϸ�47*��8~�H�11=�m۶all�BH��ڵÃ ���"�W�P7�����a�I61ݭ�Ͷ���m+�Y��'(nP�^Dj�Z��<f��dK
�Kz�`��q;A�~VK��+�ŝ�p�|։�����.�������j"l�vm�r}��pmw�� �D������bnn�BH�ߠ����������@�v���� ��<�`]3Nլ+lwƎ�`yi	$<��ݖ-[���\*�>�X��ĐW@R�ř3him��4U�B!�lg���RCV�n-T�����c˄���y&�
�!M~�С��vtt$&�'����ƦF��⧟�֥���Ï@!��ɉS�����T�󘙚	��{���_�FB���[k� $cv��]U3T����1ɺa
܋�bU�t6���ݙ����Y����P
]��P�}���3Hx<��g�;.�wV�g�vC!x)�k;����Nq{�]��{7<6�kׯ��w�!��N�Bw��5��\���4E-X�ӿ�|=���ՍU�u����~�p9y�$*���1v�gfC5d�:r5�m �B!�l,[ڱ8;��甬 n/������fX���=&z�XUU�W?���8q}D�mX��~� �RY�ﶕd---���!�����P�4�>/X7Q���Ƣ6�*�>7��a���;#�5򜑵s\�e��J����Y74����/Vc�5Ie��N)��.�[���YŴ�>�ŕ���_G[��u]]����}�D[}�}�}���OP]S�~\��������O?����&V����;3�����ӣy<�gD"(W���U�{�������̿r|��Z�~��)�����<Z�[��ۛ�.�p}[T�������#�{uu+++XXX���ړɤ���1�����_Zw����f���Td�]�u/�w�{#�(���W��.�HDҿ�[\�Q}�}݉����aK�Z���]������Y�}��>�G�����ޡ;�:���8�������Z(�?��%�����<�W5�w��7�"Y>���%Q�����:v옴����V�}�q�z�{R�鞨?�ݖ�&�ֶ4��PB!�BH�HԴ��&�c �)��v���	��M�����n3���Cq�c�X����>�_jjj"�_���k��� }����=�
z�xݢ�����(X]Y���rd5�d"�k_^{������ĩ������~��[-E�r���Gտ��ﰨ���������BT��(�;�]������wͺ�$l����5�{��>�gΝ�W�~�D26�}�om���D��X+���k��}+��t�[���7�O��ߋB�a<,����k��}�nN��g<��v�4�r�E�ruH��}�ʘΉ������Y�nVq��b7����*k��mSUU�$���]�+�T~�r6�����ňn$���w�ٍ�G��$��P�����_����q��vm7����϶�rmw���$���I}�ɧ�q�Vd��}�	n���3%�g���~�ڽr��o���!l޼�!�<p�@$}����,v��I�bB¾}�Q��B`.~CĵQ����� 777k	SKA��]$����#[�kpp0�sT�����mC[+6@��\�Ų�{��)�Ւ��}� ���N�W���"�z�O��#���k�`jb2�����v�yyT�^������Ͽ�.Q;E��ԩ��y�pp/��Ai	z��P:��Dn�U����R��|�{J21~lI�gVA!�B�8L�֡�HI��~W�2�2I��	��5i/��Za�r����bbLU>M�M#�(��E^H/r���\ZX����`a~>�y�J�%���'VX���os[�&�~bGQÉ
!8�����{V,�~��_�3Ң����Q�k7E�Q�����wET�u�yT�]�-��Q���|�b^��~���c##Z�������B��'#��[Z��q�!�wĵ_,R�f�g��[���7��Q]w^��[�P�ɟ���&����.���6�,�;�n(����L.�м�	Ʉ{v���E�R^��͒���L��M�t���=}�tAn�p�>~��+D׆D8-�{�U�3q��*��<��nt!�W��V�~w$q�;���+����m�v�s��)l��󾯬���={�B����B*��������0�X=�u���"�����s��С@7��?]a�:6�6�$\�d�W^)|I����y��ڱ�S&�MHώٝ��+���f���d4MB!�BH����]�ِ��c���:�q���Xq���w��ق�4B��1��[1@~(�k����K�v�\����=�qʹm�@sDF-bUĨ^��Zߵu���O�V���ĝ/��z�<��Y�5S���znڴ)��+���w���i��(��s&��!�0�پ}{d"o�;�k&4bb�x�Q�k7�/�u�7������$����}��h�o��cwa�ܔ{����E|߶����Ezr�n�Q�ۛ��,F�ޯ���"��
Y�pV/�>�k��f��ayk�5��֟�5�	QA�{��oj��̤ˑ���>�%������rbv�s6�-�*iu��)
�C�������븶kŭ�۵]W܎*�Ъ
���^q�P\W؞nUL p�i�3{���;�F&�p��M|��� �BJ�,��y��v�����S���k���\�׵�J_��p9��kr��r�gx\��M��Rmv1Jʐ��S)�s��[�'��"�B!d��;��k�k������]�.���1F2��������ҫ?��� �1��_����7B����Bc,B!%���		#K�0	����p9w�\�Ϥ��<k�^�r�l9֚!�f������������c�P�^d����.�q��
��w�Ju�g?$�f�ʗ���*��
s��������Ȉm�����.(o�v�ݩ'�'Z׉�OѦ-n��2�v�+E�.�7	�=;v2YE!�d�;x ��p���GX�+l�4_�4��q���v?�������9���'I����WɈ��zq�J�a[�{�aMd�T��Ĺ����B!���Gr�~����s9C,Պ�V�6e��^X7q	��Ͱc�{q���N�{���σT&_}�-�_��/���BH)�|�
��p�r��=l��pe`�f���(Y�ݡ��S�S^� ��X�H
܋��J-�,�jg�ZZ�NɒUގq&2�9��t>=A���A��>}:=[O,�C��ɣ�i�����ϵ=�l�s�R��pm�ŕ�k�3ntr��x��!��br��I���ݻ�����}��Op���U�k`���1}	�5�T}A�~���L$<��މ'B�/�}����=�?^�u`0ۗ��Y�B!��-H�����]1nH�
้��L�l�w3���se�6q��s�pp�1V����afz�� ��pӭk�Gcc#���@!����,'Wi�X�L��c����#�U2�P�+�>Ǆr��Z��~��c�o���d��DMH
܋���NVIfWH�U�6庸��*+�6I�*��7��y(N�J��Ϝ9�/��$<���#nܾ�%:7��m"s3n������ڵ��~��u���θ��U��s���9��BH��Q{����g\���w�avp���ؠ"�u�8U�Z�����{��A�e���8v��\
�O༗7]�w�:I*��==q�>�����ZOT���@�B!����L��)y�0�����2�aH�t�C�^�z�}�fXSS�D�c�0|ч���A*�o�����.�O?!�RL.]��/�}R���L.b�0���*�ڠΊ��ڡ�nh(�#����87����.�N�ցu�����.lopϮ��#Y%��B]ˇ�p:0YA�I�M�B,�A�{���crr[�l�4d�rq���B]ۑ��µ]7�0T�b�����[��_�B!��>s�=]�u��X��ZҤ/�Kخ�U��
�u��Kp�>p��/�K�bYk*/^Dmm.E��RP��v�N�q����*^�&�$B1Q�B!��1y1W�����c���X�%z��q��l8��ȭ[��'q?|�$<�zzq������jkh�E!�����bae	+�� �K��p�����$�_�P�;|�y�v���=>�������v,�NggZ����\�:2�Uָx
�K�� 	��??��פ�s�k{�ܹf���l,�k���һ���S�i���z�`]ߵ���.�Ov�܅��6��΂B	���ڵg7����"B&���g����µ]}�c}	�5c5�Bܾ��De�qHJO4!sa�?&�wU�� �y����Q�N!�B�F�s"��Ȏ�u�|�g�c�<c�9��YV\j}A�99{�,�!39>���9�X�0�������|�">��B!��ҕ����; ����4f����ӧO�8q2�r���G��5C�����sʜ��m������Jd��I������ֵn2���ǒ�̝�D��!����KKK ����?���ktm��C66��w��K��nA�ܮ���������_�
B!$�ϟǳu�v;*�^A�P>_�W�X��\S��)"Wӗ�^3N՗</�z@�E�?~����>kj
J�v_����w��{s�`�B!���j�@s{V�uC���ڡ�.���Y����ns�8	�i��1������_�L�W���ʸ���́B	B{{;f��Ƌ�r���y�U�=}UU�����j���f(�*r�MH���朼�Y;\ۚ�:����@T
�����:tH
�Ra{�����]X�aKT�	��pI��9���'p��]��x�ۋ�il�ؔ~l
�]��R����������W�c7�k{����õ�~@2�D��m������4!��B����܁�.�v�[!��\�+U��Y�v�SRח`]3֧�^���_􁄋H���	���t�槠vbp?G1.�LTW
U��z�ru�}�	!�B!eGCR�sҺ�z�g��!nי��^ ȞBf��ĝ 5L��.�M��A£����
��{���K���A!�A��t�s�ʦ��H���ק�Sq�񕂜P�ږgܭ��j���1V����%��x�kSҋP~�z�܀��aG���Ǥ��,���r��=|���8}c�ϵ�&{+��u�ܮ����.:w����,�k;4��;��z��@!���k���E!�V��]M��K[5�J�\����c�����..\@]]]�q9'���!+j7���*���Dx"�ԮJT-���*!�B!��d��˙-��������1VX�Z�c�ر�'O@�cblK��hlj�LV	�$Wӆ
333 �B
a�֭����d�
gnv�SS �"�Ž�IX��(�κavlI��f��S�񾗸]l�+�k=r�
+����Zv� ��p]��V}q;g|T�wy���q�e���jߙ3gBs�'9��.]�\|�v��Mi%���%lW�mD�vY�vmw�'D=5u�8p� ���A!������M��<�:�h
ƃ�K#���+Ϡ y��Ԃ{�� ����>�Ν��3a��{�1�u,m}N^��c/[�-;���֘�!�B!���*u��X��.zOIk�^�XY�B��1�}w\j}A�9�)p�ߦ���z�r���{x��u|�� �B
���Kx�A*���^��9��vl���B�9��.� U�;_��Hyc)Vx{:Iͫ
�KDMSV�G�3.d"w�s{Jq�{$��[VPk(��a�$xQ�����mmm���,Hxt>}��5�ڶ�L�!�ѐ�����;�%n�ĕڵ��f������v��\�u����;cG'�p�����p�	!�_�z�6����"r��Z�d���ǪE䚂��"x_�{?�����h����Muuuz�W�u�Iw�ò�]��6s�nNBw����Đ�����nY?M��}�B!���N��*�o��Z�9;�P��������X�:FPs�BS�~��i����	�ߡ����i}�C�`?z�ihA!�G�����ԝ���n6bl%�U������k��K��9��ݜ�w�1��f(�mni�� �N(p/�h#7���\��}9��L�?G��)�r�~���>-����A�嗇?���˱wm]�q��������g��ݻ �Btعk��f����ڧ��������XC#������=b}	�5c�7SZOW����A,--��ˮ�ϠH{Q~I)�~2������`D�[*�R�k�T7v�B!���1�*4�n��씭^�9vȎ5�.�	�y�f��H�ެ����F���]�t	����7���������R�<�|�߾�z{z)P$���0�9x����G ����&�'@�E��~��ٲ���ϡǵ��}O6W������ؼ��%��\5�(�!�.;`���R��UI)�D���6��e�&�T��Ν��=�~�-.]��h���+��ݍ�8�g�v�k�@��θ��9=v��	+++ �B�q��E|q�kW���Ї0�8�u�8�X��{��vu���իWm��qHX����r�݉�֖w�+���8r3)Q�!�B!��rM��X`B��Tܞ�j����9\�ӕI�PF�k�^X���с�'O��o�	��������@*�����3g���߃B��¥���ӏ �EW7H����M�Y����vh�*�堮%Z5�*lU�P�/Cmg\�����D<M`oG���t^�v'����r�qHh�x1���O_����a�m��qrm�	��Bt��%�vq���|�����]�!�+��oxl�n����B!ċ��N��}�Z彟�`����u�0E�rm� ��^36��[c���zzA§���X�ڧ�^��&��x�D�غg�q� �B!�D��r6)��ұ�ȇ�P�\�Y>f�b�w2[��Xs��,��p���w���7:���^K��Nc,B!�hjjBcs3&&��M��'�{@�G��k�^X���v�p�to�ku��T�5k�K�ء��D����v,/�ۖ�9�e/h�,_��DUF�.v�~�A���^{�5�޽ �������mM7���{����3t�
tm��IK������ۛ�smwƮ��b�Νزe&&8� �"���/�ۋ����m���f�J�.��F��US��WDD�P���ɮ�Z�_�!��{؈�����c���8���xں��8���.�[��ּ@MM5:�WQ�	�B!��x�h,������%�mL�{�|�Y\�X���`���\#T�;}�4H����anv�mm �͝{����+��OA!�xq��5|~�k259���i��Qǳ���L��V�j���������N-�@��
�K��Ў�ܬbօ�蝛ɑ���)��־d�*�{��R�S]]�^.��#H�|��7����6�h�p���@۷k�K`noL��Qe_� ��|m�4N!�7�?����~b�q�øy�6����B!D���7���/鿕�����RN�
[I����
=�] �s��q�ر�3&�	+���'���8���U�b���}3��B!�R)L-&Ѽ��+�9�+����v����w�=��y�2�	.l/A�hlڴ	SSS �"\�_;u��Y\\�J2Ac,B!�l߾�s�\��}�>�v�±c�bQ�Y��RS,���*c,������S�ˠ�����ԣ�Zȶ�eEoC� ��eq%�r�&��qHh��@�{����ap`�v��
�%�k�F�[�^t��u7vC3�}<�bvmw�K' �vmw��NJ���j�iU:���NB!V���Q[_���y�}�R��`=�of��ͥrm�=Cf �����~��˴[٨	+�3'%sb�?�˽]�(�Kr��- �B!�T5M�XYQ.I.K����O�0�a��uuu�x�"�{�=�p�������������[x�wA!��8����C"���	�+W��W6���U�}&�ڡ�fX��۩�U��,�4p�+����)�uñ��b�A�����5�U�{��z�~�K����˨��E"� 	��~�	;w�;E�R�q��=�k{�/k\Vd�+X�'lw����\���a;�1��A��;&&'q��%tuue�S!�B�o\���?h���ڮ��{��]������j������B�.v�}^�+d_X���=�[-�U�Jm�I�#�k=��B!�R9���v��b]c
����cK�gѻ�R�>��3���Ħ-�A*��=�Gc,B!R�;�_:�M�Fʛ����̓�ϙ3g��q��AZ;t�3M^cn�~���i��z��;��D�Z�Թʠ����M'p��iA[v[gpd.�TZ�.�px�JTY�K��`1����;w��ѣ���A�廻w�߾��˵��h��rm�;.�k��|1��a�yč��.k�����7��'��B9z��H&��J��߬�߂�f����q��k;�b���ݝ�A§���ϟ/k�=8��ck��)�ߪD�s»�:�I�B!�T���ؗJ���e+>\�Y 3�rcdk&q�r�����_D��=��4O;���7ޤ1!�b��}����>!q�H�G8�_�t�,�����ܣ�@5Ô�_�8����p��9����ж�S�v�l����B�������ڵk�G���4�?��GC��.C%n�=���[�@�n	v�����
�!�X��%�)�o��Kس{�mۆ��!B�l���q��Q|�ݷ���������O�k���Bjo������0H�\�z�����~I喰�`q1���%�rb��t�dv�+csk+F�� �B!�TO�8���=!VR���+?��1N\m���n.�o��E��A�F�ݻ��� ����'Ξ.�$zR�|u�[\�v_|�9!������o@�@����y����*v�����❃E]�z���\+?Kk����\��P�U�9f�A�{��C�R�YQ{\��~w���]�*����%Ո>���G�	���j
�ڮ�]�.��G̸����ѵ�y���!��7��ÇA!�����m����\�R�]�߬�ڮ/�WtԵ�G�����g � �K2���P�c9�R��3�N��D��q�,Q�MR������M �B!�T��ܱ�3�Rw���l�m����i�%0�@:ò�8����7o�w��H�,.,bx`;��!3��X1رs'���A!��ٽg&g���� B�}XY^	�7n�ǽ����Cg���果�Q3����Ա�(��*(p/1�S�x%�t�u��-c������nXE��$��+��rHZ�9s&�=::
.�����G����R�q�v���a��[cumw?W!�7J��.i*����ﶉ�)<x��� �R��y�e�,�aii)Ӡ)��-B��TDnh�>�+4���⸶ku�!6���>b�A��U�L��G��\P�-HU�})k�,a�tfL%1���tp'�B!�Y�i[Lz���&�X�9����Z3��I�_C���/\��������!š��9�$����۷��7_B!���g;y����bҽv�H�G|/^�����<����O��v�f�|�ܭz_��˹��|U�Z�)9���g�xu[�2Q����3:���[��������|���U�sP(V?����~�:���?��K2����p���k��ն\۝q��yqum�[��mn~[�oC"����
!�T���8s�Lf�A���L\�3�
q{�#��5�_k9����a~n$|�?�ݻw{Ɣ��]�a��[�{���g�9(����<@2���q�0B!�R�����%�[�9�P��5C���j���1�#[�0�[��".��+W����333 �������hhh !�s�݃�k'=BH%s��U|��=b�Y�g$|�oߎS�Nž��2�Eǘ�! ��VTKY��)�ڡ� �g�������F�:�8=�JT�_�ܾl�5a�w�A��;2�X3��ﳾ�D��O�SђpD�����KW���umO���t����� �v�u&��Xw�8���>sS�Ӹ~�>��CB�,nܼ���vu�V1\�u�TD�K����
���E��N�h��V6��=_�E�a<T����2��}.Y��҂��!�B!�Ƀ�$~�^%��*~K���J�n��r�X&z����uㅸZ���}�]�p�q_w;
B�cc���CGG���A!��زe�U&��@�I�����E�͛7�F�&~kva����׏EU�f#��z�1�}R�uºs|�to����ӱUHœ$�!�Pպvq��MRً�)�Ca��+cm�&���FLZ	�HX---��K_?���c���cma{���[��pmw�\۝�b��rr�O�Ə?�B!��֭[�Z�ᚙu;u�Ƶ�_���Jqm�s^��p���++����1X����p���f؝�������e]K:Vqkh�B!�BH岚4�ھ��Z�v��ʶ�y�C�9��V(#��C?�/^��="��>����x1Џ����x�o�BHeq��U����A����.�h(�n�7>NuFk��Y3���녩u�j���c��6�oEr��v/(p���Z���Đ�[���%�Rz$[�ʐ�z���(��զM�p��y|�� ����������Eumϴ���~�9�D�n����#��ڮ�ƾ\�3�rq����,N�8�G����$����cW�_×�~mk7J��U&��~b�	�5�T}iƩb��p
��=G2�	�;v��2�A����ջ�d�-9eMbI�S�Ñam�2��z��;!�B!��r]���`���f8����s?"�,ֱ��6��ʵ~(��jjj������	LON�c3'~������c�8y��!����ܹs���O�����gld��3 ���؈K�.EZ,E�Q����=w荵���c{���U-��#��=������2J�7ð'�d����55;U�����F��^�~���)p��o�|����ۨ��˶�@\n��\���vC�\����hS��u��>���;��zWKP�OA�^$�?4��׮�?��?�B��F�={b�E(�k{i�tm�3�Z��=��A��\�,N?�e�$��{tD�V�H6����u`�nI<�`��B!��Jgp�[�IW�Pe���:W~N��-�-�1��0݉�
΅k׮]8y�$~�����~��/�!&��8z�&�;���� B!���4��a��b��Y'H4�U�6oޜ}\��A=�5�t�Ϛ�l�m�S��貚�������sB�Kc,/(p��Q��-X��T^�r�7�C��ڮ��.ITم��s�HI��W��~=�8�D�p�3��T��Va��;�urW��%m
a���zn�q���nm���Rk/��S���O ��1ٶ};[�1�ە~L�v"r_�u�8U_�q�X?��f���xz#�Pi�
�q�fқ�c�9+���Z���M��K !�B!�΃�q��*i�P9�VQ4wn�X�B�cE��^�c	w
ܣ��yN�;�jO7Ri|��W�}��{�]B��ܸ}��1�������^�h�|��vlj��9�e�l'{���:&�kcFzu�ǣ����X�nY�8��I*���ʍ!�pf���	,G��I&�.��ڀI�W^yǎCWW�������%������Ghjj��MMN���3WlZ�G�n����&q�����]]Y���:mq;4�MNL�ɣG�P�y�N���_����S5��u��&#C����M͙�aۖ�X\\͑aii	��ш�V֮7�:�n�a"�+�򽟟����F��ƣz�(����9�����!
�|�b����Ey�WWWG��#����I:|���ct>���E���	�ڃ��/�/`d`H+�Ϗ���}a�����K�a�����|<��q��E����C�*��U__�.����7�����Q�13����)t���M�Ei�ʑ��6mںvSB!�BH����Bk�&,�Ϲ��b��]�9e]�\��ܬ�X�T$�1S�!W���6���?��?�����e�����W����U<�|�S�O�i�E!�s����_�uTB��vu!�J�o��ѕ+Wʪ6����Cg�����83^wX��ElK�f�N����虯�n�l����� b��'�����������^Du�7n��Ӿ��� ���³������[�nͶ��ա���'��m����U�׺\����l��D|
۝m��%�F!*��ԑ7.=�U�q:�?ѿx�U�����֖Ʀ&4�����5�g%��_��&>x��P�QN*�OM����;*�{�ｘ\ ��('4E)x��q�E=�,���D�������x���������GCs�4F{▲����g^�[�N�R>[[D��x}�ucSc�X?��oU�����ٿ�`��u��j�
�T������U�^4�{�8���y^b�������R'��Z�0so�qiQ��wmw�mIT+�I�YC|7��:!�B!��O��}m�0#]�YV7�������k�"5�Xg[k
�8��\h���ɓ8p�@��D�ӢB�R�9G���w=y��E�&�{MOLF�W������,j뢑MLON��i'�@����I������ً���qP(�OO���Q &{���"�?��u�hff&2��(_�����f���龣�WG�ދ��0UQ�ϼ����o�78j��KKi��dD�
G�;u��l�~r�+��mog7ZZZ������{N��G�}��}ٿ�8؋r�z�ˌ�UR7�cV����I�)k��CО[�-�x��$?���/ëػ�Z����ڐ�1�OPْU�$U&�S��:]���V¥����m�ė����s�AT����;�=ë�_�����'himŎ�;��Tn�ra;l���vK��z�f�]���wm�~����Giq���һ�[�����?{z���!l߱��}ss3�������_�ԈH��+LĄ�(����Ć�6DE��H��6��>��Q��"	->�����k��bBUT��$��;��؎;��ц��zt4�ɺ�m����Ԧ�o�7m���� �����Ɔ��;Ա��k5|(��؆�����v�4O@�ZU���d
ɵ�����yU��_�de�(���п
�y]�~]��qpf~��o�xٺ��_g'�����	�2���9U
�	!�B!���:t��d�>����+J��C[�P���a�%����V��K�-ꆿ���\qQ	�L�IT�CAX�]�s��lڲ9���م}�"
��ж�#m�Btv�ȡH�^^\���8v��'����]|6������o��_������NOv�Sؾ)���(_{��������UD��E�xtt�w���~�ܹ3mQ���OL.ؾ}{$�G��������_�/���q�5�߼��	TUW�csD߷��G����pZ����}�5>:�񱱒�CT��B��ؘ�����"�EV6FmP���U/��f�w��f��f�����༐ns��|P���ܾ��S��v�f�ܽ�� O����_G�&�N�>��_~/^� 	���|�����.'[�v�8/a{�5�Nw�_a���=q�?|����	������/`�� zϞ=�A-!��򦩩	5uux��ܵ����ԋU��5���}	�5�T}iƩb�ܛ{�>�$D��֭[%wS�S��:�0Q�:�e.=�tWt����B���d��9vB!�B���X7!�����e��k��TW{�����Zfxe����ʋ���~��߇"�%n��>���A��y�s�\�r_ݹB!�}���o��}����S��qㆴ�k�������s��V�,E��1����h$?���bM��:�d�-I%)��
����$��%���P�Ф����7����˿���X���O?���\�*s������jm����S�i��%q�#g�İl�R���
����ڮ�?4��7o���?�g�B)_~�֛����E۶�Bq�ր���rm�o�!��:��ˏ�}?�5�V024�^�D��˗�u����%���������/nwO@WNZ_���&��6m�1Jq;!�B!$��������0/]J9�Eu���=~mrg��~�������uD��s��u��El۶-�dK§�yN�=���hV�$�ejz�+Kطoz{{A!��9x� ��3�fg@����e����}T�ݻ'O����|�j��14T�y�8����LB��z�]۷�M[�<ŉ?:P�"�ӵ؟JJT��;���0h��q:��?�z��R;5���n�G��|���~���Ɋ��^<a{fO�v�c��vm׋�o�~��_A!�<�p���v#�v�j��-�����#��=�N,]�����ڱ�̠;�LP鎩�"vU��S�nYfp"%�=�dNB!�BH����fg��C��f���E�.�D|��nh��+�������o������I�&��;B����!޾�&������B!�X���#���矢eKq���y�,�DÛo������i��ceƀcP��W��2>�2�2Rr��bm���������k�ASخv���l��s�����V.\��]�088>�}�x����ۛm�k���@��|�����*�X]]EuK+^�u���� �R^lݶ�mx��'�8L�zԮ�b}	�5c�
��k߷��--.��.�QWW��7o%U�u���+D��ڲD���������B!����xI6�+B��6���E�O����X^��KL��=::?���(����՟?��CB)On޾���|BTt=}*c�����;g�e#[�����5��
k��W��{Zȶ ���=D�
�[�05�Y�v?^OT9f|�$�,�KTb�������I�1���+H4|��g����o�um��!�ǵ=ۮ-l��	��.?����m���x{���$N�>��1;;B!偸Ǻv�>��N�!��[>b�ڮ��^�O�(Z�,��$\Μ9����E�$��ߩe������ͱy.Qe��&�Z��0�GB!�B���ë���5Jw�����nuz/h��y�s\j~����իغu+���A�gzj
c##���K ����2���������CB)/Ξ=���aeu����uAQ!j��s�Qj�:}[k�~D����c򹟚������d�uC](p��T�SC6�|38La{ʲ���̑A�~�q�.,�T.I�k׮�����|�M��������H�mO�V�k��+X,��!�S.J �W�w�������Ep�R&���_��?��T���ȧh����+c}	�5c�
�彗D�n�k:?��[�n�����_�eշ�vջ�:s%���}=Q���%������@!�B!NkÅfa�53�rpW�-EtS��^�e}|d�V�1�������?�D��_S�N�t�t���k�Կ	SSS �Rl߾����	JD͓��D�[o��6�3��8��c9J��;�LW9����ִi��Ԯ�B�{�<3p�:���N�LA����vd��m�~0-��/�rJZ勿|�2�mۆ�Q�����;hinɶ���n\O�f��P=�4����u��T�����K ��+����1��w����� �oΜ=����-,J���;b�R��5�AE�J��d}�_�_
a�5��y��@�A$����	��V��eX6KBʺG��Jم�9�v���t�Lb7���Ƶ^�TC!�Bq3W���3c�՟�"w�)�Ic,/�"Tҷ0Ƣ�=:z�07;BT�UC��[x�w�H$@!$��������x��@��ٙ���;�16�r�r�N��>����^3L�h�U��\�а���wo٦�ֵ�yo��!34�ĵ=�XY^�[w:���⬮r)�\�D�awc��r�|��5i�/^�Lݾ}��@��O>�[o���\�e}躶G��36����{��^�����M8w����!�ē={����]�~��-��N\�����Jsm�B�h9y�$����������n����}�� _UM'I%�?�$!�B!DΓ�j�:�����=���Rr��1���Q.B�B�oܸ���v��̀���o���Sl�ĕψq�|��x�W����B!��7������� �<��n)��ҥK�5���߷e|l{ _[W}N���-�6�8�ч�0�6#�8���n�۝��P�9���n��#I�8��ݹ�5i%�U�G���"����Y鸶[�T�sW�D�n1,����u����	�}��NNM���C�@?!�ċ��f�:{_��ƱGo2S.��R���`]a��X��y���KÊ/l�Ŏ���OOr	�(�կ~e{���x�ee�?N��a��%��ֺi様�'�B!���H���F$��������3�R�k\����]���j���؈�7o�?��?@���Y'N�=BT,,.���'8��ݽB!���ի���/XZ抾D���
z�w�D�����$�q���S6�i�wp�isU�>k�ܓI���a��w?P��ˍhO%��\nP5�C+A��潅�^D��7^,7�s�N��΂DC���5]]UE�vG�b�J ���b��n������B��m|��o�νo{��;��G�.?@P��f�����їD�n�_퓇2����oF�V��>v�O��;Q��-Έ)G{�M�0,ն��ۄB!�BPײ���y��mm��J�)˖�TW�W�U���v�a�%���_@�aue��$/C�xi�6�ۿ�== �/<���E��/�?~�D���F����h�홱��9�E�����؆u�mY�ُ1�7�����q8��MU�Y:Eq���r�Z"ws�92����{$��
~��,$!��ӟ�����|�G��\�%vmw��+˵]���}���������?������B)b9���!�v/�!��#���E��+�8ߗ�^Va�G���,��@���ٳسg�g��tfȿ̠�s�}����h�zgj�zc��B!��f,ьF��[���m������].�Uó^hi+c�B�V�߾}�6mJ�I�h[���He�������701>���9B����x��~|��� �1��|�$:�n݊˗/��Ԫ������0Z�����f
ߝ�*���c�?�Ը��*�>�G�����ݛ�8;c������w!>���vdȄٓqKZ+��7ޠ�=b>��c9z4�8�����rm�����@p�:f�?�z9>=�S~�� �-Ǐ���,��MW%����!��*V) n�%"�9qK+��{ih�����<|�	j#��V�;�s��i+t������p�#;�=<C� �7�f����{�^�VK��ƽ�ݍ݉�vbw^̾x���b&B3!͓v�Q�>�eZ�k�&	z$  A�{W�ŭBUefݬʬ����/�jԭy��Js���s�)�d�HK*U�x��!�B!�D�^�6e�H�z㏀k܈�5δ)�R�m-&�1�'7���,�1���C��>����悐H���%�ُ��}�w�$��(iiiرk'N^���D������8ǁ|���4�2o�.@U?����^1���|,�K�W�Ⱥ�Y(pw����/n{ج����e�C_|�"wu�*�Ɛ���'�P=��6`Μ9����0�xX^�ڗ/1g�ܘ��]�M����Ǉk��\�Ip�v-=�=�^X�7�x��� ���EE(�5%e�Z���H��vӱFk���<c�v3�{Y��v#���x���9���}{��i!a�FLL����Jj���dc�IS����I�B!��ȴ�� w^��8����l�K5�W����A���a�%&���g �QQ��wa�u��U�ܽ�_ !�gٷ?.^/�#b�G�C��v�ޭ���6'�#!����7����}?+j���h+�)��)��z��Y(pw�Gi�E�>�c���Y� T��Ǥ��$�$I*' j�|̉X0Q��g��@����;����o���=�M"n���Ʀx�˖B�k{<b����b�Z[�|�
446�it#��X&M���;w�ҵb��>bM�nFDnu�V"��v�ۍ�	�vQp"αc�_��l��xc��n���i�*�2���v�����m$o��aB!�BH4��S���6\�O�5'rW�cy�5ƊD<��֭[1c�<}�����Ԍ���@H$:��PS_�U�V���� ��k׭E��j���h4�֡���9/^�իW;*\7�����:��"R�P=����V}����fL1��y�fL�}yUKF�B�*u�* tO��v�!�U	�U�b����`6~׮]����o*)F�˝��p��1LKV%µ]���wm�k�ŵ=<ބ�τ Oߵ=vQ���*�ݘ�]���<t������!��� �<|�.߼&�>'�>�8a�nl�&nE۩)��4,��v3�CCC���q�<+����is2>�9�f�T�d��2�Q��1����HB!�B�1��fb��|u(�)�b�(�+���C%F���˒��=�>���}����q���rl߷�D���gشn=�͛�/^�BHbBٔ�t<�k01�x�#�r�С�չ��x;]���5�Mj =J��q�F7X?�"j�{T�{�:�T��Xf���!��d����^����Ny���U�N�}j���B'�ڑ�mn�>�+V���r�D�����W���9��=�M"n���#��wm?�!��C�jU�gY�� 1�����<~��N�'���O<G!�~<���]w���X����ܛ���8����}V?��}�arrr|�&�p�j���w�M�,�h�v�k��e���-�`*��S�N!�B1FI� �e�M����\�C�?��?+�*7��K;̚�Xb����T�ėښ�l���) $7�����{|��mmm �����0w�\�^B���܂���d���2�j�ڹܡv���Z&V�q�WeN�4˒k|÷��l<l�s�&_
��v #����-�*JVE�K�G��{Ff�8���}�h>�}�(pw������������E�Y�|_����JodZ'�P�=��F�tc-�l�[v�5�i׼�ux띷}"w&�	!�^v�ٍG5Ot�>"�[�{��3u�Y�����0���KkS�ڱA{Ճ
gٿ���k��?>���KR��c��̩ ��J!�B1�Ǜ�I����d�f8������?Gͱ��3Ɗ���֬Y�%K�����9*�`��� ��._ġ=������!�{�:�G�ӟq����γz�j,_��Q!��}��Ǫ����FK�~�K'��D�pR�,x)n�
��N��姨�۵bwY�<��A��H�j<�1���ѣG��}��\��)����K8z��qm7gBЦ��.�í���b����q�C�h�hÑ#G��矃B�=�]���him�%r�]ۭNr���| �Y�c����(���z������ ��\߆�v��]�n[Ǿ�`eG�� !�B!��ù����3��&�1�7���R�n�^D9���1�[�F������a�?~��׬BNn.��8�]������>�]	!��CZZ��ۋ�Ιz�"���N�*=�Y�1�'��v�e�ƾ�q���h�X���$����I`�06(pw����lޔi��lS�u���4#�d�li���Zwc����&��Ν�6�ڵk ����w�>Lʞ�j��k�,����7k�=6bl�����"� ;v��M� �_���
&M�Cy��`������=ǲ0�L���=��d,�X��	�c�?W�=q�iӦaǎI�l�z�����1���&�F�I�op�m��={R6*�� !�B!�%�#؜y�(�&���ci�o�d�e4> p���7�d$�:����A����p�z1:��'O�BH��I�:{��e�ST�>���IOO��s�U�n&^YT��֬�l�^�m3j����,��vǘ�B���t��#u�%���jS��91Dsc���?��b9�ÇS��0����z�
�8�{�k�,.~��&D�m��H����v�z7�'tlooÌiӱr�J����BH|�>}:�/^�;�K|�������o�F��ٯ7�,K�v˓��$J����sb �r��1ddd_�A�K��c�*6�I*�x���fܭ��Ҹ0�e3
f�[Oq;!�B!�m}#ȟY���Ni�P6&��C�X�E��z�@���y�E���F�\�t)V�^��w�8Ǔ�GX�j%2��@�zzzp���m߆�+� �_�a坲���
���x��	��l޼�gώ����p�5Cm�r�^�6�6b�fl��o��"��Q�+�;LIS
֤Jfo踸�;a��B;1xn n�|N2�1Ĳ!p���'tR��(�??��۷#''�� ���!�iwm�d"�x�}����D�eA�M�{�n�6�*���	K_]�;kjj@!��yyشu.߸�{����?҂0�L���=����cEK��g �"��9�����h�7��D%�Bz��Q-�P�^�:$
Q����0���lp�AB!�BH,��OW���:bw�R顱����^�Okw��.#-��X%%%��$�exh���ƺ5 �(ͭ���?k׭��;w@!$>lظO^֠�����q�#����=�z�pݙZ�dRw�=�,�dq=c,��#�!v"�G��B����wy�}�d���9�EZrP{�Dr����KB$֍��DVnn.8�O>��9���q�����.����n�/c���gM�k�� ^��a���>y
mmm ����8p� .]/��`��}���/�"�޳L	����k�o@Ow7���Y�+V��K����H���m�)$j(��*!�HH�r[����sa��aޭg��B!�[S�T��+?G�zC.��0gw��X^�9�w�cEBoǏ�w��]�#4q�G+���אEwb��Ϟb��7�l�2TUU�B�5�����A<}N�#b���A�|��Y


|�H��zN�e����za�M9��d���7깷��}yW}��.��=#��E�a'���=�8/uc�$���~'����᷿���c$����Sضc������V\��qtm7ؽ�X3�?KBAo��*V�����>CGG!��#--��A���Ȅ����X���k�õ��q�χ�.B�+V����	��h�����>��M��
�V|w�%�����~Λ:��B!�Bb��u���ahpP:�Э#*k���X��|�L$�R4�l�<y2��ۇO?��9����X�v51ý�R�ش��ݨ��!��ؘ�`>�f���;7A�Y�^��{���&M
�v���>���s���wc�B�����xQ��
�]��L�1�� u��;1h��nwc�s�7oƒ%KP]]��=��z�
����{�W��k�_-�nr�k�?Ԙ�ݺ�0��?�q: ;��ϟ���c��>�%�!�CL�<r�(n������$"Q�k�p3�^��Y�I/��L3�q̿|V��.��_���q��!G\ⱏX��$�cb�CȉA�Z�4I%�{��e	!�B!V�)�H�tըH.��0w�)�̓��^n���)xx�P�j�u��A
�]@��]�<I�.߸�};v�r6� �b�3f`��E�2z=%�,�}}h��q1�uC��bm�5>�0����y�D���K5��[�m8�������a,����aT�\B]�@����
f�!~��Ē��YN~��➥qq�cݵݪ�ݲ�\1#,�o���=�|�u��4'�/!r띷�O~���^B��o��'p�����5�&�>b|��X���@��p�/qQ|/,%I��Jt��?�?�T����f��B�v����&N� �B!�X��/EQ�H���jbn`,6�	�uV~��'�1֎;�`�<��9��|.YB�r��>���!����B�1�M��U�����AH,<,-�{�x�W�n�:�E���G<�5�Wcmх�����h�KV7�����އ@b�w���gLG_k��ҥG����$V����7'���}�{q��{1��ߧyG_�K]�#�=�?y�a�����u���c�x�M��w���� !�����>|w����G�n��#ք�fb훸eQp/uV�nf�/�>GG[;222@�C��B�n&�H�����S��L�J����x�"����=/� u/�� !�B!�%u�845͜)�v<3��F'�P��l�e6�ic���4_�����>��T=x�e+�#�.�$�_��;��z�Utvv�BHd�L�����Q�NbF��?��FF:%�Ns��	��-L�b_�YG��S�z�\?Ԏ���\]w����t��S�j^M\B��$LI*�L���.�7e���n��G<Y��s�b���x�"�����slݱ�Yِ���F]�ÿá��c��ܲ��&��8pm��3����A'��!΄#���GœG���R�Z����d'3A3"r�����'����`Μ9�����S�$��D���&vW����\F4c���"D��B!�B�!�F��)����lX�*Əh�����,3�R�b7�J�(�f�������~���.�Utq'1"��/._���{q��	3z!� ??��n��ۉ*J�3<L���dff�СCq���p�j��6��=l�x�`�P�f�j7P7̙:�&��«�K��rG
�ͻ1��F�n��T2�����#��D��}9r�w ��.\����7[��ь�{��%����>�X˂6;��E���_(��^���o��6~��o��&�����h��P�&�>�lTn&־�[�?~��f�����>�v�<!]�,��6�x6��2�����ɕ�k�����t�U����L'B!�B�u���=Ҡr��C"�%K�kW�JM5n�����i�������vK�,��͛Q\\�,B���k�"3+��E\��~yGĹ3g���B!j&M���w�ԅ/b�"��+�@�g׮]�={v�'��ݧR���Z[�Yo���=��ڃ��9`��:����0�`:zۛ�UV�Ė�j܍A��/N$����;�����A���>����|�D��܍ݨk{�
~l�[��$�wܵ]�5~�fD�C�x�X������o@!���;��--c-�����eYDn��e�����In���@�;�н��eӏ;f)�V�v�x�b3���%�ԛ7�jZ'���$wt�R��I*B!�BH|�Y7�]�)���?�OQ,�_c,_@�^	���=��N������V�_BbA\7??w�����@!�Ovv6:��ϟ�=?+�%�i>�Ę��ѣam��cmsbZ���u
ջs���5C��g1��vχx@�����E��^Z,��Eqc�o���ɛ��S^3�ѝ�H�X�����/~�؉��	!������$F���O~�W������>&O���P[G��e���g0'�3AA[ͳ�x�|������Y�������756���I���Ϫ=�����:;;���S8�p�ɲ��>G��]U�H0���I��Ku�p�;ݿpA����mN��g�ZWW���w���n��_<kh�;w.N�>���n���L%ikknAEY�$��5Ȉ�|hh�����}Í������*M���������6<�|d|��M�ZZ}c���\�k�}�aY9i�k�S�ց��B��-\�0b�[� ��>B9)�#c&Q5���DLR�%��\<���B!�B�E����NGog�����M��#c�~
c2��ݯ���?�3���@�%��>)'�Ă�}q�<�3�N�B�_����~����cuM2>�����G�A�gƌ>�d���ǘ�v�x�`�Pk���F7�R��s���@�3���.�F�0�MN�]�<Qnj9��DKq��B<����7�|?�яl�U�����8%v����I�����~�k(�2E�.���/���g~���@�x��x���A����Bܾ{�^��5]#�Bܾs�n��j�k�����.^����	v���:�����N�BS!v�9s&�����X�`�B��-Z�H�����m�ԩ����gw����&���ů����.�5�7o�#����aڴia�۝�����������U�����"��r��@OW�o2��ysUǤs��&Y�qq�㇕X�|Y�8�n�=ߚy~\Q�E˖�}�ZĽ�l����z��7�|=88'�'�o��_�ͅ{��-R|<���86��KT��+]�ck]a�d���]�WX  �B!�ďo>2=M�b������*V���b%&�[1�
_E�}�V��ǤI���[o�׿�5�D�E�NM�w�K����6�G.�~��Ήk�=]����Bz�3����v<��v�o�����C_�#�;�مA���|u;�͙�ǌ��D7g�`��N~vq��ߩ�8�D�fE���ɿ}�ϩ��g�E-�����}δOC��N��ă�0�r'?{�������@<�4�N�1���8u�{��T���T�eJ�kH
kn�g���rc,��WR7l����.��;�;u:��[�&�B'�|v��p/��Tcn)c'����b�,I(��b�m۶�ҥK �"�O~v�'r�㕈\�nx�b-��M�����-�M<D��_7&�[p��ߏ��|��������'>%���Ğ�{Q�܈��F$�>bM�n4־�H���f9v��#�T��J�N�c֬Yؽ{wB�Opy�"1h����OTI\%����1�x�����Z&�!�B!��v�5�q��fp�S;�[5�R�����D0�:q�>��c[�s�D��Dw��n�8@��\���'ǭ����ȟR0:�wȨ��ڰaE���G[Kf)�B���=-3�֯GZjjPl�H��)��D1�͙����3hr�͙�9՜9�(d��/_��ٲՇ��{q���O��H���.����/�c��E�'���-�H��Lu�z��gOd�BH��uճ�0��/�Vp�K����}��~�1V���s�=�w.T3T�Q��1�2c�%3��w�>���
�]F�'�<���'�70{D2�Ŀpc��%n�#ل���w
��A�����0s��O�H�����kT�gYDnB�������Po��E�v������x��i��W>� ���7�$�!$шg�����Z�Z�1V'3���X[�#���m����H�W�> q��+]��7�|T@خ}#4&6����0�N4׌ս9�@!�B!�σ��������A4Escu�ݱ��v��}�c-[�7nĵk�@�E|��K�cˮ �
���y����|q�#4Bq
1�c��=8y���Pz�$.5Hba�5��q�ڳ>��-��c������H�ʺ��u���i�9/(pw�j�ؙݍ!|�A���	-Q�h���<�"�1�p����}�۷s����"%�"�ϟ�G|���"������n��ܲ���=]�#�
��Gϟ��w��~�{��;!��W���#ǎ���J�����o��C�v�N��Tzx��Q71B�0?~ܶD�'\*7A��U�1��2�è�K����B!�:S� ���0�
M�U��KV��#�B�X��"�����
c,
��A͓gX��uL)�
B� ���;��{����/���B����cۮ8}񼭫Ӑ�CKc�^P[��F��mf�k[<�kfjC�P�ި�=d�%[���0��z��n�Q��=y`�0~P��2�G�7w:�:[�KHg�x�Dd'�4Y�I��<��#���}lB,"�U����@��֍�س-^�x���k<֨�]���U���vƙ��*�4k�%�?�����?2aE��g��G��~E9:���޷�>a�n�ν���ͪ�^'�i�z<��}�}x����I���͋�f���LK�GNRi7�n�J6F��3	����Ƽ=!�B!�D�f��2�jW8��]5~�*�6c�hE~c� ���1����x��СC��w����z�)�[������k���p`�\�r ����ԩS�e�6��������xp�v	�;5�]�v9^L�˻�
}�f�*ǵͱ�c��� n��O(pw!m��O��.�r����'�dN�D�:��U]D����h����\��%|�_�?��'��݌��M��M��]۽�8����nQ�nU�3� ��{����'x�����Ą!d\!���@ɃR�h�V�zIv�v�����Ǔk{�����3���n@�W�;�fv��ٽ_�{����х�z�*��^�|<e�A�Cj��}Q�N!�B�����/,B_wG�^u�g��MV�OM�P3��� l�ceff��Eݐ8O݋Z4��c��Y �*�y��8�{/n_����fB�x���k7����gm������5hnlqo��6��CR�d�Z96�dm��@�z��,���Z]7ND�����	��wr�ދ�Y��=�|�"x��$��41#t�_(�N��O�$�Ѿ�Ν�={��̙3 ����c�޻�UkV�^�um���ܲ��h_&�tm������̇�U8|�(Μ<���6BH�#�m+W�����>�{�#��!a�{��i������6���,\�;w�t<�����;�skfPjQڄ�j�\fp,6�2��Nè��핓�	!�B!�ѝ^ xZC�Bc,�8�;6�78�	:�k7��ϒz!����X?��}���)�y�<fZ�C�q}<}��n߉���h�X�2�����kW�&�/Ľ���� �@h�1V�k~n]��?F7Y�ea� K��sPgn�%�`��|>��m���������>�f���=����y��jڵ'�p�Ԟ�A�g0����,nLB�9^��:{�3��o~�+�����sF�&D�m6	�-����(t�*�7k������I5>��KW���KBH������������g�DVV��ݾ�����5'��X����:+X����[|&v!---���.�ݯ�$KBA?I��믄a�A�ds�2�YY�(m���B!�b/��S�.-4>���YR]1�״)�F�>���-Z�l~��y��hk���O�p�����>�{z�C��ւB���3�\x��2�'�+����<�9s�D��K�ﾌ�{��G0�VL�����by|����zz���ݥ��NA��Ew�G��tI�~1��+^+/����$�ō�-I(3���%K�����yZ�[p���ڳG�M"r��6���{\���&�k��}���'��q�fL��B��RBH�1}�tlܲ�����s�(X�	��X;~�X;D�n�|K6е�-��������`u�������n<Q%GZf0l�-sb�oƔY�42QE!�B�������K5>��_���Һ�̥��XƏ���ޢ��Eܿ]�� =��?�_��m7#7/U�U ��de��#� G�k��-!�bhp���jS�6���g[<���pիmP��c���jc,o�q��n�?�mOG@�G{.�����A�l��B����8�\VA��6Y%�I��%�G_a��I(#m����{����m��᷿������h5#"7kB�'�n�#X��+ݣU�[��b�~O�?��EQ0� �/s3!$yX�t)�,[��7�����9f]���l�-�,
�a����"n�������(,,�N��]����*�P��u�J_�.KRyu��a��&����Q�)Vʠ�;!�B!�~z2��v����Fc,+�ݽ{�����ӧ ���ׇʲx}�*O�o^����M[6�Ƶ� ��dc�ƍ���͒; $ޔ��bp` ����زe���D�C�S�G^�Y� +�S�Q����q;�q�w��50�ܹ3��������_^=5���C���\\���$2	e�~�ڄ;�~�����8O_?N�:�w�v���0'h3#�7�=��{]�-�e�g�����ô�"���[�㧟rb!���Y�ٹ9�~�V�ͨ���}Ą`�L�����{���!����_��a{ .1�.��DL�5ow�]��:	j�T��������^�8Z7IHP)��9��(��r8!�B!��ō:`c�W�����>''�]���4�fcb\���|�T��c�+K1)7�ē҇�X89�M�fHI�s˶;PS�5�/AH����FuE%�{��W�6�X��5?{D�!�,���ߩ=\'nY�&l���7j= �w�8��O����_|?��N�HM�8����)^���T��3����D�{����<ߒ�?��A���3g�}�v̘1C�nYDnP�����x_�tm�EDn���ٵ]Fsk�s����C���;�B�Ȗ�[�34���I��#���'�eJp/�G��6q��� ���;v`Ŋ�LDّ�
806u�1�иX�̠�Z+
�h&������ENCB!�B���;�ɋ����]��.��V~��yB�T�X�7FSN2�1����w���Cttt�8���������[AH�yV��=�8v�8N�<Ś!!��ddd`߁��q����A�ܿu�7V �@��,V~o�W�⵲V��������(3���L�u'�KVV�+���j�ws�փ����ur����OXɜ��5#��&��PF�I�v���~�A�K�����_����#�fYDnY�����{]ۥ�1�#��u����C���W?���)��\Kq�Q���C�z�-�-�6{�#��D�v�G����:\���.��� �;����1����!a{�g���e���#��x����=c�8>$�B!�$�o2=-Q��'�j�򕮴�v��Ke�%q��7Oc���|������A����'X��2N+!񦥵�/���c8w�,zzz@!n#77����]����A�4����������#''��Q"�����ۯL�ѸeE�!���F��ZS��Yu��~h2X7�
�]����Sg���>b�J���'���a�����8�zÖ�H�$�D����o�>�:u
�<,����X���w����ƃk{X�)�[���iFh�?�wE>��	���@!N������.-AOo������{�(����#Bw�����OU����K�b���I��2ۗ@��
��D��I߽=4��q�,c+&���
����I*B!�BHb�V;��y)a�LE3����+]	S�ڡ�M�E��<����������A�G�ݹv��1=�#����/N�о}�}�Y3$����ӧc͆u8u��y�;ㄒ��A�Cvv�ou)N��}Lr$ZW��C��[��Ħ�𦥥�z-�vA���y�7	Eڂ�$Aeĝ����I��Q&q��dIBY�_�N�>�Pa�̯~�,��ː���h5!"�,h3ڗ5�^,]ۍ��*���
l߹�e��� !�8�̙3�q�f߼���g?����k�E��)���XcǤ;�\�ܽ~�Ͻ.C�*%���̉(#}�Ƨ�ve�JyA���uAol�ua��2�G!�B!��3�E�ԙ�io
��[�9��;��"#�/^�={���ٳ �����% ����乳صe;�rs���cB�ӈg������� �N�+*����:�9s�8^�K���\���\+��:4.�7�RQ+4�J��I��0�b���;���%-�k����w��ܣ%�����;Q��x�NBE�j_[�l��5kp��]w��ڊ���Б#0-"�$n�&X��ںQD�V����x�={���,��чC����hV�\��sg��kWl��X��3u\��Y^M��'��cǋ��i�c476�����;v̱���ɱ`ZJ-l�:Q��k��v���ݣ3�\=��nc�h�t�!�B!�$���y���'=]];4,r���2�:�{���z!��Bm���.����p>222@��k�ū����X7u
�ܢ�-!�96oٌ�����b'��(�{�=����h�dqf�kw�����M!n�]��v�&�����b{֗3�+��w��=�2
f���eXaݣsb	W?�C]��#:1(^+/�����b䶄S�m������?���QTT�j7%��E����`݌ͭ"r{�����g��x����yy��W?���)���@!v#��v�ٍ��N�,�c�c�>���wjJDn��-3�e��!Bw��]044��;% ������ɓ���$t�ǅAo�_^0R�J������T��&Q�?u�R�N!�Bq�/�p�0#�=NwL��*ꆱc�j���Ac�H$��=Rێ;|�eee �  �Z�i=��;��0w�<|��~��BH����ۇ��>!v#&��!q6l��u�\&>�_���S�5\�e�ʺ�n�Pn�5�̬,ܩD`lL��I@EG&�y�GO��,c�Ɛ�
$�:��׏�,3�&{�6����uuu �@<D}�?�����l�~�,ڌ�]��n&�k���ѵ��n�а��=��8�֛�|�2�jkA!v�������Ni	�::u���V��-��V���#�c�*�wZ�]P^r}����&D�Z�e�I��D�ڳ9 nW)��^mJ#b�}DW"KT��v�N��	!�B!N14dO����z���Rǹ�t��HĦ�b6Ƃ�f�+�E�ь��x�wwQ]Q�E˖�`�b'/�j��юc'��ʥ�hmm!���ԩS�e�6\�z��|$!����Y�w���������g��иT�0 n����uEO��u`��B��]8�F����$��q���axpP:$�r��U�%!qf�z�'��Z�$��"�Hm����dտ�˿����wKP��._.0(h���n&֭"r�5a�u�'�mW\oVWa�����b&�ܾB�7���Ǫ��q��˄�V�#�'~Y�'�e0N/v����l�@��Jwq��!��&�M&�H�{ ���:7�cTqr14N��kU�uΞ��B!��7�=ãc�C�X�՟哂�b��i�u��q|�{�CSS�;��;Wob�у �nz{{�ǳ��e�F�44���
�b+V��܅�q��Y��Idb �gw�����e,X� ���O��_|�
d����B��x��[h��0*��G��+�	�I�H�tx����$Kss����. ���6�̠�cPaJ�'���}��_��������|�����_��A,ڌ��ڮ�}�D�H������>m9�3�O�����o؀Iy9�t�N�U�E���8�f�\ۍ��t6��nHݾz��3�!�_�����dqF�b�?�m�ra���"'�d	�@�*�p��!�B!�8˝�A�3k����-����X�6co�����'���+�{hnlD͓g��x!�q=�z�V��;v�ĕ˗]��%��ĳ��m���݁3σ�D���- ���?DzzH��&�{��d�uC�M-n�b�*�Fwo�7�
bi&�O��Ei��vC�{�PҒ��F<a'ˈ���������� �r�^��()1h&RR�/b��VPP�w�y?��A�CkK+Ξ9�c'N�tm�V�C���#p��ܪP�L_��S/��Ѹ��fL���WG ���?����+b �w�>�l�CՃ��s"�k���_�E䉼g�ӋuZ��b���Ghn�ۘ�عs'V�\�x�I�����jq{a����D�J9�V%���8\0z� �B!�'�򔼙�4ר풉�ac��B~d�h�X�#S�<���~򓟰>�2Jn�¬�����	B���
L/���o����g���B���L'j�7��AKk+I�}���.��(**��o��*��5G�bӠ�*k�Z��Y�v�)�:�Rڔ� �C�{��m����S��nԉA~�z��jf�A�����῀(�S\�p����׾�5�����e���$V�]��s愽g\�f\<h�>�"rsBI#���M�k�n1�3��ׇ�G8t�0J��Gee%!�,�f���-�p��m�Ȟ/��Gd����b�pm�߅��J�v?(�S�.ĸ㣏>
k��9�	;]��*�vu�*z�J�ܮ�T�������B!�B����t,Q
�u�a���f��]%nW���| ֕�RR�/b��6e����������e�)��-�@H��Xg����޹y��� ��X�3w.V�zg/]��0s�$��ɂC�� �BL�����vS������B�H�uB���R�Ľ}dă��i�={@��$�=m*�=m:'Md���M���*��ܕG漰�,V��={6�?����7 �A|������_����k3'h�C��V����wZh��߽�Ǐ0o�"��lN~���zL!FX�a��B�ɻV�#&��c���g���uZ��a{���o�D��]�Y�[�nE�8KDYuaP�ݵB�p7�do�I+ɘ;�p6�A!�B!��Q�kLEO��K�V(_�9��]��]�f�ө�j�,7�#�Y!0A�W����\Ɠ�GX�x�fL!�b`p 'ϟ��u�`�ܼy�b�l�i�f�>O��x�$���:�<y�.rss����#%e|�ڍcƠ���b�L��;�G2�ҚQ�O��gO�K�'�/F�'/E�̠�Q.������BȍAv���Ag�1*�3�L.9��.����1̙����ӧ�y�:�l��Z�v+�v��:�	����õ�(VcM�������|_^����zB��y�سw/TW���$ª�ܠ0�L��ޖ��E���+W�G����5O���1�Њ�$c�����̱�0�O��{,5(OT��#{�g��!�B!�;�)��$]�Z�W]3��*q�3o�%�xʜ�̗,��xc=z���oA܃���}��8꫃�H�߹���g���c��aOO!$y��]�UZ��f:���#�w�qr�y�w0mڴ����b� ˨�=��9�{u�J��l�g��VL���IDϠ�
g���^:3DZ�OKsn�w��KR��D�(��jwu�j<��#�-[����ǩS�@��'��5��X���U�Dqm׏�*�4�+y�D�N����(�|��֣��/^!�hY�|9�,{Wnݐ��`�>�3���NM��w����>�$�y��� ��W^�5ܓ8���=.���.pa�*I��P��_��/(n'�B!����^��AX�=�)�gtKS��,Ky��*1�(�!c,_%1�'�1֧�~Jc,���֎��X��� $�445����m�&�44��� �=����-�]7�Z<q��J����.233�կ~U����2��ޮ�!d��F�*Ǹ���X�U�[jj
�׺��?^��=�x�3	3��qcО�"i����|/��.]zP�:D
��qɐp�������Ӯ,Md��������ڨ��+m5g.6a��^㟕���c�}�׾@���x�+��_�]BFIOO��{��ՁKׯJ"��G
���&�>bQp�����(/����Nw!��(����j�ō϶`jʰ�]-r�sb��̠*Q�k�d	G�B!�B����"w�,��5�L�t��v�1���?&x_+� +P;L�G`�4Ǣ1���bϞ=8{�,��9�� /?�$q���W�,ŁCq��yB�Qغmj�p��y����,�d,7"V�Z�p!R\^���z!��+��������^2��G+L�m ���u�DA�{�q�n������`����L��=�DMU�R	&���v��]y���q��h0�%����_�[�nEqq1���u�&�oڈ�sd�.Xw��܍�{��;-44��>����щήnlݱ7�]�s!�Y�fa�捸y�.z��4�Z��X�����>bQp/u�}��*&�܉�V�8qnOR%ąA!n&�"�۵n��=����6Q%^�}\�!�B!������(R
�5�X�L�B����J�fGc,sm}����W�&"�\�s�v�B���q5j�j���A�=u-�� ��ٳgc�����������ϯ��������HKKsĽ�i�{�`�P�!�]=���y=��a+>k�uO���DA�{24i<��ԅw:��6z�S��cnju�*��+�,�"%%�NVڄ��իW��r!?��O�������3�bM�l&�����E�����~ݚ�эn��L���g/j�_P��[���3!d� ���m�oz*.^�M��*"�����5�v�2x z�f7�G܂�7ݸ|�I*�"�����׉H 9���B{�
���#v�NbJ7Y5�^^��V�\!�B!���[�CxgV���B�B��\4�{�A�ܹ��X��6l؀͛7�ڵk �O=ƢW������é�_`ڴ"̜1uuu��#B�C<7�۰i�8y����y��-M�|�F�*Q+W�tA-Ͼ6-�1�N�*Ff�5���>�[[7�5���srsq�nJ�,�
ܓ�[�X�ꑞDF��*���RS� xe	+�ɪNb��$g�hۮ]��v�Zܹs�]tuv����~�#����(��(׏�*�4g&VGi�H�v�ۧ��]�mj���D�Ç(/+!d�3{�lظ%�eh��м�ዛ��`�����@�^_�"�:)nO���������V�1m�4�����9 ��;����1�9��O ,Y�NP��T�x��)y�J5�k���<��!�B!č�:�7w<-�U�QE2����M��KE�ʣ�8�B�1���ד"G4�(�y3��¤�1!���I5�L���Ǐ�ڕb����2q(**¦�[p��6ZX�!.���ew1��Di�dq�-d�eDܮ�#�̟euC��6l��6�L�z���$��˃������=l�H�tr��	���0�wJHuLX�/.�3��III��S�m��o~�����W�`���X��rU�U��u�]�qfbM���n<6>!�o���
3f��{�_��S��=:X ��?����];����W�H"��G
���&�>bQp/�ݕ����щ���d�V����#///�:Q�[���GPЮ�h�*܅!���ޘY���2��p�Xy�.�B!��r�)+��|�l<$��׮�po7c���Lc�`�pX\�f�޽�.�q���ؿ�8M{{�ϵy�u�N���K���&!����͛����;����D&���cxh�}�U�7n��"���m�q%$��fo�ڡ|�T7���s�(K�jo6���$qP���4x� ��<z����KT�%���w�M<X��*g���X�7��T��$g�h�޽{�~�z�ɪ��U����ɾ����?���dggc����&��ScF�,i5(�.�}�}�b�pmׂ��^C}�[/������4CǪG�BC�g�}��8�&7����{���1=�y�������A������>4����N���=d:��D�ۋ��w�'?�ܹs�_0eU���^w,^[}oD|�~�G��zrL�"�'3��x|�|˂{���H��Y�C����^�v1���;y�{��\sF���嫾���YL�Ϸ����|�AR���+���x�0xF�v�dU`l�5e6<��B!�B�͋�al]8}�ac�Hc�HYF����BE�04�U&�1����K<��,!N#�7��F����� ���������B>v�n�D[G;q��h��qb\�o}+�M7�ڼ�-$nW*��Q��d�MS/��#�b��?�O���'�'
ܓ���L������4�D���:2DXrP�.�I#P��ĻM�ɪo|�����D��p��X�����I����_��~��_a՚5h[⩽�c�]�BCsar�_cC#���W4Y���s>�&�(�_}�&�F���C_���Ի5�_3����f<,`h���f*�;�|b_%��1);3f�D��G�������a���)�K�S�&�����	Ŀ�D�ۋ�wuu9ҿ�]|�E��e}?~�i3fh"L\Ǥ��~����������1ԻQ��{fwW7�^�F�ܙ��V��������z75�J�w���A��I�^q��_ i�o@��uю簀��)��8��dF��G�½=???�z<��cuaк�k���y�0q���0�f�]K!�B!�5e
2=��q͈'�_Q�
�+��cj��zZ@�~�n��ٶo�>������a�W��\��_[�I$⻘�����Cff&2�2�������K̩��յ65;ҷ0g���v�'?������ ��.��I�c,�� s��CYi��n�f�:V3w'����)����S�]|n'��-��N���N|ޙ�f���?�����z�"����;��u�H������<������N��N>ߊgz����/�v7mڄ����ihk���HY���u@U=�#��j��U�Eݰ~� �&
ܓ�!�Sfb��VZ��s�S%�Kj��nR�;��ɇ�9�M��G��x��/]���݋ڿ����i��x��C'It��e�{`?fΜ�{�p�"X6�b����q�f�XSn���vE��7o��˲k{�����X�h!�Ƅ[�:��;8���nX5N�l-�����X��5�~�5dێ���_8w>�I+��y���)D�ĩ�����z�ԩ����gw����&��� 77ב���W��/]��[70���",ze�"��}D��:q�l���T��
潦�C�8q���xa�����X�u\$j��;0s����K�DQh΂�p
���E��uut���b�@�ĳ����IN ��k�X"�/**»�;!D��mr�2{h���'����n�:��'NC�S&�!�B!���쟜�.�덁d��ʓ���ͱ�c!4nK�1�Q�0����QRRb���b'p�o'��K�V�j�:ߪ���af!�"55ͱ���=-}b~v���v���E}����i�V4���EM�-����+8�����E.۩��^g���2�q�ϙ;��ǵ���ى�ӊ��{���D6��n�\�T�n��G�ו�ܷ��W8��}������ʱUJJ2��bkS�P��Ɵ��a�X^hM�e��X�U���6=�^�n��'1�Z��J���*wo�IpcP^ �\��v�z�.�nqO�c����g�g>7�Xl�^~��?�G��3_b������L��Gp5֦�jE<hW�����YEL��'���ǻￇ[7n�ٳg �����BlݶO^<Å�˒�����ucm���\�����	���ĳ����:}�


��'B�J�_m�%#�0����ܽ=����PlM��x�B!�B���a`R�l���E�J�4�X�X��5�Dc�KoGmr���X�r%�޽k�����@��8�w@ ����
��.Ƥ�I���C�CF-�Uu�8�@_?������t��<�^�U�cŲ�غu+.^�w�q�b=y�d8������0fMN��g�Y����_��,V0u��9�{����[P�Ԉ��!=+٣my��������t�ã�����	�����ֽ�<��F}����V�x�v�=_�����m`B����s��͛�����o�&l��K5cY=c��cfM1�h.�[�aBC�{S�:�����6sDof�Ȉ��.�!U�Ơ��f����2��҃���-vɪ5k�JV����щ+/a���v���Ċ�-
%%����֦3�N����	֍��r�]�](�|�ů��UkV�����܄�!�;v�@Jz.߼��9o�>bP�mUDnq2�~l������du�n���R�6���1Q���ߟ���^Ŧ@������ubso�_�L������B!�B��Ҏl,��)�cV~3��q��1��6����׾�sqO֜�x�v�u�߲	���Ux��)��ځ��V����B܍xذqr��q��u�ĵ�D����n�q/v���k?���ǔjc�`;�S#��)�>c,Ot��h5Ļ͙�GAw'��=�iB!�=m�Y##U�qii~��r��W�Ƞ��KP�(]��	�ɽ�*;X"(���r/�X�t1.^�{m\�,�]ۍ�o攰Ghh��5���j�}�����a���ϝ� �� ���׮��ٳp����$Q�Ms���u3���gY����d}�kkiEEi9�{㇩S�_O�v%�a�D��P�,I%OV�h�T�IޢM6N��܇�U8�.�B!�����i����KU7�3�
��\��c�Tc��v��A���?���L܇��<yT����A����_bƴ�8r�*<���O@q.����v�=4��p����z��U�O\�ƍ�}��q)j�ަ6����m�0�s�Dm�f���N
��O.,'�;�I��a��)]R]�D��=#�H�%�RG�Ґ�ٍ!,qHP��B�<�@'9�U�L`�d���d��9��[�S�H�u��<��{3��pm7J"ŋ���b���E\k+?BvV�|�-�|�ׯ]!�9DrJ�ۅsJ��:QV�#�����w1.X7k��j|B�D�{��q��˾{
q'B���$q�)����R��Lܮ��
�޵������� ^2VV���vK��@!�BIFZS
��i������\�}uDci��������!i�K����<y��o�!n���	��;�W_Y��Ǐ�Zq1���@q���l޺/�kq��9�v�)VSC#�;c�?��?��V,��D[�f��B��@c����f�W}����"9�k��aTƺ�SP���� ��ga��f�J�
ڥ��90|'pj��؄�])lW%�?�x�2'�V}�))�#v��wĤ�o~�����{w280�_����O���(n�n��Qpo�7������X{>��(���e�1etp��{����[���!$q��Ԧ-���َW/���"ߟ]���$�>b���b�xI&Jn�Awg�{E�)�I�ͽ=� ��ݱ=��gD#^� ��}t+(��gta �B!�$)�^xpdj�aS��C�HZ��+m�}/���$v?t�~򓟠��ĝ<,}����a��f*U���jlX���Y�Z\L^B"337m}�J���i4D����6��Ь��lذ۶m����6�b��$j �K^?Ԏc�v�J�Q��cY��8��uC'��}p�1�R�'�T�|!l�.3>���M[nP����]x���0^I�8MV	w�d�͛7A�I僇�z��vlGB]�-�!�7�k�^�9���X[��h��@���ڪ�X�f.^���.�	�������� -7���v�;���nE�nQ�oJp/s�}$�h����*�2c�|��I�|�2�`{�}E�JW��˪6�z��h�v�6��b���B!���dpH�2-/#�ڕ㣴�13��1V�+�1�J�.�zi�%����o������K�����ߋ7#��7��ANNv�ۋ��6ܺu+��ل$��j�*M���wn����$����bN�p1�����Ͱ�TW4ڦ���	M�0�qU�֯*��ca#���0�
�c�	�A(p�vc����l3��.��������P@W�.���$�HII�dU,�/~K�p0�n~��O�ʲW0}��`�;D�	�K�Z��vut�H�k{��Ok����{�CO._�ā3!q&==��؞_0%奾s���ĺ�[8&��7q��}��n��$��y�*�������k7$��a��L܎��֍Aw���pQ{$�B�{�Yٸ�bJ�!�B!�$��2�W1މ0�W�b�f�Km�%��+���X����5�@H2��ۋ/.]��Y�q��Q��/�
Є���ŋ���[v����d����hkq/;w����S�f �NUU/���V}6�ޮ��5	y��9(p'�����M>A�'w�̔��7-$r�:1h��&�$ɪP�&$�NII�dU��۷o�m�/_q'bɶ������w�Y��.�[J���`��X78���%�:�o,��1i��E����:^�
��{p?<�����E
�	���<�n�:L�9����QE���H��b(6A�,��6��G�!n���=��,\����+�O����\����bw��zS/3�	�q=х���[�y�4��� !�B!d��݃M�����ݔ1�����Jc,=���X���c�X���h��r��}֜�(�>�$��u�mū�qh��(�w��� �ď���c�����EN]��$�u�x��Ľ��poW2Q��k������aX�F�nt���E3��1��NC��8���a�5+�C��ɪ���tq���a"��;C��]�'�+�N~qJI��*�HV]�z���&���'��޻a�%��\*��Kpo����=�v�;c-�<�`��ء�!<z���w� ��|B���~B�#�߫׬���p�A*�?�[� �X���G�������H�RU�u/^��q��������lU���D�%>a�Ulc��["�ܮ��
X��#rU��p��]8:�hːs�F!�BI~�S��i���@Q�c�4��=c,��n�cź�-[�����r��K8��qdff��d�Ae�o{u�+8�~J��E�K�	���ٳ�z�4�4���s $�>߸\<�j��C�a�ڵIch����Q����]o�g#��hbv�6<:��(=�ag��}��=a=���iyfj���+_�A/9�"��.�ިX%�!Y%n>��S�@�˗�/`٫˰b�J�k���5��5Ｘ�a�-V�W#�|��B�~� �zzp��e_;!D߽z�:,X���Kq񪿸�k���ݢ^�����c��@?����K��ĉ��۹�p�v٦��$���1���fUy�3QGB!�B�8��fǦeE_�Yf����3��h�5����ŭ�kضgIF*���q5^u9�X��ܺ���&B�3s�L�Z�Mm�>a�x�#��W}v?>c,%�ahe�-D�KV3��N�Y�ꘞ1�Q�vaTv�Vh��k]�=P�>��Z��^��*�I�����'�ҍA�Ȑ���C���_��z�>Q��dIV��_�%Ο?���A�����	���?(�2%�M�D�Ƅ��q�5k⳺�m׺(U/���E�,nPݟT��N��&:;;�克 ����o��������.����^�b��ڮmM�k���v�`7���d@�"��y�s�&�����}ɪ ��۹��m^�B&`�sc����핊�#�6¶����@>��@!�B/� ��gc��ቿҚ!��h�5y��O���x�R����OY�C�WV`Պױn�zܾy��� �������Qn�g��Sd��M�Ҿ��eY�,;�c���q��/���؎�؝8��L���d��93���{���Ξt:�N:��vbY��K�}-IU*�JU��J��\.?�  � ����"���G�x����� 9���b�����D��+ݽ��<���X�z�Gk�ۥEvn�3�Ҋ�C)��)�v�g3�/D��� �D�H5+�`��ۢ��OZ0��!_l�A�f����]7i%��e�{<q����*7�G���UW]%94��7��_�����/��u�"�D��BGG�e2�Bl>8�����N	�������8�4����*|�s����7TTT`l�O�⦴�7�xf46���Vl߳+���2���Vbszq��JG>�z���br�T�;r!�M�7�X��vBj��Z��tdJS0����b��jZ�х�B!�R`���z�~!?�����X� v�1Vas`Of5�c�D�s��1����u�a��p�i���@I��؈�7nD�`?>ڽ� kH���뽂�˗A�a^���O��y��g_l�6�R�墢�^o�g��a0h<�sZS�@@�W�{w���������Z,vE��R�����E^�	��)��JrcHra�
�%y��d�Sɣ\o�_�*�{�=�K�3g���͸��{���Jڋ�����|ݹ&�bm
��Mn]?��W���0F�Fq��	����?�2_)v�څ˼�!E��1���P?�ǚO���3��v�1���,��NM��4b2�(6_�#^���ε�Emm-H�"��P�B,���gv��y�Z��yq�F�v�k�z^�ae�E0M�*���'1��T�"WB!�B)$����]2��I���=G�X���2�J���X�.�!��o�=}F��!ċ�~����|���108�y���BG)f�,]�U��r�@?>ܹU:V)S�ٺ#�@��	�=��.]Z&WV>�o�fR�����M������jf�C���
������z����ۓU���=��'� &79i��&�Dǥ|��.�v׳h�"|�_��~�3����?���˖a�����������.�wYh�/�ҍ�y��m�%���k�E_��rF*6�Y-n����Çp��,)d����K�Q�O���q�rk��E��[����O�]���sy)��������[o�m�����Ė5�v�䔁�=�aKK���Q��!�B!����bv��Xq7w8c���gܮ
c������ ��`� 7��7�B
���{��sX�z�}�~\�Љcǎl��-��f��¢%Kp��6m���Rp�Q��i������eŽ]�|�'�C�,���0]?4Y;*�u��818-�� H~@�{�S2U���ɪ�"w1\�_$��;C7�&�c�)�zB)[�qbݲ[�pq����_�o�'��!�|�[�����9��`�����m׬�Ӛ�զ�^?0�.ȩ�/>��y���a�����ށ��tRP��J�>\��Z�;zXz*W��d�?�d��"r��#�ꯌ6��9�k���]m���H~#�^z�%Kb��K4e6/q���:�%�ԓ����h�*���LRi��E���aFz
�� �B!�7�xtQ=�GG�`��wFc�L�#c���?�oZ�O�q�L,^���mg�i��y���{11:�=�w3�L
�sڸq�ԧ=ul�B
��3-8�J�C/��SOa��ٞ2���z:vŔ��a�����ڡ���F5���8v���|��d{{ ͪ0��.�~�	_0&f�%	��4�*u�F�ae+Y�̈́�S�L�>]z�����	���?�^x�%�a�
�ӵݮ>�{��$`��}����̮K��a�|�{�MMM��� !^D���֭����y��؇#'�&�Y{��(�\�o�x��yā�#?�#�ā]{�����<���X�~��	�|po�'��H)� Q��o�>�-���a�RI��I��h���e�!�B!�����Fy�%�X�s;���G�~���������߽�PW_B
�ή.i����ͷ�
�M{�bdd���ո���ر}Z:۱��QR������} �Ϝ9s��/9ku�L>�^�1���C�	ݓ5�r�0&ne6곘.���a~A�{�ڹ�������ك����$�Bw��2tc�qdH�dU6���O�w��Ο?�ߴ�9�?��>>�3-�����vD�^wm���[�y���Mo�l�,�Rm���¾ҙ���'M�Խ�FEY9N�l�ɓ'A��5k�4AiyN�mAk�^�X��Xy���J-��{�)�}�ۂ�B�ZO�A[K+H�#�h�$�	�l�Ǯ{{bJ$��F�����0�1���$UM�\t�0IE!�B)l���4�ʫu�1�3�<������oS��x����(-���&�CCضg�T/��ƍ�,+G��f\�� !^d���Xy�U�Ǟ��z�K+� �P#p�ڲM�	��G��\[[oWD�]�v��G@U+L]?��M�1S,�1��}��{{Ee%>��1�o��@�~��[�J�)��~_�''��&��a�
�'A����K�4Y���TF:B!n����?��?�?؄EKc�k-���
%��R��v�kW�����Ѷ̶ɰBQ+�f�oZ��-�^<*^��S�-R�왳���##ؽk]H�!��֯��s18<�ǏH7)Q�>�bi�Ϸ{�g�<b��e�v%�N��m7�����^:0x��|�+X�p!�ە��H����FCjTI�vy���:1�LP"�������<*��v�B!�R�L�����)^?������Oc, �q�v��͟��2�^�c�n��Z�x	n�󓈜p�������|F�q�o����8�u�wn-
C$BM�wahp$�Y�v�4�"�|��煡'h�Ӛ��S�b����b)F��/D ��F�A�{��7´�0v�KW�ʉ��rP� B�ɧۡ�MV�א���BHV-��g>#%�:�������o|�hll�ϳ�ڮZT��6E�&������oI�j3V����Qj,�rO�4U���O݅����̩Ӓ�;� �M�P]�\�Vzr���f��k�Dd�'��Vb�;�d�oˇ�H1�Qa疏�kz���~멧�r�y!��dc{�c:S8Iܮ��R�ۓ�[�a�:���%Q�<E�k��p���vB!�BHq��Ӈ�+@c�,�;��1��h?{�����V��BG�S��ڤiZU���:4�O���V�ٝ�|bѢEX�j�aߑC4o#EG���p�����˪Q�����^���d�ڞT;Tc�9�����n��7G�A�
������*�9(�$��~�b�A�4�A�/6䠺c��t�tD�2�:�|KV9���M$����
$����c|���QVVf۵]��]�M��p쿤�6E�N�����ܛl@:y�X�vZ����ON����zά���#���� <���>��M��u��cz�t���a��#:Ǉ3�Xqm7� K"rf�C}[>�G
�=[w`xh$�� /����c��̼L>�{{��<!.h����)�d���B(�<Ġ)E���?LRB!�B��+�!L�/��.�˥������_2�jjj��i�i"�XÞ�E�_���G:����D!1q���*i����h�8�ͻ���b�Jw�<�>��O���ow�������{�D�PF�h��aXs/��j�����z�B�.�����?ͺa>B�{s�/�����`�5�����!��SJ'M���&:�������7�x�t����~��t�w�׿��x��O&/4-�Ά�n��4�u[hh("�)J5���.�V�m��-�+���%iz�p�M���;48$��@H6�E�֭���p��N�=cm�7����c�"�/�k�<bS�o���z)T�:��� ���k�Ib�̈́����:��x�ڹ]/I��*���!ɪ��rl:�$!�B!��8�W��{�<0�.�F���`h�+c������?����m��s�Ayy9)6�;;�I��7�p=�**q�B'���9�(q�x�f�̚3#�c8t�(�'�AH�2>6�[�J�'$�Zqݟ�v����2�A�0�+��>y4h�+�,d79譈�" �P�^�Oգ>�-]�V~�4i�x�Jvb�L>�r�A��EONViV�dU����J
 Ye�3�=�6mڄ��Q��g��&,Z���~{t�a�N�VbÆ�����Z�����.C��~�ɭ�/�&����NMM����uY��r�ףzZ5�FF��>��L7t��^��ƙ��%Q�����2kǻ�Xk"rz�{1X1]�!l?q�(�wx饗��M�M�{&����b����KR���A'��.'�􅘺\\}!�B!��������+c,@NI%jl�f��q�F�w�}4��#�Ò���{>%��	)F��ư�i�����7�r�UT���'��؝d��.]�s�χ��ͭ�q���;�Cwo�D��<�裒9����ro�ͱ���o�����C�(�iͰ4��u��p����|��gWG ��Sc�3 Rz���!C1р/�qc�%%��	+�EiE��e�7Y��g�E�c�=���� ��w��-�̙��+�'-�&�4g%������m�R��wuL�jr���N����T��܅�p*����PYV.9��kj���I�~^��j�_��RN�jF�Ʉ�׹�^�"�:����t�<����h�;�2C��سmgQ~w��O}
w�q�#I�|pYH�n9A��t��5I�ԉ�p�~U�k�UVU�g�~A�[!�B!���zMcISd>����
7�>�@����r�E;x�6n !�N�+�$�7g.��.�����y'���؝XF�/[����I�X�ζb��= �$8��	=�.�x���z<��3�y^�f=�@�cEEs�C͈ϲ)VP6�ү4�vy�ى�VL��'�C�P:�
i�$j�k���C����pc�I�>��/)Y�JX��(�udP�.�UNF�ɪ?��O�x�"H�#~�?����7�BccC|�%���tm7۬\�������ܺ�X�����
�m�A����Ϝ��WVV��O��Or2���!2��m�5kP[W�`�s�l�؛gW�n�rʵ=�eC�  ��IDATl"�hvV\�m��<��I�����9c疭�����<��+��M()�U"�M�v��
a��>2]�Jf0jPzm��ALU��w��uB!�B��=<<����$S,=c,�h��1���W�sh����vyޒ%K��O��?�!�7h>z\�s/]���(]�.J�@��o��NT�����?v\:��8.[���,FYE9ZεQ�N�mgZ�z��wx��g1o�<�_e۽]y�'n�d��%c�`B�nb��f�������3������C����>�H6�Tn�"wݡ#�/�$��am�V��*A]]^|�E|�{���9�?����k�c�tm׏�Q�F��3��)�76k{�Y�Zm��a�R��Ǎ����S�k��0k&���g$q�`� �;&Ő�@\#,\��W�@�*������V��m����\�Qlѻ�[�͇�H1"����;���x�'�|�V�ʻ�T&�ɖ{{b�:Yeֹ]5Ġ҅!�A1%����"��FB!�B�a81V9%�jc�tu�lc�j���C����\��ψ��=���������ދ��1Ca�E���/^�w~�S@(���}ӦM���(HqSSS������u�>�9׊-���b̕���Ň?�Ċ+��SOeT�K��u�Qc,����P[;L��:�X��1c,��Z����%�-@�
܋��ȕ`�z>BWΩ�L#t���nꄕ։AvqW���ɪ\~�G�������&o��ى_��Wx�+_V��s)X�"t�G�]�����iQ��uc͋E-�+K\��b8���A��	ާ���{�/�������L��ۋV�Z���֢��.r���.@{�<yL�wξ`��1�k��Xܛ�u�o���H�p��atu\ �s�Ε\����5�v(��:�v�ACq{.*�{䚤n�|�k���B!�R�l>�e�c�k�4�Jz-���o��oA��8>���<� **+A����i\�-���k�P�󣵵g#S1��q�[�h.^���
L�p�T3���3���a�G[9���>W*������;��.�굆X�{D�ڡa-Pa�7�
�`V�.^WT�c�y���
܋�-�{��k}��bP3̠R �n��$$Mʄ�ϧqbP$������gD���^�VBtA���� r���;��[�����m����ܦ(|W��&�oI��qk�@�4	J��X�b��n�����/_�bD�+WbF����bht��OCkg�&:���E���?�u�iIpo2�h[0�dl��G�����8q���I��ӧ;�(��N;�ɚ{�2)�K��6NVYua�'�8:X�0B!�B����mQ�n��c�4bw��'̱lc����5G��z��v��	�FGF$�����#���LNN�����kq�,�7��q*��11>��ǎa`���BA���\�e���O��`?�> ][B�#��w}�U��p�w���]�˧z��y	�XZ#,����X�L��)��Xf���~���H�C�{�02F�����@ii��`��L�������3�E�Ps`)��%IN�a�d�ӟ1Z~�u��/��/�_�
�;��CcC#�\{M�B��D���y���T¾��q{NE�ľ9�m�n�z^ @[������r���jl�č��sg���҂��)���q�L,_�\ri���111��p�+*f���)TTVi>�}���:��z}���Z�����C/و-D�z��i�.o�O|>���u7�ү'����{����A�.r�J���k����B!�B����YS�?��K��X�:���$��{���2�L>c�������̋{����8�w?���FB�#��:�IP[S���\��i�G�J�X��� �`ƌX�b���H紡��<s
m�1� �����	�w�Aow�w#U����5�\��ݪ+&���Xr��ԵC���|ߙ��M���c��p@��-�cK;���C������t��M9�pc�]܃A��#����� '�r���g�NV�Y�׾�5lٲ��� ��?�9���k�7^t��E�n���: l7h@6D��m���m
X�ؤ^7���b_��p�#!x畹����U�#G�_S��u�--�����K�`��E��������L�'X�=��Ll�]�5�F�k��u*�ccر�#���1�}�po��XIy!���v�$U($�0Ӻ0�I��f^���H( �B!���D�b��]�˰f��a)̱����V(�˥vqW�3"z�Hc�������_�"�����;�4�Bm}V^}!�14<��C��kkj�d�Rlhh�F�LM�|�9�;w��y���Ι3K�.EeU�8�a`x'[[1<2BHv8y��ZZA��3�<#�`�f���:�նd�X��XH�������+��~����aY�bwӽ�P�^Dt�Q5o>ƮtYrP\�����J=�bP9��t/��;�3�5k�{�9������4eee�6m�B�%��ɢ��,>���w�ug䦭Jg��{^�x	�� �F��H�~�/]���oɒx1��]]FEe%�	Xu�f�M���˗q��XŬ�5��vll�CCL�-�w-��ݗ��|�8�n��� �`��=�h>~2�J�D�'q\�~Z�8���A��zD�]�s������0��!��Abߋv��@����n19��n_�����1}�tL��������t3���v��.��1��T���+ǻ�d�F�.r�oE�n�M��K��S��>�om3�����,�@���Orw*-+��Nd�os���������GǤb�@|���?�-n�O�8)��������[�xN\cY���K�#�<�6�Ny[�VL0�ޮ~V	ۣ��p!��
���$UM�t���vB!�BQ��˟�1V�>-�1VT�l��́1�a{�c}��4�����CuM5�-\ B�}���p�d�V(t�.��w}Rʣ�ĥ��R-lpp�Y���1�|̚3%����.vb߱C��i!� j���s���W���<7D�N_��gǽ]Y7L)L�%ʦXAS�v���B;���i	�^��"cwO�Er��/'�R��eG��|����&��uqϕ�SɬG}���=
'���q�����+���9���.M{����Gy�Z`$������5W���wm7�֡�!�Z��T�i�]�N��c�����I+�9�6��
���V�]���4�DOw7��\��Z�V:���(��X�����]m�R�F�G"�_[�����1P?��lX���Zi��l ��K�q��qId..n ���&�����ݾ���*��+�G������}�s�Wr��Z��~����xי'��kkPSW����$��X�Yc����H��`�KǠz��T@����`����+�3}�F@�̊���M����F8�Ϟ?ב�&c��nth�sg�&��1k���>�{��Bߕ���/�;���DaA\c��8����ˆH�h&I�n�ׄ�2V������\�ɨPP9Ԡ~�*>_����` 13�X!�B!DI�H��K�Rc	w�ce�|�����/������4�8�-�wy%��v�m1i�s�p�� �PQY�6Vĵ�n���Y������S&9n}w��?�c����������TK�!��E�cU��,zr�ꄢ�%ȔN�b�h!�w˨e` r̷���m�ω�o&�/j�������_�W���n�ik�h�`�
C�Ҷ��Ν��߽y@4	3@7(��V<�������~w���3��[�}�%�n����[�Ш8Q�sω=7��z�B��]i���KU/L̯l��+g(n�
��AܺbF�.K���T�ܣb�`d�:2(;���KVes�����ꫯJ��'y�o����������+�����'��O@���N�f���"rk�o�?:<X�8+�L��+�{EE%*++��f�j^�S4��k�v���(�&3��+ȸMz����{yE�鄁�}�m��ݕ��'r�����G��6��:=rðj��(���W�Z����@�#�@� zzz�iddN!@e�_r�����pK��{����>�E���A��1�\���]����>k�D����uY;��ņ��w�l_�=:�a��5۷� ���K�.-�l�,e\t�v��dD��lr8��vA ��t�	�cI��>�w?:�;l���k,�z߭�y})�ͳg�v5�de�v>cڽ=6���$��*Ɂ!:iE��$��������vWL!�B!z����1V V7LU?�c	a{�����(F�{��wq��������<y*���+��/r��K)��-�N��>��&'DoKW������^�u�m�������{�H�Nolpe�Ű�+*���5�7{�T/��9v��%��E��!n_�t)�@�ubT��.SUU%�g͞���ӥ���y2�y�"�"�R_YU���d���f~B0�c��ݏK�p���qe�mE�ߊ�]���l��w�b���d�)�Z��k,�n�n}�[n���w����|5�J���ͱd���$Kq���$+j���1Ɗ�����`�>X�8X;�
�!G�����!���?���p�Q��r�HJ��r`�M7݄�~���oA���#G���������z�E���X'�Vb�������� *5n�Ia�c�{�";�s�վ�7u�Ŀ}���|�t�;�Pŉ���͑\�++*�s��	G��ztt��C����G� ��B�E�_r���	Q��|�+���ҿ�����$�q�t3��i6x�������]e�x7����oؤ��n���y�jl��z�N�8	�=6l؀/|��8+�[�[�:Ie��Ҿ�s`�wb��C��z�Ae�J*T�-A0L�vB!�B���@7/�����1V��$9���1�$nE33�ʤ�X5�z�W�)�l�,�##���|�{]sR̈z^��sҤdxh K�.�5�VH�A	)�	����w�=�������n!j�bD1�W���ɓ��7�O�c����Ckg��������f[�v���}�פ��e�ŝ��:���/IȮ���'O�eqa{L�n��5{�BL������{+/���"�dw �.�����dG�ȁ,:Y1iQG�����&�|YMV	��^�Un��|7q�۹s'._��->ڴӧ��M��lQ�h2�����+J�C�����[��Tp�Dl�ž�D��/�b��e�J)�5��
3������ʊJ���J�!�B�'}V��"���yrrb�X��A�?��>��3:6*=�,����P^8��ϕ��I���p]�c%�)v���X&M������@/�.v(D���a|b"i߄��kD���Έ������;�~��|<�3]�8��	�{������R��g3I���Ʉ��%����u�$����=��r���$F��t�I*B!�BIő�,	^�7�ҩJSd�/�c�����X�e�&�oN����!�7Z~�7JN����A�E_��ݱ��y!��0�j��@o_�2���^?���쪕(�N)�F�����X�(FF�1<4�9*�ΝB� ����	VuM�+�dX�_q�E�+D��}�҃��˸�y�4!$�׃��n�@_?��xꩧ�v�ڜ��-�n=0�g�?�V$�+m�Pg�gف]6Ē��)D��I1�`u�%<z	
܋�։�莊�S82h��"	��dU\�HV�fC)�2���7�l�s�̙x饗�_������_Gn&k��ڵ����I���R�l>֒`��\G���`s�Y���W9�g�:6Wb_��2g���H=*T�S�Z;�E��P�1S���`�[k��m�d����k�q�̮Լ��j�N
���H1#�\��n�����x��'�~�zǓT�*t�&���q�*[����uA3Ġ��_��K�w!�B!$�k��F�$cɓ�'��V����"�U=(�������،�v�؁�/�x����8R} �n����F��z��JS*D-D��b��Ƃ�3���e�ҹQ�ʅ)���d�%�#1���wq�'����K|UU��'&Y�xr*�y����Fϗ�u�q��(zGq��Kzo�w%��?��CW��x�b<��s�y�VC���V�ە�X!�)�~�Pֹ*G|���5���V�۽�E���)<��cÃI����{�{�Mwe��D�yA��Rw����7�)^7�͛7c��� ��?�9^��KX�d��ޒX7G�vg������x\+���%v�&"�����V�j���k��U������w�&X7[د9�ۋ�W�v[��l�uC��<R�g1L�f�x��z���U�vNp­��gI'a�����J��Jvo73̠<�`ii��� E�N!�B!$F�T=�Q��9V:S�`��/sw�c\�1Ɗ.J��9e���.�3f���/��������h>v�Ӫ�j�� �x�Oˮ�@���^�ԅ���B�8q�(Z�O�xq���o|uuu�����=.`���R�ci����J����X��@�ܣ��)��i�������i4�1p���INFn�v]�u�U@R�J�ٕx>��r��_�u�߿ccc �B�����_ŬY��L�Js)V6�S��6g=ָ�&��C��
X͋}aK�k�]�q��H�wq@�������e�x�V~W�`Wnk�7�k{rX~�G����	l۴�c� �C\����zWD����J$���̹��vaH��-���3�k\����@!�B!f�{Ac5`lx(!P�b)���^�1��ϸe����cӦMضm��8�t UUӰp�bB!�hi?ۆc�x�x w�}���Vn�e���bv�~/3�v�1��k��KY3���f����{
܋��<�d����+�U�F< �۳�������U������իW��_�2����{����G���x��WQ[[�i��͑�=lO�l_�k뀸=�"r���V�����>����M��h����T�:�ry���3��W�v��k;���?�ÃC ����ý�ޛ�$��I,{�ǧ�=�F��MN�IV��T:�Z��f�A���� �B!�b�󁙘���͚bY1�*)�E�U�Cc�_.��p��X��� �B��lہ��
̞;�B!2��.b��] �D�����+����!�S��S,e��h��t��F5De�P�ό� �۽	�E���*�5���]$O����:�g��R���v��L���~�����q��i���ׇ�|��x��PQQ����\ۓ�s)V6��-"7������������žV�e.ΚX8sa��X�������a��ߕ��6����V~�6����aa���k���#���Jw�7����kI�܈�3qoONRe$l��Q�$U
a�ֽ=���oX��n��B!�B��H.�Qc,�!V@�⮬�5�*)��W
�i�em�ʕ+���O�����A�����ܲ��̽��>�B!}����6�:�x��^z	�-r�F�d1�g�k�Ɏ����F~N�O�ޞ�n(���x���v�B�{��LVŇ����]ϑ�L�J�R%�����&��I����
N��h���Ւ#�[o�%�{�=:;.�g?�1�~���;#l��،u@��h��ľ��Y���m��0ڼ��l�V���	������^lA��[i�����ۍٷs:�;@��8����X�x1���J�<���0�k�U�Ĕ�}P��
��������~l�aF!�B!�lD}�+�)�9�d�{t~v��
]خ\�����1�ɓ'A����$�o��~�~TVU�B!����0�m�,]o�a�<��cyU#tG螬�1W+�^KN��XA���ں���L6���ޅw�JV�\܅�ƍ���=�^���&�R$�"�O��dUt�ۉ''�if�m�݆�~������MZϴ��?�',[���\۝���X-lߴ�7��{{�v��ۮ�F����&���kr�s"r'��v�wk��Q6��Vb�濫�!r�_�gl1rd��E��wY�v-���/�U*�I�D
�Iߍ��{�*e0Ġi�����fD!�B!���#�G���Ȑ�+��{�ߘ)V�+��9Z7L���XJ�,�C�	����䋉U&�4����*����9�>����>������B!�����}�c�c ޤ��o��&�������۔8m\�Y���a8�di�g�1V(�� ��
�I,Y5�#��.��d*Y�%����LV9��ufs�x-�U�w�Fww7�79y�8�&&q�'oW] �V�l>֎(�86�bes��D��������m��:m����(6����m�B��F�����Z��-�.,	��g��[���z!	N>��c'@��HN���ۨ����s:I�ny���$�R�0�JR�b�ȅA<����/�Z�	!�B!$S.c�ܗ�5�`�y���9Vd��+1�s�1��}�b~��4�~趉�NlS+��y���7��&��ضi�._B!�±}�bhpĻ<�����,�����ν=q��5���5ŊNA�Xto/\(p'�3Q��MV�M%�"��KViUJQ�V�+pqRˌ��9ud�d��ٳ��o���.�w�|�������?�c���X���D�v�f�i��L�+��ޮ�c�~W����uLD��_s��n�3�tm��`�����4�Ʊ��A�ͳ�>�����4I�F+�:�T�\�U&.V�TF.��K0�Mq;!�B!��a�cc,��{�f�_���{��`d�'��5C;�X����5�c��{����ě\��EYi��Z9^� �BH�#��?��W�@��ҥK��/���F�fQ��W�g�eT;jꅉ���a-��
܉D��*����bSP�̴�*�2Q�x��,�>�Kɪt��A�ne�C=��۷�����.���@MM-��.S�/:#`ͥX�^�~[-�+�����V�����LG~+�`�X������n��vm����$X7g�].?�b%��vs��m��=M �檫��W��U�$��I�l���[���J�����	�S	ܭ$��\��~|�B!�B!Y�+<��X��XA��(F{���BP��McA�WU椊�kƌ��7��w�yĻ���`���q�]wH�!�B
q���m�|Ļ�7��M��չ^t���&��R��bI�B�u0>�s|h���3"�
�x
�Ie����]�*7!|ɪHg�����i:��{�D�^�J���U���Ӊ#���t������Ž��	��� ����ǴiU���cr)^tB�k�]��{��&l6�}�ޜ
���/J5�]mÍb�z¬�݁�꜈܊�^g�#�{`WD�����4-�7�<]ۉ�K�]ػ}����;o��v�m���&��-7^g"A�c"A���R��HRI��{Ҁ�{�H7�7B!�B�;ڧLc��
c���Q����'p�d����K���{�̱���?�x����۱7�~K�\!�B����۳m.^��6�>�(�㎼��Z螸oӘc)�!��hv�g��=�R
��5�3��y��
�Im�J���6Q%'��	�H����d����OV%92@-p����J2���ϟ�W_}����@�Ϳ��_QVV��6nHZ朰9sq�mn�v�[�q��[��Tp�Dl.žf�d�N��ڦ8��wuFDn�����|Ws�����r�8ЏP�m��]�c���u.�6O?�4n��Fx)	��$�n�*�dօANRE]�e���I��PZ�Öv��!�B!�;t�g�.�1��n�o�ҭz��n�1�ۗ����ۇ�/�x�s�gQQY��7n!�B
������<��Y�p!^z�%ռ��«�_�O�ꆖj�s���=1i�i��ۂ��{{a@�;Q������:�{�2Y�OVE�4��Һ1@�Z�O�OV�M,�˂��Gy[�nŖ-[@�Ϳ��/Q�+���I�s)lvB�k�]Fq�Xu��ir_Ym���vY��|�iC�����pm�ݼM���X��p��|�� �"r�ǻ�8� G�Wa��}���:��;��=ر�c�:�x�U�V�^P�s:�dkv�sI��bBJ9A�LV��T3��UtJ���qo��%�B!��Mv�O�E��a��{�W3�����;i��+�l�o���x�����~�9<�s��I�����ցB!���}�z�������ַ��А�5�t˳UCL���̛b����X�b��a����D��� ����Ã�d�*Qe 4�&�CJ����U�ӑ�L��� �K$'�F�*%�$\7��L����W�C���������%%��\���gl����R�l/V�����\>�`�fŵ]3ۑ�J4X�Uf��ι�g.87�Wf�oi[0 ��y'\ۭ�Zܛ�3ږ�8������I���1jڏ�o���x�W\o����4I�+g{I��ܓE�	�3�*���b*+�cS;!�B!�8���#��qwq_��c�
����h�Pi�U��7�
��c�Q��*� \�E}�h��>(c��O�6����k�_B!�x����Ա �G���y�y[#�E�j�PO�.&=S��#{�����t�b:;E��B�w�ĩ��\��ڵBw=�A���/����dUII����ua���P	ܕI��]۩�p=��F��-�׿�u�����@������?Ǔ�|�פ����t��D���;�M�5�"rb_�X��]q=���?�"�,�9���J��n�9q���ݠ�s�A��{�M9"Bw*� �W��~�SSS �����-����$��$���'N*�ۍ�T"9��T	*Iܮ^0_@�aF��N!�B!��4�R9�+G�N���A?|¡=�F~����X%P>�4�����(���Wu1a{���HUK|��7%c�K�.�x�cK�?_}�ZB!Ļt_��s�gA�ς��+��լ��ܮګ!����(5���Za{jS,1�s(a�%Mi�Iu� �f������$up�����R%�dwI�KT��jGw���&��bw��aMG*w��y�L,��f��_���Ȱm�6o#��_���x�٧q�իuc�
s&��Ю�X�f��ka_e��ᤰ\�R�׬���j��:m��m
֭��M���C#������k{�D���\�S�n���~|��QV�۫B`ٲex饗T�
=I��<!\�bJ/nO���VJ9I%����k�������gB!�B��D��zMc�uÄ9��K9�s�K[/�k��$���6ƚ7o�d�����f~� n���Zk~�gB!����N���e�#��_�u̚5��̰�����L�Rdc��4#>��
c�c#3"��!]!A���`�/G��D�2Y%��+�Vqa{ܑAt8%�$UB�LV�"�'�d�{�d�]a����pQ��\�Z�-�y��8q��� �F��ӟ�+�=��+V����;&`�)��6�u������V��K��������oC��9�v�+p"���*�ǻ����o���$C����������� ������QWWWTI*�r�	*��[rp���bw�[{��������1YN!�B!�9�1֪es06xEe���i��^����!���	��XJS,�1��^�c�|�+���L�6m��}�; _��Zy�U �B�w8}�$�D����� �������_�fX֖�SlN�{:S�ĨωZa(6iGz6����6���V��*0�.�zX�b.F��S:2(��j7B�`<i%:�D�x-��:2��hE1R���9%����ƺ�b.\��^{����(J+ ĉ�g?�q\�n[D�+��v9&`5�}K^'�������)��+�ς�ּX�¶��n@��k8���`�ǻ�:���-���m����h�ُ�5Df����� ��3�<�[n��I*��4WG�n�y!�����`�A�}մj|p��vB!�B����,p9�K3��n菊��џ�I%nO�9I�Y�V�n��i�,�j������-;v/^�>�4I�,[��B�Μhơ�� �����曖�J���Ś]nv��{0�Y��!idg���Jc,i��K%rW�cB���5��@

܉!�z����r�SP:2�ĕ,f�
��Mv0�uc�%%���:�*ّA+p�]4�*iN�U��`%q��#����	��A��,r�`�U�����-�mp-ę+��t�Y�w�x�岀�8.�b_+�2km_; ���k��v9�]ͭ���n�̩k��88�������ׇ�� ���5k�}M5/���F��Zn���6Ġ�켠�'�0��I�v����{������@!�B!�@�K;��v�g�1���}��?� ˧�WL���W/E&�|��!
���Fbw�c�
����*�r�عs�⭷�¿�w��0طs�t\�XM'wB!$�ii>��{���G<<:s�̼���V���Q�c���P
���c��1�^�P;�s�h9Cq{!B�;1��?��W��ؕ.]G�N$���qd��yr�*1�`A+t7���Q�N5_���l���7��<x��� �G�|����K_yk��F7�PD�+�ѧD����E���C�{���W�u��p�v��3�[�+V6�x.E��(�7g�K�s�u���n��X'z1ؼ�u5}�W���͘���`����_��_cڴi�'����̓X�$�4�t�Jx�T.�@za�2IUS[���'at?H!�B!$�$cE�ϔ�C��=n��u����c��d�1��պ��>�ܹ���oA
����cb՚�A!������q��px�'p�]w���Jl��'��4�X�eP����c�ҍ��c�%�p8���@��w��m+pCyX��
7m'"'���x�*�Ŝ�J�z�DבA%r�Z�''��dU>&���,X��={6���oKO���G���;��g���O>���U-���R�k!Ζ��b�Y�w�x�eUpos��ͥ��l�>n{_g_�O�v��լ�����>�um��_e�d,Q��݃m�6cj��х��/��k���I*�$���~�Am�*�HN�sa�'��΅fE��c�B!�Br��+3Ē'�{:�n(��*S,�B�����tE�P������r~!���Ki�u��9�������I��ukA!�������c���R�PI.�~n���k녲9��ڡ�^�1�
&j�1c��|�)&z�&y~��E�<Mq{�B�;Iɥ� *V-�xO{\Ԯus׊ەw��Ȑpc�&��Wrr*���:����qd��i�l:6�����;��c�ᗿ�%Ha ���L}�Ql�x�����be�dEDn���^�������|��}mM�6g�ޜ>4����޶ۇе�|�ۂu
���s�2�o�SS�7�t�|�ɬ$����R#'����ҭ]��JNV�D�DSHG؞�ĠMRń�u�x�,�AB!�Bq�1V��K�n��
��_g�gq��5�J�F�!�S}��^W]C�Wa���Ϙ1���|�M��A
�c!9��n!��>��&R8���I����Ei��~��f�6�
��^����>�cik�w��β��� �	�$-�;JqG�/1�b�Ay�A����/��Tn�!�*��]ב�DUX���I��7�M��qdx�Wp���>}�p��_���w"w%9�Z�sB�nMDn �5)nwFp���v�ľf�d�q�b�����n����k>`�_0����k;1I�������X,$�O���|�;(//�]^Lnj�:Ae͉!�vl�b0*r���%��)�o���wB!�Bq#c,��]�n�0�
J#?�����F�P��k��O˳{뭷⩧��O~���A���q�n�B!�=ăg'�),��ylܸ�hͰ�u�dQ{�z�~�P�gu��ص]�*k���a e���}���B�w���� J,B���:I��jWԍAv0(�3�UQg����]�l��G֯MT�'�	�BsY�[__�o}�[x�7�.Z`��������ƛo��;#`ͥX�\�Q�Y���j=/`5�]��S$���Zi�~��6~���bs�Ј�{{�tm7�`��v�tu\����I׺���u/[�,��'+�NmK;�t�
�e��^�*�����$�ERJ���k�K�vB!�Bq�$c,�)�_�K��Q�ea���]k�%���
c,m�P�0(c�+��n��Ċ�/���d�u��Q�¡��q��s���@!���spOΜ<RXlذ�>�����/��-+��"we�PY/L�9$��
��k���:bd~ii)6��"�
�.�S|p��5T�9�+n�:2$����z��%�����h+w����\����zo��&��_�%�������o�ѱ1|�t�: ��爀�R,xs&�7�|���Ή}Ͷ������y��.m͆�=��u��+�����ݬ����Vb��o�>�϶�i�.隔��?>�����a!�I�t�R��k�JP�qbH��S1��ƠLRE&��4PiGQ �B!�7Ic�%��1�{@��T7�w�)�v�gu�Pk����'r`�#@;e���u9e�%�����o�����)N=���Il��ƴ�"B!�dq��o���i),jkk�Q����t�Z�0�1�y��u�䑟�\�U��ͱ�
a�4?0�����f�С���bl*��i�Q��j8�V�.�W��ew�h�Jv0��'%��ve�
��]�ɪ\
���v2�������СCػw/Ha��O`|l�>p�o-�D�+�ͥXY'>+"r��\��Nۣ�z�vžV�e>�����~�Nã��'���9�v�v�}��v��S�n�ph�>��dѢEҨG�>E�n�\�q�Jߵ=�HR�9190(RF�ve�JρA̯��g�P�N!�B!�����x�1a��4Ŋ����XZS,�޸n�4�sd����+��v������/����RX�4����>q�-�<!�B���.ݳu:Ν)<^�u�^�:oͰ��fo[	х�V����k��uG}����+놱��beU~�RP�NL�Q[��c�#�"w�$����/;�xMR9h(r��EJ^A+�R�28�Ȑ/ɨtɳ��r������y����;�n���y��O���-��gE�j�bs�4l�M��6��V�����8�؜>aAp����ᰅ��S���u��������o��\�aA\O�������.a֬Y'��rc�e��ȁ�8A��� '�B�2��/�HT���-��!	!�B!$? CUQ��b�+�+����퉺a��ݠf�CΡ�1��"y�mx��gq��alݺ��h?ۆ��n����#�BH�ײ;�lť�.��C���裏:V4�L���rum��K�~�5��3ƒ��Q��ͱ�������%�
������&�Z�0+0 i�4Ԡ$lW$��L�����rP��Ҿ�R1���{ul�����B��n��Δ����WU�������S�o���\پ�nuuuV�u�L~���5׮M�ʐ��t^�DӮݖ4�ר]`��+���뽒r�[��Z�|t��ȍƁ�}iV`e�fE�����FG1<4�.f�"l�t�PX����a�m����i�im���4:2*��=�=o����	���<r��:��M4�Jd��GO�ޘ����H��^�S�2+}~�n�/E�r�Tl��N�Z��u���`�+�b����z��0>:�����vڝa��M���D������]����9��k�l^gX��k,+�^to�����э�n�J߭�ع]��ҋܵ����%�롸�B!�B������z�������Jc��џCIuô�Xr]L!vO��X�XW����"g����hmmEW�Z�%�=�@n�[ۗn��gc�Bl��͸���#ksy��t��S汝��m��}ї��}�������&���}����u���nQ��;����oK���?55��[������y��k,e���k,+�~�x���9k�z����5C$��qm7�9�9V0f���W�����Sp�Br���������MRi�Ը2�_!|(jP)r7rP�����EC4f�+C��*+�n�,XIb=��طo��_�E����/���}Y�499�����>��]�����?��+*5K�_B�~��7�^�i'n�߲r�'�`�B]�ё����x��v���7���k��� z{z�l���Z`��TN�G������P��l���S�V��}���`�X�OXqm�zq��3on��n�l�Ѿ:q�(��vmR��m�h[��B�~��5�Ӟ��ŎNT�֠���DK��6���i��/�z����+þajr
]X�|���M[��]��9g������/]�m���J̞?� ��};v�|۹����5V��3� ���<��5���w���%���S��1�KR�3�q_HNVA����MV�0TTV��y(�B!�BH��%8=5������]���9��9�P��n(f)k~��X���&��9���K���s�J��~��q�����UUUp�Wrk�⻋I�?r��l}����ܼ˯Ziz
�{�q뻋<nW���P��k��藄I����]��pd��cc��OF�\��B�.�P�P���y���Hn��&&091��b>���vdx�"FI9{����-��ݾ�rs�b����)�73�7���=˿���3g�̉x=_j�Fˣ�Sl�A�P[7T��
�{0.n���H�4�slY����v��^,P�N,��W����h�#r�&��	�`l����];�`ԕAߍA�����G;^�s��s�@�溲!���|�M477��ѣ ��pr��?� O=�4jjd!�� �쵣ia{4�\���2k��7)̵)`�&��<.ulvž��F��]������n,�"�p�^���� ��+�;�Ě�m�A���m�9�sK�7Ļ?ކ��N�¤����***t��C���Z�`$hW��]�b�����T���0IE!�B!�ȡ�SX�|Ƅ1���]�k���~1O������亡Rخ�
i�Os/%yh#c,%�P��.�m�뮻��#��?���3n�&���_YY���)���NcMNM��ލiiFz���h�.\ 7���K�-��~�i���]�~1��˝QSW�i5��w�L�/a�Ⅾl_ț�.��;257���Z<P4k�W�`�q;<4���lK _��X�K�󸅙���+�ছn�k�s5B��DM��+]�PL����>k����55CQG�m���-��˜���U1�ۙHRiD�r�J��roW���C&;2$�1�ܣ�&�2h�UN%��-�E���jjj��|/��2FG�y�8���.|���{<��3�5{V�r�BIkbes��D�������Vž%ڇt���V���m2��"xgD��*��kǵ�(�����dlV���~�@a�;ǖ�~���+ ���&��e˖e%�TxI*��	q{����=�Z��J����B!��Q�^��5%=�{=IخqqOvr�Gk�:"�Ľ��nhd�%>�}X[�g�%)o�sQ�溲e�%�<'O�DSSH�!�r?��p�=wazC!�b�+=�R�pb|�0���[�r�g+��Z�\/���OV��ʚ���];�sP��rr�N��zv�L��͝�S�;P�N2bsG��E�Qr�J�ZύA9�V�.'���jG=7��]�.|Њ�ԮF�^wY����k���^�����0������ɧ���K�H�r+V�k�V�bߜ
�3�K��7�6.u���������pm7/X7�!��|g�0�������i������N2B�/l�`��/)\�x�	�{�YO6���l���H��3IR�LP����TCtU�` '�9� !�B!��;����a��˧c��4��5Ŋ������Fu�0QKT����ʆY����+z�\��X���*|��ߖ�����A
a���p˝w`�� �B�y�:.`���%CR��Q��~���9�fX�c��v(���^�P�KYC��S�c鹷����q���b�w�}c�Nh�B���K$��!	+��]��Ҋܕ�Ɏ�"w��+������1q����&����СCؾ};Ha21>�������_�UW�6�9���,��͋E-�}=/`5/Vv��<�Bd��F�Έȭ	�Э�߆�ݡ�Ftc-	��f�os�o���=z�{�c�G���.�AO�LfՁ�knV�T�T"A�.I�/xOva���Ӹ.���uU���p�CB!�B�'�X�����u:"wm�P�'L�*��N�rmP9����]4FQ7L�?�Xn	۵�W�Z�7�x����@
��T ;6��o���ZB!����L+���#]k��D�S��=���Vb�yz�v�	�z���=Q3L����Z0�Ҋ���~ljRg���$c�|.��ά�7�qq�KX%�%��q��,nOvd�{-�,����NTIsJ�;2�C���甯���s����R����?�'����q����/V�k��6)��"�Չ7ܺbSU����}�����.&�Ypm7�k"�|�� ��+�����Z����ݢ������B�SWW�����AmmmVSVב�X+m��3����+�Uz��PH� O!}Q{�vщnﮎ���B!�B��d��`½g�5Ø)����]��=^/L���X%I�v�~5��a>ce;�����/H�X�6m)L��o�n�����ցB!�?tD�Ha#�a�ﾜ��|.����Ê)6GY+Lc���#&�#?�������u�)�f,��e�ۋ
�I�L����?�HRe��.%���VF"w�9�SB�r��$�WFu�%���Ƞ]�f�w��믿���1��������Q�uϧ�cS�}���Xk"rb�|�ڊ͡��t���Z��I�$V6k,�\pn��r&��k�w��������e�:�7P��.gN6����ܷ���׽�W��zb*�r��JvbP:�+]B��v#���{{E�"t����B!�B�ğφ�9�059���c)E����h�P�9�1�@�.������9�����&���p��a��E��FGF��OH�!�B�k���p�������ǫ��j��M-�Ͱ���A�9V���ܕ5�T��t�XA��]���V�k���X����b˹ ����Ã��+V%�����=��23�`8��F_G;�h�N^e#�n���(3�'l1����������6t_����(*�˥yFb>G��a��w3�̱��^���J�v��	��	�ai[�b-}W�������[�׹��3��G��C{����S �ϓO>��~��y��2�l�!�I*�����Cl*++æv?8� !�B!�x��`���P5r���ݴ1VL�.�eq�c�D�Mm����Lb�~�h{b���|�;x�W088R���i���(n��(+/!�B"װSS���v\��	R�̜9S����:�uA��p+V;O]3��6�֥]׹=ͨ�qQ�A�P�=K��X��������^�t*�����\��{ّ!��J$�tE�vHI*��=�z�A�d��$�2��x-�\9}�4~�߀6�O6�'��<���t�[+���&"� ������w�/�5�&�u���Ní������[����r�x���,<a�m����{����w���� R�lܸ���ZV���в�^��&���ۃ
q�����
�������1t9B!�B!����|i�L�����6���}�Q��N�F"�T�X��f9�m�+۱�4�J��5k���������2/Y�\�Ѕ-����.�}~B!����0v|��|ȯ��b��e˖e���K3,+����R-��#��L�5ĠB�n\?L��{]�8�R�^�P�Nls�7��V.�ؕ.��=#w)a��ۃ
'�dq�*a%�MZ�eRՉ�آ8��`�Y��累�z�-���p��"�bg��������U��X-��M��mǰ]y+`5�]�tmOw��5�Z�}mW�l.�9y>
�a���U��w�߅��p�\ۣ��
�YD�>#�����G� )|�����i�\ML�C�l%��\���r�jjJ5��n:�?'�T�Y!�B!����f`U�7zߧuq5B!x7��^�pq��C��aJ�;27��D�^�X=��?�_�� ��@_?6��'�x�- �B���������s�<����h�{���Ųe�5n��n'��۱c�]����q'�7{��&q��-�Mb'��E��"�V�3��f4]���$H |A���_?��_�8$p�������E[k+H���_�:.��Ҵ��n�ͱɞ������fuC�`,���v�>��m���u�4�g34�Wx�X�/͕�U�Rܵ���Ƞ�T�X��Q��-��`p�V8�PY��;c��Rm�o߾X�r��v����w��Ԅ훷b��Q�>sf‴��m�}�2�[��X��,>V6ҩ�W~LV_B����#s�C���+2�po�`�}��������{ة9��^쌥���@����U6 �=V�Z�4���	SV�K���"���=E�����,�=�\;��t��B!�Bz.�;0w���W�}ƚa��^h������#���ڡi0�keU�ĤC���lƺ��;QQQ�6��nZ�[��;�0m�t�3�BH6q��!l\�!:C�&��w�y�ַ��[���`�a����OP���bi���������G��8PFs{�C�;q�ږN������D�J#H%�&�q��,�A��h�*%�A|�
�{�w8!�!6���Q2��7}�t�X��>�(�uY��{y���ŗ_��˗şH��ܢ6��{9�M������u�Z���������mwbnw�p�}ú;�y�������/,�Mv�Fs�&t����8�M��|�������&.���#Luw=�"U���^2�R�TS{<�!Uz{�wc���!c����vB!�B��~$�S��Tc{P��97e���f��S����y�u%��4����R��ѓj����x衇p뭷����w#L}��+wx�5o!��l`���ʃd�F�>���BW����o��V��J�JR7�q���Nmb{����F�{A���k�s���B�܉k�q�7�돖3g�b��ԟ������}�V����U�
�J��"�����.#�����g�g�������Z�:N?����


���Dn� �7}�t�}���6����]1�K�:1��l6�x_0����1��ذ�����o�I�X۽A�^wlފ�;v�d˗/WZ:����nû��P����<���Š��=77o+�:NތB!�B!��ƶN4�����xr���.��Zab�0�3���@ch3�{��`,�8k�XZ��	vw=��9a�<���(�TӬ@���46b��s��SB!�7�b���ء# �A~~>V�^��cǦ% ��6����x]PolO�e�On������n�ţ�t<�ڙ�Nhp'.�� ��:�C��D����hnO�ȠMqק1$3�KD��ஊVF�JY�"��e��]c�v��;�@YY6n���ޱ�+�p�>��*˜���ߣ6̾v����nS����gSj{d�3c�7&�L4���&r�72Xg�8�R��p��:�����B剓 ��ȑ#�r�J%�A�Fw'��c�w"����Bz{G���`B'����vB!�B�M�q�7��֦F]�P<�њa���њa(��J���܍uC�`,q���3��Z��'B~��_�d�fC]=λ����B!�7!n�����P_[�=�~��X�ti���UO�_&���2b��j����ϝ��B;�v�(�? ?$�>'�!���U������#�\{���nLb��U�D��`��McP�`%�	k�*�e63m�Ay"C&�QN��2����~����ѣGA����J<��_��[nI�86��0�z`����n>6�f_��d�M�fa������Æq�o.�lX�3��k55�{pӈt�N��n��K�/���g�$�hll��-�PWG�*�())Q������0ee=#����w�z��L�
�E�N�@��Tک�QR�9 �(RB!=����Ĥ��<�~Mc3�����e!��<�� ����Pm�����Is7�ۭ���]��)�f&�ȱ$�Rki�e~�e�QK��o��ػw/�{�=�젮�o��*ιp9��B!�7P_[���>A[kH�p��_���Z��uA���f�6�*�e��l%K��cu&7�'3�wv�����1��D�����;'���(�w1�Z��)w��n�b����Λ%2�1���99�Q�Fa͚5��������4�����w��EX~��'���XG�v��v_�|�S����6���ڃ����v;c�,�_��~�aYr���s\q;�q��&t��{=x�?ژR4 ���}�=�`��i�������*.T�E�pT��=$-�*�Z�23��$���0�� �BH�c՗.�]7/�|?�'���_�B�;!��@v�`�)��RsR�wY���n���)����F(3����w�6�ҭ�QMЭP+7B������#�(ɗ�4���ڰ���0k�\L�}!���̉��Q�g���F���3g��{�E^���������_���z!j�F��ՎϑyC0���Vh���â�c����v�w�:UM!�G�C���������X7����V�J0���ј���^�R���Cvƺ����c�/V��x�	���7�F]m-���ӊpiĺQԹ)U���{/��1�¡���1�lӱYءa=#L�����3�1��X�n�ph���װNc�w�����۰g�N�|S�Fz/_�җp�7����%�)N�����T:3�{"����G��r��	!���H���o\u�r���/��N!=�7�by�x����n��9�f��uj���,��=!K\�F�A��}�Xɶ7d�<��c����ǎ�Y������4��c��%��+!�ғ��:���Í8~�(Hv1x�`<��8p���@7�v���}�5���p,�P,m0V(V?L�eZ7��H0�����c]G!*4�OX{�׎*E[KK��`�`pO��I�*c���@%��2t-�Q?��I>�����2]�rc��믿^i;��?�$�ؾy+N?�>w����g�a��!�ސ�.=V�0�ߵ3ú�q^��~_a��6���������a����F��{��=1�3�=3��{_��"�����q�m��fn�4a��zFTS{�'$�T&�,���He�����ݿ(RB!=��?a���*_��b�����yI�y	!���Z;=�>�7�Gk��g��Ě���,�][3��@��H�0��n��il�n�k3�ټH�|���z��X]�d�*�Lc#ν�|��B�	4�i�o����Z�d"�}ժU�:uj�jz^m�ͱ��`�?#�2�	�?˂�B��ϝ���p�Q?4u�Lo'zhp'����cx���C(� Ms��U�D�@@op��4���(X���+�����l���]w݅cǎa��� �E�J<��_��ǔi��w�d��4�:4�:4����q���N��f���Dnq�w���o�ll:Sϥ۴�[g�/�����mX���[j�k��;�)B�>&L���+W����u�(S�����#R��ۥ"U�4��؞�ܮ�0x"��in'�Bz��~��/�e�_�|!�]�&�+��	!���ZE׍ꋶ�f��ݐ䮭ƌ��Rj��`(ftWk���������;@�c����ow=/��b��+�@YY�}�Y�좺�4^�e�s�29�BH&s��1l\����A�q�*B�.��b��~l�;ce����aX�B����`�`��,�=e��~����Dhp'���D7M����q��!�A+V��Uc{ "TE�E�$m�{��nfrW�*%�A+Z)�*eI��D��y!@Y5ډ����x��q����� �E[k����������/�T�{X5|���z������qfc��ߵ������{a��s\޼V���x���3�xKž2lٰ��QYJII	y��92m�t��)��H��,}!��S�J�0Oo�U��E*C���~���
!R%��B!$�)꫾t����+#/�I������1c��Xfwy�� rB9�za V3��U�j0VHW'hk����X�]��ڟ��X���wp��!���� م����[�9w��H�qB!�F���޶Cy����\~�����Z�ϫ ,��pg���]b�2��)�j=��eLm��
M����a(�Ζ�]׍Lo'���N<卣�8�_^L�2�2�&24���P��Z�*��b��`k9���4.^��Ȑ�t��lo���X�f��4515���G8q�8����������J�6lX�([���jl����t�n~\��)B}�`k�dr\��n�ܞ^ý�qfc{\j��qf��	Ǧ���8
'�!R�?��n:z�0Hv"�'z�!,X��w1�+q�;�ӟj�E*�$Y�Q�2m-hG��=/D�!�!��Ƨϙ�}�*d"�=�ƃ��x�E!=���A̘2-5'�>�5DmV��.�՚a@�HLqצ��b������h�{�D���X�XK������h2ǏǮ]�@���صu��U���KQPP B!$7bmX�>N?��̝;W9O��Km��DӻW��k��p,+u�x��������X�Q<tv�gݐȡ��xJ]k'�F�EA]������VB�2U9�e�XZC bp�ъU�R�J&X�ZF�*dP"COHg�7o��^<��� ����G��/��u7߈q�G��0�z`�M��5�f_��d����:�8�d����&����{;��a>m��fc���Ә���F�t�%�i�o�＇��z��E�/\}�����NaJ?��7�T	���ʘ�.�%�H���`�͠V��Η��e�!�����1C��)N�*kϠ����>EJ���M��ꕋ�)M�ҳX{� �W��]�U�{b�{��ܣY���|(v�,ȂX?������ ���[���ӠA����"���$�8q�^���8���<t!�?9]Y��Y�֖��d�СJ������Rt�.hwɞ��!�j6��k����ΤuC+�X����	3;�94��y�`�L��z]��\���\�J4�kS܍b��`�&2h[&&2º�{J���H6�u��ȑ#x��h��R�����������/����V/��}�=��jݬ�ɩ��֎�dޤ��7b�D���o����W&���_��ƍ�2��mX�w���8��nT�I�r����[oU�T�0��-tuwV�K��� TI�)Yz��0�D�Z{8�!���C�����Ϣ�8uJ�_����?!w���|�R|��L�&wqJ���O�;!���:�P4E��	]��5D}�{0�f���F�?�dŮ����o"W	(�1f��=���t{3f�P2W�ZE�.Kiij�;��^��ӧ�B�};wc���9�N
�f�L�<��Z�W����/~��<���&wY�P̧LoOQ7�.��b�Gu��q!,��^hp'iaC�@��Ztt}@i�۵FwU��&3��4����V�2&1Ėu���I���ԽD���2�2����w�m����/��H���{�D���p���g^<41��-�S�&M���}��i�������홅�7��D���{'۴�z��n:֖���X�oz�3֫�b�����O>ڀ#�d7���H`���8�M�N��۵g[��s��`\����IA��v���"!����ɭW+	�xm�~W�����2Mfr���$w��	!����� n�4��5�:��nh4��ꆁP�~��#m�0bt7��wH�z�{dU{�XZzc-��K/�ѣG�_�$;W�?ڈ�'��slkv�BHwikkæ�*]EHvs�]waٲe[t�.hoښ`<+fj��eu�����v�h��n��>��W�Y7$ɡ����C�A̛2Շ$i�C�hpWD*!V)�Z�J��`4��S�-U�
G?�ӑ�`w=?��V���Ã>�S�NaӦM �ˑC�������3�2}��I��^�#ce#�}-���k5ݗ�C-�����5��ȭ�����o}loHm�o�}s~zozq�M�=jNWc�{�q��Hv3z�h��?��|�2C�21�kE*�8��Vf-�Ȕ*�!�
V�����!��^�.���/��r����q�Ϟw�ܮ"L��<��뗚�&w1��y�&wB�!|P�s��E�����=Z�D��ω)����ƚ��XWR7�c4�{���6�3�կ~'O���������#����9矇!Æ�B�ʓ��������݈s��}�s�������6d�ˌ�aX&uCuj��?'��Z2s{��]�%y]e�����d��N��+�kF����-1�A�v01�!bj���S�U�p�ܵ-�P�2E��z?���J{�;���^Z[Z���	�/�%�]���|O��5����k��LVwlvnX�4f�C��pg�|�u��5la���s;�צ�-���arw��c���w�:���S�g/�m�̶�%%%x��G1a������D*c{A���(X�ZS�۵"�jt���!���ŤQ��䷮L9���_�8���ٱ<��k�V{�u�&�/_�P���N!=���!̟2A5KS7��Le&w��5���H0���Y��vHk���ab0V ��"�r�&�F�/fv�*�����Ǐcݺu �KKS3�]�&f̙��sg���!����=�wb����\|�Ÿ��L�9�0����2�^A�SQñ��C����˳4+h^743�ñ&�D9�$54����
�@�H��Z�Rڵ��JIm�ܓ�UZ�J[�5���T��Ƞ[;�(7��8?f�<�����;�����l��	�9�kn���=�.����X�H�f_���V�k�fe�c�3�g����؞��ng�s������;��=���l\����@�8�衇�hѢ�	PZ�����خ~j&3���0��
f	F�J�fP*Ti��(RB!=����ˊѧ� �����%%��k��k"��^w����	!�g�jE׍.U8���ܤ�X��a �Zu��U�;�u�x�0~���nOW�΍mtw?��Y\\�tݻ�s�N��E�}�ںU�*�d�y(.)!���MM���Q]YB�̙��~��kZ2����mĉ��5�N��C�����3VC4{XMn���S��uC�IRC�;I+�Ot�)��RsR���L[�)Q�{ fpW��D�J+X�S�]"CT����	&w��Tx!n���s��G��ի�/��T���s��k��EX|�����wFSk�v�f�LNmO=z�ޘ�3�p�d�f�k�72�`����Fg�o6֋��3�c����7(�~���~;���j����2���==Zc{�ܞ*}A+X�j�Amk�Dc�Q��ۃ�!���g/���SG����o���lG���o�*��^���~��?��w@!$�	v{ۇaL�AC��\������E��0��H����ƚ���VX��9Z7�c=+k�^�E���'�?�:�Њl���)�����xٹ9f4!�'=xX�v�{�5��F���{��^��`��񚠾fh��n���vh��nflW�C� v�C(L�!��$�y���(\���L��	V�x���&�!�X%H�Ȁ�K�D�G�S�exe`�2饗��ѣ��/~B���ۯ����e����A����O�0�ה�.���X��պ��� d�2�D�ý��N_�ߩ�ˡ9ߖ�^:�:��CG{����@����_��~��ʹ��_F�t���T�Jan�	Vj�A}�A}kA5�=e���k��H��u(B� !��sҿO�1"�}կ^A�Y��4��}Ҩ� ��3�q*��SFG��D��^����jpW놱���y�g�����b�BE��1������<K��D�ꊓ'OV��x�477�d7mmmX��;?y",9y���B�k��HII	֬Y�	&��������Y���u�XH^C4��uB㼾n�t6�
�������C�a�~�ۉux5A�NmK'ꇍGq}��Š*T��d&�@�����rbI�r�J+R�%2h���8Kd�� 姙�l��_�2�;���<����Y|��q��Y�1�X���{Cj���+����p������ՙaݹ	^��f7=��nnp�p/��g�홅h'�q�8�x��,[���{�r]�=��nu2c���l�����a�մ�&0����S{L�����D��!㱻��vB!�����w�y-m����}��;y$!��|�8V���Eꁚ��1�]\�����X7T��dݟ��B�k*OrWǨZ�{�XN�ᗙ�l����Ê+��SOQW%
�����J,^�C�!�b��Q/\�z5�>�l�k~^���-��BM1Z������e���a0�v(��l�vD���x퐰+w����N|�CA�2y8��N�����hnOl;Mtb�X%0�ݵ��
VP��Q�y"��Ft���"N"��>466��7ߴ�^^�??�Qʯ����_���w���/���;w��硸�HY��Ԅ��:�����[7��8���6���X�n�wf��t�II-����d�������[�^{C]�=s~�m�ؽ���vԛ�߳���T��ĉ{C}}�}Y;.{���D�������jٰn�D]*�nolhH�	;7BX;.����52�N9��X۽�x�g�����YGE�P�yK{{;�|^ڻ�曻>w���i�'.VS�vq�V�w?�U(?���$���>���χ_�y�������O��$~�$�L��-L���꒰������ۓ�jRۃ�-�UQq	^>�[��B�<�ob��S�Cs��!��P�B�б(�/ӥ��?�S�՚���5�Kꅪ�]`���ؖ4�=Ffc��=7�o��F?~�=�M�DA���]�&Ϙ����5B!Z:���vnݎ};w�<�����q�W�fnO����z�>�hjצ�'�ڵݝk��a01 ˬ���VN��vjz�4��x�D	���E(Y�A�ԮNc�U@Me�Ls�D!V���Q�h��D�`%�����*��vaa!V�Z���zlݺ��~�4����k�~��t���#8������a�СhinAcC�b�غ$�qc�~fӆz���|�E[��ܬ�M��O�e����mm�kO<9vh"���"�Q���v��ܺ����[��wb�M����l������ar>sƅ�s;{��{�޳u#��}%?~apW���3��kMv���Hji��õ%������;���?݈�w񹓗��Z�\�쵋���=�����w�Z���{ޭ�����M|Nn��9�?�8�����}v�X�"T�J�� KaH&TS۵U*QJL�F�c���dz;!��ۨoj�/��!�7Y8��'�@sm�i�gY�gm(����
h�?G��dwy�P�v�!�]yN+qfO0��y��q�m����/��2� ���������EO�?��뵧SG=v�0j*�0a�d��(�DHʉ#���n������D�o���߽��o��Wj"A��|�	�Ų����c�9>�PD�د߽�Ջ0��OzyO�����OIQQ�k��s�}�W�N��D�������������կ~Uw�\&�۽4�[݆�^h��YR7��e�Xj�gY���ܮ���aHq�3d^-���؇w��͝83l,
�*t"U�wm���堚��$��*B$�=�S�Z"�T*�����5k��������S�8�i�&��!T	����ɛ_�]��߽��[���Y��`�ĉ=v,����e~�:�|\dy]m-�M+e�Xm�ߵ3����_����������ʏK�5cƍ���:|���%��uu5vL��zj����/�W>뇍�r,\x�F�k>Z�2����7ld��m��-��Ò%}�����Ү��\"�Ю�w/>oR�!.��;0d�?mW;:�1x�Ю��/�����.���ڃ�[�)�^�
%~}��y������]|�t�������Į��"@���d���0���5"��X�����^�Ҷ���^2d6���N!��FN�4*��B�ۼq����S�3�ݟS���X��������o��ѥd5C�*\��n�R��\��]�Q�K�9�-����{�Euu5�}�]K��K���������kW�~�ڿ�϶O�`��0i�d��=h�����oȫS���e����j���(��p�|�o�]h��ί����]�ep�h~����&�����3�o>�D���طk�'�Cu��v��{�ﺡ_��<S�u�K.�w�u�'`��9����)|X�0��6�ai뇪��X;������A��Y�Pch�.���Û���e�xH�w�+o�IC�\_�`l�ލBUlL@�r0'�N"�*X�q�v0]BS:�.�H�|�'��ɓ'A��J���#K3fʹ��sS�u��s���c2٦U�sdp��ɍ�V��vƆ��c�پ,�ȅ��S��/���a��zeBw~�qq�Ѧ������{�1̛7/#��~������Gj\��='�&�P%K_�����4wM�BP�jдŠ$�]��=,9(RB!���:UB��Զt�a�X՗'��w�Fh�j�ܕZa4�],�u��j�9�5��녑e=�ޗ
7�)�Wy��X�۶mK�_�W���j&~���ӹ��������cJ(Va�?)ڂ����/~����������p ��������������}��w�����w�~���`,��멯���|���՞�[=?��6�1�~�����z�j�������L�3Ʊ���3l�ޞ�vhLmO��9����kK&w]�1�t܉�W�g�FL쪩]�~P"T��wE�Jh9h����^5�kJ����w~E���D\�R�%F����jf7��6m�br��{���B���[���E�(�ŗ^��b��Rn�����F94���=0���-�Ӝ�niG�&�ݹ�&8}_9����8[�e�F���oc�ݱ�>�奸�i����])�8}�}��.��ߦws"�v�H�
O	I�a��v�@%�Zs�����TA3�*:=�?g�)RB!���&���!��~�>�-�����>��$K;��5�Xj-Q��Y��Ko�LE�P���Y0�nK=��ne~���x��'���!Z��N+uC�C͘3˓dVB!�I::>��͔)S����[�n�'�����YV7ԇb�������X8�y��I-Q���2���3q ��wN6��2t�j*�,��'��Jd�?کN����U\�
�?��63����E����+�����f׶8PV��.�g͙�{ι)5�f_��d�M�fa;�ou�W&rٸ��M�ĥc���LHm�tL&vlη�Z�0��؞Y�"Ŧ�?Dc}�!�o��V�x�aV�D��R��A�J�ޮ����������JLK���'�!��^Ms�>B!���,�5�'��j���&�='����푀�x0V�T�'j�T硽v�h�ᰶ~hnrWɶZ�1c��SO��;�Du�w鬤g"��vE;@���\4�Bz7"�}�����6l�r�8r�Ȍ�����iq{?�uCՖ�։��u�X&�C�#�v(���t�vc����y��x�?��,����N2��+B�e�`47�%��R�c����]�Ȑ��.P�c�0�T�ct/���Pv�/��2�t�����?!2Z����__ā�r\t٧Ч��k�̾��_��fa��{��[v�;}����.h�ؚ9���;1�{eX���[:�.|7�	���wM�r�-��k_��o	M~�^���aӇ�{���P�Mk�	U]���B���h�̿{B!�7��ƛ�!�xKus'����ri �Hs7���X�I�w�#!�=Z/D�(�cuM#:�ZgT��Sk �ZK�1c���):�577�#�����k1���5.��	!�":>�ٱ{��dj;1E$�?���J�{&��Q����6����X74N���ꆲ0,i�0��0�7����*j��4���ლ���WI[P[��IdHl;�(V	T�K��������YKd�$�������,N�>����74�S��ڍ�r,���_�0�ɚ��d��]���3�[k��J����X��+���m���9�����	�������c�ؿu�u $W\qV�X�ܮ�|-~M�<�d�L��`4��MR�թ\��TRڃ&	Ʉ��`%�����DWB!������{B!���� n�<�u5�za�a�N���`,s���8�%�#�n��XV��=�\�Y�F��,��1"���;v����X�t	B!���&���W�����Ĝ��B<��#�?~F��3����J���Jr{b�3��9Yr{Bz��9�t�!��*�>���dG�C�=y<B���S��G�D��0%7�dSm�{\�
 2Dk.	@fr�᷁=���'��z�����������ގ�־���wⲫ���a�Ƹ��nѰ�Yj��͚���:6`\�Ny&�a�S�����u\�n�����a��voiin����p������$cٲeX�z�"Ve���Ix=���Pe�ª�=�<�]�b�3�b0
�[����1�3d^-�ٍB�Z�Y�"���U������V�0!�=����cm'�$)����	D��\�gc�{���/GUU~��S�%�����W�b�䉘�x��1�BH�D�@�����@SS1C�������K2�>���c�����>S��k�C����P����ܜ\�}BxB �)4�����!�4~Z�MM��$U�R1�*�R�܍b��^�\�Ҧ�k��[�N�W$r�}�ݨ����/�B�q��	����a�ًp��磠�@Y.�H��W�{�Z�x{f�$�u+cM���2��-����nB��ku~#�Cýt���uK�E�7U�ۏ���)���b�x��PZZ�"��x7��4�Am1�1�*�T��)z�*3�u	R�J�4�b�_P�7��"!��t��O!$=�h�}�x��V���k�j�0jn7���v��l냱������ֺ?���f�.����466◿�%Iơ�8u�$�,���&�BH��P�l��	�Z��ERr�w��n�vm�+2�Ψ�@2S{�$K��k���ڡ�n��c�C�L:?�@k�ɨ�bHq�IF!ğ������r"�~��ܞ�"w�M��T|��փ�yDl#*X�q��`*�)L�ݙ���W:�����o��d���'6�l�~\z��?Q&ZY3�:6���uh��gvjV�6�;����1܇-��oמ�ܡa��8��Non����>aܤ�&x�=��N�7����Xa֬Y���A�e�A=M��H�{��d����Θ@����a"T�.�����B!�dy�9 �B�����e����IjpO��D�9�wM`���] ��D녝b��Z/T-2�NЛC��!~����wp����3�[��֖l\��U`��g�o�~ ���45���n@剓 $������(�V�I׼�b�Z/t��Z�Ϋu���Iz�����ax���v�4���C$24���Z�*�U�����.��VF�*jt�<9ֈ�b-�!��f����X�fZZZ���T4�����#&N���.���ڀ��l?�M�VM�^��XwL��q�o.��/���kej���*�\`�W��,�xG{{;vmݎ�=��{&�?~<�|�I><#��~`��vui�.%S�*�@��"�v�P�
T��Z�W�hn'�B����|B!�Bc�U���iP�G��`n���a�v���?�L����Ѯ�j�PS7��]0Vo�+
�������܌���/ $�'O��_�Ysgc�Y3,�!��q�w�.�پS9w"�
��r����&|�gBm�����y}0Vb�g��]�ʦ��>��X)j�2s{^׵�ۧD�~����d$o�)��T{�R"�V�R���=�⮊U�&w񝠊LF�J����6��4u����Z2APJ�|߾}����������A��W���CX�d1�,]���x�c��X�\{fa�fe��v}>�c�1�;�?��p篵G����O�9�Oc�ݱ����`Yvlފ��6b��#G�駟VL� 8e¼9�B��؞L����#˂��`t�^�2
Vf�����|0�B�.�YR ��^��B�<��m�c�C����eqC��6F��.P��S%�=�^����j�^��熁]K����������T��֮]BR������T�/���a�� ���8z[6|��3g@�U���Z�s�=�ya&����ߞ��.��l|���[�Mo%�
��Fs����}�����X�]�F����%X�7/��`��`0&E����F�{�!0N���ӸȤMo��,'S�#�����z
=��m�B� N�6~���܅>u	�͘��W��S�u��Cs���ꉉܡ��޾`�U�S��������8����?7��l�߆u۽��T%�l؄��:bq����ӧOO�8�&��R%0Ȧ֓�5˂���Xr{�ւ&BU(ԁ���d�AB!$�`�;!�?Xw�7O��S�k�Zs�����e	��j��!�`�Ȑ�F�e1�|���?�0Z[[����+45���7�Q���^�Ҿ� ��g�e��8y�8�ç>�)<��(((�S��x�j��ݮ�qs{0I�дv(3�w��a�g�4������'����2t$Id�&1hS�uFw��=�� �M��b��*Nz������c1b{�1���C�@�U�.�^���`��	���K0h�`e9S����D�v�f�����X{&r�&zc�֏�����{�4�`��-8T~ �إ��T��3w�\WM�~Mn���Pe.N��������v!P�+��B����<;�hn'�B���B�	!����#��dP�r}����ż4�]ol��H��x=���YL�`,��]��;@3+�|�>}�f��\�6l !Vi�������S1{�<����B!�B�o�۹{��T΍�Ò%K��KJJ2�p�	����$��$ݞ��w}�P��������;L��E�x�H>��g�6<�'͆c�i�h�ԜH�)Z�"UL�
h�+��]�� ����U���"ȉJU.�쮁�O}w�;~�x%�S��9y�$������>�y�`�ҥ(*)���Ooj�4]ܡa=#L�����3�1��X{�{����eq��X��4�{�*N��z���L�Aqq1�x�	�w�y�o2APJ��;	�*��=>Ml/��خM`0�����?����'U�B!�ҿ��B�4��q�1<X&OpOR3T��j��Z7Tky�:!b�X�r�l���j�PS7��o0VO�8p��%j��w�!VZX��8~�(�.^�1�ǁB���@,�%��˜9s��O���Q���ym �6+�1�ǌ횺�ݮ�AC�0h��Y�vDk�ښ�:�`�ژ�N��w��|� W+FG[��؞��`�^�JLq_�JkrH�*�4���$���w��Ϙ1?���p�}��ĉ ��k�Ə�s�v,X���,A^A^��[4�{dl�l��e"�s��e��a	{&r���vƆ���!��{�Ą��Xb�{=v��}��MM �;��GŅ^h�$�X�ռ��@�.��+�F�T���"���Ik�L�jz�Y�����#�L�Ǎ�
��B!$[ط�B�_l>с��Ek���@,Y�P_3L��9��92�k��`,h�2�қ`,;5F�p�>O?��br///!v:�����C0w�BeJ!�]��N+����*�f͚���2$m��t���=^34>:�?���ܩ��������5�Ȳ�O�hn'�A�;�xZ::�?8cC�ʇ�,��htכ޵-�)��P���U@��`$`1u�A�e��	M�`TwSH���̙3�ar���0�O{{;>Z�>vmێ��/ǌY3��s[&r�f]�fa�fe�խ��0�;4�[ܗ=ý�qfcәz.ݦG7789&��~��.��f*O�ĶM�QW[B�K~~��V���.�,2e��ӻ�m��d	��vm�*X��0$�T�V�b�s�D����B�f��蝼4#��/��gF�A{kK�F$�j��j�P��	&w��'��f�Xq �eٝ`,;v?�n�رc�`�{ｗ&w�-���W�b̄q��p>����B�3�MD;�lS��	�.S�Nŏ~�#�9�3C��5?�ǥ5�k�>���±��:��%ʺ>��]��V����Gqi_��@. 
��;hp'=��:0y�8��>��nP���UZ�*'n�7��L��/�݅��S�7i�AU�Q�<�&�L�D���Ǹ���Q]]B�CcC#־�
�oނ�/�#F����p홅���7�{a��s\޼V��[��L������?��8u��aℼ�<<����k�
=�`2�{�nC�%s�>�!���O_P~N��`��BU߁���;B!�d'"��K�-Ŀ���B���]m�01T�܌�P7�>;>[��2�
�S%K������̞	u�t�Ǎ����TQQB��й�>�Iӧbּ9�/( !�{t��cώ]ؿkO�7EHw������3fL�0��a����%c��~���C(V�wy0����ʼ!K�-���<!co����^.���MMq�J���A�$wm�{N ��x��>��*m*�����tu{�pf�N�����?�r��0���׃��r��	����)ӧa���0p����c�3�ݑa�5��Dڞ�<��ƙ�������;iin��m�q����q�0�?���4�[�7۝&0��e��v%���ԞL�����ە���!����ۮ[�la�ޣ�`�!����߸B��-;�_XEqa>!�d/{���:e<�Շ�����f�7�'����fh��R܍Y1�ciɄ��߆�I�&)ݟE���#G@Hw�X��8\qg͛�IӦ*��B�#>?E�p疭hkm!N7/��:1�C{wM喙>'��	�R�V�>w�:���s9�'`_9���{hp'=��N`S�P��iR>4#�
9	�2�{d^/P���`�&���U����h1�ir�c�x�b%�A�hr'N)ۻ���c���X�|���{ީמ�ٙa���{G����Z6�{`7k˰nq��1Lv�	ݫ�����ػc�"��sB�"η��s�!�鎹=~�]\�R���L�jZ�i�n�T��&���"!�8A��ʧ�-tt}�|�'��7��}���_�	�~�Y�w����_��&�!������N\?�?Z�u�B5+Y���n�} ��]�����h���ac�Ygʔ)J��=�܃�Ǐ�����ֆ->F����1w�M��z"!�d�{�ء#ؾy�π������z
'N�V�/��������N��$5�d�Xj�0���I��]���X���
�8Hz����(�1u��Ք'��V�X%����8���9�J�v0�� �"w���I��t��V^�IB֒%K���+W����8A����Y��b΂y(--�-���t�|�d�S����N�
Lm�w#��X�����W����m��Q��}س}�bZ%�rss�b�
�r�-i���%@�"q�=�*uCb{A��`0�b0��U�*jr�J�����in'�b���\<�����O��W?�ɽ�Q�ؒr��#���_��t"n�����N�4�BH�'��ځ8��L$A0Z+�e���؀��YMs7� -P�S�!jk��`,��.��Q�JT�զ�g��]K�u�M����E�g�܉S�q�طs7fΙ�1ƁBH��'���ͨ��!n0b�<����M�=��翹=;C_?�����5Ci�g]8�y0VB�g5���i}����1�Iz����8^���#�T{*!�!���vP�̠m9�#��9�85���b�A���"�6�]��={�Ťt����ҥK��U�V����8E�mo��	��맜|�_��Iױ��,kbVv`nwj"��Z�]Im��/k�쌵g"w�n:֖a��X�7b���:S��Cm'�k�v���6�ban��������7ڻ{�^'0����*��bP+RE�������B������oƷ�<^�hH���܊o]�3�K:�W-��������]��Kp�˒�y��x��� !����Dc'��GIC��(7�Kñr��Xڟ�5C���`,�SM0V$K��J�{�:�v~�̙x��q�����
�8������w���D�n��Nc�'[Pu����0���'?��3,��2��矹]�q�E��$]�Շ��vyb0��n���b��>w��t
�W1L���I��#E�lh1:�ڢTb�A�@��7Ot7�1���@6U�ʌ�q�B�v�س�@FK^��.� ?��z�j&��'g�� [�.�.Y�9�梠Pot7{�[7;5+����Dn��k[4��7܇-����ü#s����-ý�qf��	��mX���]c��r��EsSqq���_��=3��[hr2/O`�$.$����`��)D��D�Ǳ�iڃL` ��}���W܌���Oi3A�tt�K|�g�c�3�FQ�y	A�����bǁ�8|���cz�㮛�'#��>�<:B� ��=�{8����FK��x��f���.ꆱ4�@@7�ĊeɃ�T�;ľ�Bc0V�t@�	�f����E&��gϞ��E�{uu5qa�lmnAmMf/����B�����ؼ��� !n2r�H��>k֬�4����n�.Q녩ñ��v�`,IH���Ϛp�����J��$���Nz$g�;�?8�:+�mL��y�@��"�H�;���@�ʀ�(�R�úm�m`�û�e˖)�=�M��UDz��＇�?܀y�b�����ݳ�v��iJm�gwf�wÄ.]�����n��L6�Jj�a��QzeX��=��;�8z�0��؍3�� �mĹ�+��/|�Ss�ߦt�捩��H*��v{	r�J���T�����.��&����vB!�����/��}�y���n�����U��o��Ƿ^�t܀�"<��-���ߢ�ݛs���"����I���N!�͋�}���"��lV/���1�����������Y���x�~���?�ɔz��ǔj������<� *+�2K����c�c�ј5B魈.����у�A�ۨ��~�ۓ�W�P�&�hl7Io7Ȓ�u�X��a�@,Ӯ�Qs{QI�t0I3�x�ǲ�T&L���Cq� Z%3�'$o;(0
V�w�f02,����{��ݎ��t[�{��ʰr�J��y�E����6l��>Q���-@aA<���,l\�Ԭlc�w&�L4�;�8�ܮ����.��9߳�v�64����P=r��v�Qn���M^^|�A�x㍮�ۍ�mJwk^���x
�F��el��.�$0���*������c9��B�C��u�͸������3x��MX>w�9ﬤ��N���~��_�ۗx�}�B��������BH[0���C1-|P��5��ljv�	Ħ9ڟj�F�{��]�cA�����fBݯ;��t��Ν���E0ֱc�@����N�ʹ����w���N<c��ъ�묳�J��݈�uA+�zc���.��Sw~6�
F:=�u�P4 +dRC4��,�ak��.�I�����h^��������Z#B�[�	V9:�*� V%��b�1�]��F�X*�X7.��{o2�kq[�:�s�ӟ�T��z�xA����f,<{fϟ�$�'`��n��끉<�؀a\��lӥ�s+���zps���7녹�+�<1���<�@Y9�l߅��f����/���W��n��W�(��{=���ęU�������Tg��P0h*Pi�j*�(,*�ߏ�	��^Zۃ�#(��EIQ���N�4�� _I�����?�u}��T'��~H�����7��>~����n�h[ڰꗯ(�8n R�����I���N!D��:�)�ǣ�����sN�4�d�H��1�]npW�\�`��~���y&w;�t7k�"��g�Q�܏9B�Fkt?k�L�;!��&��VU���	�x����s��i�|1�gB���v5��v}�c�C��Za(	��Χ�ʻ>Ob�g�4���0��}�KK�TY��*P��D�J+\A3/o;���݅9��.�H�q@k�Ӧ�G~O���3S�J��%{nѢE�`%�B�z�xE[k+>xo=>ް���ż�PRZ�Jj�U#�w&r���S�}u����wj���rhηe���ƄNs{z�>��+�w�0���/),,�#�<�����U����N��V���I�Z��?Sۍ	:s��H��;$U�����6�T��n���w��/�G& Һ���)ǉ�{�o�w�M�q�d-��)����z\~�4�:y�9��{nT�_�g�N�̧���������@QA�r��?�W.��vҜ��;v؀�chn'�b���N�2y�j+����Qc��!��}h���=G[/��]SY0V$K���&w-^��O��c	����L�%ޠ�G���sgc��� ���Bu�i�پS�����x�ĉ���'ONKMЈ�fu���0,Ӯ�����e'�]]�a5)�J-1U�gY��!���2v�'�A�;��T5�pr�Xj+3Mq7
TV�*y��ؼؗI*Cm�����t���y�#ar?u����v|�a���>c�Y��x!�W�������s{�|k�1ۗ����������n�Dnzs�l}�XK���7������!�|�~�߽�� �k����f�\y�=�ܞ��TI��p�Zv��Z�d)�;h"����N!$5w��_�Ζ
�n�-�oj�W��/<�K�Γ���܅n���v�d>�+N���7�+nH9v��H4�B1��%�h@�r���fh�^7�[�j��z�1Kot�&w7넩�%B���Q1������8v���2l(��>KIv'��L���
{v��	�S�*��&LH���o���y�f�7��S�e�X�k������
:���ϯ�㩿�����
6��SƢ���i"C���wS�;�r�$�AO<�A]7b��2\��=7w�ܘ`u��Q�%��o���c�X�d1��8Іa�y&�a�u��pj7kٰ.]����2gϠl�^�W�|F����s�W\��B������ԈT���!s�J+LY0�ǒ�%)����
B!���;ۻ�K������߽���<��OI����V܀����m ���]��c��Ǫ/]�����N!$)u-!0
Ãe)k�v��j���]��Y�*)��h0VB���jlW�[�N�/���4�O�8QIr�X���!^r��
��|G	Ě:k�Mԛ�!�/�w��cǱ{�Ԝ�!�@t��cǎMKM����0A��Y���!Z��v���h�0�P;4�ծύ��L|�w�kx�"׍폖3�1I�n0���`�vИ�)�iE*�pe��5�DЦ��7��H&�C�܌3���z��I�(߷_y�?�/���l����~�O��f��3֩�ܙaݖ�܃�\1�K��oB��=}�V��w�Q�b��$�_�~x���q�d���ܘ�S�O��0H�Z�E���ݮ�]��`La����ۧ"��3�B��_X�֎ ���������N�����4���ן֡��߿i�o���wᶟ�@s;!���l>�uS&�����f�c����������5Cm�PE1�#^/�w��MF�����3�Nh����0a�y��\��v�!^SW[���>���1e�tL�:��� ��t#jGR��gAH��9s���>f���xF�c>�}0���.Mo�P7L��Tj�A��v]r�!�=g�$l-��������	���������Pe�� �?��Z01�!�t�9�w5�!2&"�DZ*si7��axw��.�܅`�o�>�.�:�<DB��ys0c�,�(����v{���p���Im�n��e�:���n�po:�_�:��CM\�EKAB�������SO���v,JqSd��Ю�W�)��].Ti��*�H��TJr�=s�Q�R��b��P��B!�m~���PR�o��-L�:e�_on�|~�oo(S?L�"���vB!Vy�<�'BsC��f��J��n��ꂑ4wm�P<dI��pT�b1,.��7�H:���:"9T��V�^�m�x�$I���c��]�2s&M����BB�״���B���ݏ��V�N,X����1b����tڽ��S��I��G���#?%��!������ϥ���r�<Hf@�;�U�h�x���T�,�4[�}���P��� ��RD,$���S""��j����=��[�L�8?����裏b��ݰ���^�_�Ȑ����}��/����/Ӈ�݋��n�vqb����رe��<


�4Jm�mhmnQa�/����@юL�������K�HuHb�¤kwg�_��Ȗ�߻��MҒ͎������^�{���ֶk�B����ZT��oe��mZ��L���=?h�������[�345�Q.
��ٵn}]]�{�F�����������~~ר�t~���گJ�wQ7>|�r�5{�l���q�"ju_�R���ZIo�	VR�J1�����O`��O�hn'��"��_�"�q�y�����{WaK�q��G�܋
��k�I�>��N!�.����+�ci����X34v�R+LU34�
��X���`d�z�|zM��zQ'�Ώ=ZIr�ᇱa��.Z[Z�㓭صe;�N�ig�D��@!nS_[���p���rBH�Y�l{�14ȳ�^wֱ�]��!��k�� \��j�0E(�xN���R~��ۃ!��X��aA~>^?Q�u=E�d4��^Ǧc�v�xt���B2$���%�OhD������dE�RS�)�P��Qѩjt(_d���v7'�ūQ�F�駟VX�֭�T�W{{;�@��kէO455�����b�����W�����br�N����c���	f�ƆT�>��&ꖛ{O%&r;�p��;wc���}���t_�Ǌ�QO����Im�.��:�|.>�z�y��k5Mm�"��M��X7X���?���M1ۢ-�ݱU'O����O�R��0�O�:ٗ}��SG�c����i�o��={#�T�Y����������[+����ɼէ�
?_��������a�ԩ%J9]�+,�6e����zc���	T����`4��O����k$�B�����9~>�P~}"t�A�J@zk~�w��𭫗x�/��	!�t������)�?�1��5ø�]�hpW��S������jz��{_�g/�2d~���'���~�-Q��
�;��p*?�R��M�i|X��K�1p�`���k�+�P,A]M-���ǀ ��/�kk��RX�]�kp� ̎�MMhok�e��&���v��3���]����[�練�������x�
D�.�����~�
��-�X˗/W�唖�zV���:�fh�����O�w~քbj��S�������ۃ�������	�ma0�hp'�����i�`45�F��I�)� �A�BJLd0�S���F#�Ơ���v�����='�-p�c�ڵ ��{rߞ��cА��9kf̞�u��P����[2پ����Ec�sý��`q����f5��e"�e��3֡�^:�}úW&x�}�<v�w�E剓 �ofΜ���Ǎ�(e�?�z������v�Im�br׊R�H�.����w�e��`x�"�k�K���F1һ7| &����f�8��߯��8g�8e~�#hmwv�!�������m��y��U�{��տz��TaΤ����t]���w��{x�B!�{l?с�J0��x�Ϥf�c������;�k��iL'HHqWuUu���Yݟ��V�q���S�E�z�)���˰BQQ�����g0�x��_KK�/��;,ī�����S����~H�&MH08
��`��A�?�������%�}|�����o�L�J8ըqc|�����1b�(��tS���;aN�����<3���J�P5�;��~�Z�� �>� �k��ʕ+�s&/k�n����)��Wk�zc�$K��9U8V�`,%KIp77�kk�f����8;*hn'��W"��=�l�����Z������[�փ��t)�5��p¶R�n�ʭ}�5N�??����U�򗿀?�9]��＋M~�ig���ٳt) �M�f�p���������>ֱ1��ذ�����5,��?�7���nѶT$���݇��f�	,\�P�ap��ᾋR�Yǩ�ݙH�OmW1ڭ	TZc�^���/%���)��U������V�T�wq�����7�oI�F�?؍5�Y�cU��D.Y8O}�JL)h�>T�����n��靈����X0u4H��w�~B!$�y�<��'CSmUb��]c;��CM�;��c�t�h��R7�uYqTc{d^����v��v���5k�(]�_x����7Dw��mĎO�`���4}*B1���������v0����?�y�X�B�Q+Sk�F�7��KL�>'Io7�!&�
�܃��ꆚ�a���c&H�A�;�Եvb�(��<�|(���bL�����Fw��] �'��6�|�i�ܭ%2$#BV&�܅P%�-q��?���񝶶6l߼Uy1�ƌ��c%w�;5����%��7����Dn��ō�2��2����p/�	��v��'��Q���U.:	��-[���]���:~	\qaJ�,ǖwjR�%$/�甶�Am�AU�
�No�̫bUp�$�b�e��Ogn|f�L\0o�]�[�<�I|��%x�[WB�Q5s�0��W�;?��l�s�wB!�������b\1��m��ρ�4�d�CH����XO4ܣ(ݟ%i�q��B���0��Q'���Hk}������~�;�'B���W�<��S�`������!�tv�8?rL���3�$�����{��r���2�&�t}o��.ϒ���>�=Y�0e0��Ƃ����=duC�(*.��G���UC�o��Nz5;N1v�xt�ԋPI�)�p�D���-�F�2��(V))��id�jt�orO&�h�$�Jy�.�G�5x�]w)���}�Y�)���B}]v�؉�fb��4d����V�E�'�'�NM�Lm7�=Sۉ�3�gp�� �U���t�ȸꪫ�j�*%��M���8��(#n�TZaJ�b� P�����FD*5�!"P�-CJ�{|Y�ʤ�`�����r�n�%���י�U�u-�6fH���L	����уAHo��x5!�B���-��#0��@��s `�t����;�6��?��v�x�+쐰)Ф(�B��=K

m�(P6!�UF_(e�Zx�{�@�jl'�^v�x˒��邏�Nw��>Yϧ=t����$ǖN����~��.���.�r����z�\�Rc���,�ǨkkVHu�{FF�=�\��}����7"$��t���#??���M��((*!$��ڵE��K{k�t]B�]���wu�	'H�J�T���H�z���js���5������ĶөNm7��,�d���a|3X5�y��EĞ��NF=�Z�qt��q�zC��l�W�BZ���G�R��*훟^��xc�\����G�h��=�w�#���>UUU��[�p8@�]�7_}--��J�ݎ;`�v� '7W�o�Dn�ֹ��#Rzhc�o46V��ǆdX�8��qY} z�&ڰNc�9"ma��.���2m�ؚc�=�w�����fn���%�Sjc�B��S�������*c�,X�*Y�r���z������6�#������� �.�BC�NB!�$��nr����m�n���Ak��-��;?�F)�J�{���9��+6f�D�詧�*%��~��� ��U�W�R�k&Jan���ːckV�B{�2��-��͕��~��1�Z�:��j���v�H�۵�X�����r9�����⚤��	��4��B�;I	���Ay������-�He0���*�H%�*���5�GSp��������xΜ97n���Zlٲ�؍�M����ه������v�v��ﯲ%�Es{�l�&�P�F�0��s������P��sń�:��ƈ����eXٶ\*�����;"���:�,��`�[Zm!+ZsY�<��T�R{Au�'�����ss�6yA^ă����CNB!��	�BI4o��0�y�;ש뀊��1���������u�:�ۛ����,cy�%O��x�8�s<�cPYY�����5Cb;�T�o��
�k��8��@������X�b%ּ��bG���p�Wbƌ1�Zs��Hj�ʚ�|�.�U�X�Zb8�}�X:�C���ҭN�P����k��R�.{C�;I	z�����b���`e*PV�m`*���J���Ms����F�cl���]�]M����փ�_~96l�W;zBd�貖Vi)(,@�6۠a�f�W�������O�z�&���uǆdX�8.���s��	=&�T�gk7V,[.-b] ރr����w��K/�!��ւV��UȲz>�ߢ��L��k/(�	�In)�3��R�v���BO�H`�HE!$��ݴ'r�(KB!$q��<��/�@_o�B�АC���v~�� /ݣY�k�R������E��?ۥ��qӧO�m��&�׭cj.�B��b)(,���F�75 7/��䣷��m�280����ۉm����u�]�)S�Ĵ>hu\<j�њ�_/������ImW������|Fv���nnn�j�y#�/�e��aC�-`%��-.T�5����/@� X
�J)X��ƕ�MeP
Wfo��4w(�*��M�b]�	��EOd����cB�������e�]��K��;��݃%_-��¢"4o���n;���-]F���i��9>&x��qKm7k�1Li��v�0�=|�����#4oڰ�$eee�ꪫ���Zq�����]ml4��R��U��v��@��\N�}����J��A�sB!�G�G�X��Ԗ�B!$Q:��bk�f�y��B4����c��=�=�����I�}j�A���)�rh�/�@�Sit���]�Us�ո]w�,�j�--- Į�tw㻯���K�Eiyj��P[_��lB�ːÁ5�V��u6���J��	�+;�#���?a�ĉa����E����KknW��C�P,�ڡ?+0�%�`��X.��v��azF:>��!�0�;|%)Ň+�0{�D86��ܮ�` ZiR�I���u�X�V�T��<���4���(�����p�B��Β%K@H2нu+���KiWV��m&�y�IRjS�Ck�𘥶�-�38U��4���E)aj_�f��!��d�n�V���x���^j�����`)}A��`�^Л�>r�?��X�r*��}%�x��B�mX��wB!�$�[\���GY_��g�1#��%hQY3�z�6�][s�Q��)�B��f�X������<O?zsk�4i��\q�����A����"dG,�|��U���Ԁ��Zdd��C���ڕ��޶��C�t�@,�*//�g�/�u�X���vm�0�P,�`,�v������N�E̵&s"�v3�$��%)ǫ-i8��}[:B���o[���\y���c��B�ʠ��'�*�փj��ԂM���UTTছn���_����$��:���O>Cye&66�q�fz���10��*�=n��n��ذnql��|��z�ƎV���NFF��T7�k1�����-m��"}a�zr�����S���z�vi�SJ�{VN�\W��B!�.���!�B��b�f5�c��=�.h1(K��[3���:���ʘi�w����1�����B�[�|��u��7��k���B��;,�Ų$�KL��Am�DT���|���!4~Q7\Ѷ\
�FSB���3g���/GAA���V�%��.�c`n�	�r[�k���c��vhhn7Jpr�=��[��E��I��y����<X����J��nx�O����4�X�Oe�o�I"��X��V�9z���+紛x�1�X
V��ŒX%�>��3 $ِīu�勏?���'5���	E%Ŋq�G��Je6N�=��qFc�����c��n��ݛh�z����X�zM�d�0m�4)����4,q�l�h0����򺜾�m+,�A?�]���i/('0i1h R	��BW?E*B!�b�Z�	!�b^ku��*�u���C���5��!������2�u)����%5�x�+**�7܀;��=�I&���޶LZ233QY=�k�Q]W��Z���#o��׮ê�X�r�����d���y睇��,[��=&�㭝�_Ԛ��B���cik��`,o(��klw��U�v��aA�x<�B�I.xuKR���n|�W��ۥp]A*�p��U��,V	dQ)M��}:��JNv����j�{�D�h��q�O�`_NN�ϟ�	&`��;!Ɋ2ٽ���M�k���q�����c��nuRc�}�&���Fj��?{LL�LmNOw։�����ظ1ed�1g�\p����K2�O�*��#��/LI[P�����e
��8e�ܮm-�Kp7I`P�/hD*�s[�к�׺�B��'߷�p�ٙ���#�k6mIr�2p繇c�m�a'����7����@�G]e�GG'}�l��!���<��b��ǴF(п߬f�4��������r0t�?�!�z�@]���=�Z^(��D�����/DYY��>����Dh�"�G,��?��k�뤄wa~'���0���9�Ծb�/X��dE\��{�8��c�^��j{f�en���]��6��ە�XnˡXz���ڡ���:uk��.����C�+,�K#�{I6hp')˲�NT�L���V]1*����m�4����܁�7�1
C�R����^�M��2����l���O<uuu��k���B������E��s��P�0�#���jT�}�V��0�GhX�:�;����o�T	7����[<߮��X�j��l�`�$]�k�y���SNAzzzL�'�s�K���\������j��G��On�����U"��e��n�d�����	!�ؓ�Vlĉ���^r��1�p���^ŏ+6���ń'.�5�Mi�y��0��'��+A�AfF:���8�gۃ�Y�ُ8�ƿ�bF>B�����K_"V#���v~V��KrW�jס������v{��k�ꚡ�h��U'�w�Phg��~:���q��ף��_>"ɋ�庇�ݮ���	���mvN!�����DJ;;=�ф�^s饗b�̙Q���K�Q=�c��+���._��bOm7KnW�إ��r����v����>Q;��sNI6hp')ͧ��8��C�jJ�zPF_��jS^�
aK��.��
V����Oq��*2���.�����*U�NBT4+y{���X�`���J������B_~��i����rm�D���kF[7����n5���o�	>$úű����n�\����p8ذf6�[�5+Wa� ��Fd�ꗿ���K�~� PE{\,����v�X5�M\P%2�ۇu�)��]���t��+���:K��2<�*>Q�p�B�	�^� �4����C�~�4���l.�۹v%+3g��6��3Es;!$)X�Չ��ZT-�s����4c����.���P3Ԇcy����n�S�w�ۃciI�:a(��QO<�����Ϣf�b�
���q����"(*)���jL��W&B��֮-�/�lڰ��6jkkq��bʔ)q�Z��N�v-�ڡ:�s?�uCM(V���q0�6K�jk��±��� �k�م�$'4�����a�T��΍~Qʤ��@u_��� h[z��i��e��PR�;�b�[ό�ڡ��nr�Q��<y2.\����
_�5m�٭[����>����QZV�ꉵ���AyU�d�Wb��n4������>Xk��,�M�a}�����ذ�׮�:7u���LHUU.��2L�:5*�پx���=&������v� ���D*���/Py�+e��^��P�kn�?'/o�.y<L�!�b��o���n��ogs�?�ً�4�B��o�:1�i"�|u7+FwM0X�л#���B@��?'��]�Ь�w��W3\�d	M�X~���())AgG�dx/���2�z����v��[�FJm'd���{H�6�|v�ZKs�q�P���P,m�мn�2�҆b�B����N�"B ��5��6��I��+U��$�E+�0�"��}���`B����h=x*}���Ms��X%����C3�kG�ūP��<����jjj�$��n�	���:�dTӱi��|����kJiy��Q3�cǍ�1Fj"w�1�p��a=s{��{���0��jl2���#	R"�}kg�n�
BR��w�]�D;�x
Tј#��h�M��ւ�@�1�����{o���T�P5f�i|�[��A'!�B�I�ȅ��<�ڌd�o.�+7nAuy1!$YX$��&U��cm�Z�aѰf���ѕ�U�۳;����L�J�Q'�em1�8����>�pz���n�[o�BF#BOl�o���Za��T��B��RVY���dG�΋���"k���~O�hgƌ�?>
�^4�g�:b��|.��]��9�P,m0�����t�nn����j�B��$^Bl���W=��9k%����*x��r"��\���5�q�}�u��X�ǟ���=R�)�BT(iV�H����J<�� $�G>���O?Gn^���0���UU(X|46��`հ��<4ý�qF��&ڰ>ڌ�=���q�zlX�}���}��� $U�5k.�袸Tf�!J�s����MaP-r�A��ւ��԰"}����R
Q��T��6�7�}#��B�>7�y���H�oq�[�bnx�m�t�)�\�B��yyYfO(B_owj�r�P�ߚ�D��Y�v�_p���9��Dc\��D��0�766⡇u�:!J�����SZ��7+;�+QQU��	�_�ZIN��X֬Cff&zuDBF3���8��q�YgI��v�Z����q�z��X?4�2�
��w~��c���f5�`����b�cYL\.�$4�⥽˅�	Q5���]Z���vT�����e��*��8�4�!XY9o��ą��~�;)��[nA__I%���}����,�WV����U(-/Hm��z�1�plH�u�c#5��=��� �1�c�Ftl؈�k֡����2�5��3ΐ�F֎��9kn����ܮMafn7N`��/�]N_p��a��E{A�6��V��	!�}��7N>x���>�a%�uv#�8�\����؋�~X�_�T�]"��d�1�����W�������.0���=�jñ���r�g!^�[����#���پX�q�Itk�Bk�7o���q뭷bpp������U�WH����PJu/KU�.DlJOw�T?ܸ�!
/!�@nn��u���^�*�C}��h���S�������"Ky_��XN���kvW�ӫ�۳�2�r1��$?4��`�!�Ѐ�ͭH3Ɠ�` V�&'2��Fw��.��`8�g�����'��ڂ�M�b]�q����c"�C�>��={�l�����C[�H��t`����"�Uƣ���W^(X5|Gj"7����#2�GjΏ�	=&x;!>�uut�c�&tlڄM�7b�����Ÿ��q�A|��.������v�X��Z�{k]�
L`P����)�0\�����k��R�S%��dg̘��S���C!	f�]�p�)�:�1��'$�9!z\��[җ "}��َq�!{�B���n��3��e�&w����f���3���LMHr=�J�gar��e�/�j���lΜ9����j�k׮!��0�eyK��-�A�V��ld�XcKǁ�D��Z+u}&$թ����W^��w�=�B�}ў#Q�v�h��҆b����͂�ԡX�ڡ�.h��4����{�EF4�����9qDs:V��z	*b�S��%b��KRʖ��o�R"�ț���b ���c���.���eeߔ)Sp��wK-?��CB<�+�-���b��.�,az[Z��#5���jV7�8���!�{��a=���@Wg'6m��Q���7�	ѥ��W]uv�qǄ
Tf��������J�*����@�m1����HYp9-e�*��v������ ������=��w��ڎ�&`��d�wG�Bj+Jp��DzC�k؍��~��vb�s���O~�x���ੋ�^��t>;p���Ď�� �$/?lt���%=��:`�:a`��5C�����<4A��?����h��徽����w���Z,^���2���Lx���Eiy���-+��!�Dh�;:�)B�F��M�08���(�k��p�e�I&��Z�:.Z�vm��(K�*�����`,U=�gl^;42��eKa3~Z9BF��$D��G5U��s��T��R�J�������+�7Y(E*]�J�S)�x�e�z4��X	V��UUU��o�=��򗿀Ȗ�-�������,��t��Ri;N������î�bal��{�a�1��s�HU�ҹ]�G����� !$83f̐��E{d��can����ZjĩP�����~mr{0S��1���Moţ7V�9l��{B!�_Z��;	�/}��:�����/:S�ƃ�6�Y#�G�� 7��^�����؅�]�!�=�p���Nt��>Y�ġM��l�\'ԯ%��k���>��B����]{�x���2N�z�vκ�:�y睸�;��/��At�Uv�/��E��]$���,��} �9�]��E���M��N��c��y睇��<�55�v�k{ј#u�P���n���2�V%�����b9��|�Js;]��N�B�yey6�.BOw�D�Ȣ�^��g�˻\���ъU�M��f3�{��	��OolNN�9����㦛nB__!�8X�r������zM�e��U<��8����=ѩ�FccaBOVc��=�-]]����eC�0kBB#=='�t�͛�����Tf�%^��ܮ0�+D+���<�!P�2Kn7j/(��>arW,���eO��øC!$:4M(�3W����|�[�?�T����1���&r�ɿ���	A�}�t5n��� �BF;���qԤ	��X�>���fx��ݟ[�9����><����5�"\�{2���!�FͰ��@JF�f�m$��� Ӄ	�"�f�vm����e�}���R]���XZ�R�1��L����������)���#:��J�%���.��9s���h��b�Ϯu�`�ve��j(�Y0�6�ݿ�
bb7^�˪��R~��>hp'Ā'�A�8�S8 ���P�KS�������,UG���
c�,P���9!�����E��hr��>�v�a����5�\���vB�#^�6�� -J���%A�d�X��YJJP4�Y��vӖ��~wk�vC[�ű�2�'��]�����{�G��:r۳e+�n���(PTT��.���կ�A�*P���]~U0�kZ���0lA�
������ �2c"ڻ� �2�ر�/�p
�\��o��9�r2�ĥs��@��6�C�:�w����x�6IلBH�y�5�3q,��v�
--�k�i�z�<�}A�?k���Z��/�������j&�h���_��ט8q"���:�]��s���i�Fi������,E%|vv6��D���oDOw7�:;%#��)2���𨨨��W^�}��Ǵ��ݶK0sD�����ܮJm�1��c�c���=�C�3��v��XP2/��LF'��&Ą�=.��[�F,W��C� �X�6���Ղ�b.e"����6-M6��s�E+y�d�����'oO�:w�}�dr���/A����^iY�J�ʼ��P�
E�C

QP\(����&x�8Sۭ�C�{�v�Hi
==�[af�����7�������&\u�U�i��l%P��øP��򺮹ݻmM��7��t�,P)�����r��	!d43��/�x*���)���鹪���Km)���~J
rq��g��2����t�BI���7�a���dٴ@���^��$w�~�����q�F.����R�����ќ��|��gt>y{��ƽ��+��,YBHh]U$v�EIfV��I���zaq1

@�|%��[��Xb]d�I���~�	�»t��W���.�^(cen�GQ������B���:�X.ej�y�0�۳�v�����|Nq3���Nhp'$?lt���%=�*Jm`N����|��/Zi�ӛ_Nd��vЛ� ��!~�E-Zɷ�`r6� ��������]w݅�z�=�X\L����[��X��_�
�'h!7/y#�"�!g��]n��������L��}}�"��==ҿ����[f̘��/��������a������]O�ro-^{As�rqh��J밨�!�$#"�z�M�y�
�Uc����w����Z��$��o��a_Z�q�>�Qz�#��Y?�e��A�=��7x���BI5�����
�3�=�X�j��f��_3LS��60r��8&�V"b	�����h���U3��)�w�y'���?�7� !$r�iO��.���-d�����/�-��f��ė���vw�{d������&��E-�9s�����/�M%��>;��ܮ�'Z��ܝ��v�N��J�зx��c�����Jt�3��^hp'���t�Цzu.W�K�~#|��P�o��`�fl���7�+��������Oo�H%>�s�����oFg'Ӫ���P6��[��S�}
û0���`�V��fdf�9�Dvn�s�G��s���TJmY088���~i]�O��}���^���vB�A���֩����N;YYY�5���/��v�5���]��`��n����&��c�{�b"V���s��[��-!�{�v���sמ���c-#���{űx{qn}�}|��*Da����_�}v�έ}�����G߃�NƤ��].}h!��Te�f'J��c�`+���*k��BE�PB�ˋ�-Yc�e������J������'R��=�mr�Ƹx�(����p�u�a�w��@�>��Atl˦�}�Y�RmP,��y��37/ϳ^�/ൺ11F�Ɖ�܉[����W
����ꮄ���7�v���裏�y�d��vh�q��9xoC0�{;Ak�=+��5À`,�SSC�	Ͳ�%�^�Q�U[�@�h�wB,�j�s���ױF��e*�Vz�)��g+!N�$2$���q�h�Yfs��+��3g����_=����]B����,X�OCMZ�H{��͑��"R<K�d*��ʔZ ���v�ȭxM��&�1H�H�AE��.}�Y�*#��Q���!鹉u�����W�ş}A�:!I��s�E��?�y��P�&�x���B�B�@e�^Pafwi��J�IW��i/�_T���sC�r!���b}��/x�⣱�v�����k���w�F��؊����}'����A�Fާ�F>�de�?��{��F>�T�b���J����.�6v���.���翣��B!$��z�J���`\�Z/�����a���W@�PO���&�a���4���]�#i!����-Z9o4��OolFF�Ν���f��r�JB⇨�uun�=�����˗j��6(��R�07٢F��#m���ъР�җ� ,����R��>)(�uEB�ŤI�p饗bʔ)��&���1��8��]Q?�N8���~0�q�g=�z�P,����,����~F��!1���8���]�+-Z�'V�o4�}kҢ7�v[W�&�`s�aV�D��~��q�}�a��x�@I�8#�p�8cFa���"BF�3��#�+�ۥU!�9�oҪ͉��[!�mq��c�f8��RA���a�}��%�\������Nњ'�sDz�`�vY�����[k�����ւ���ZAʡ�^PY�Z_�A'_�	!d4�~s���	\u�/qƬ=�JflS[.-�d�5���6����p�AR����;���Vl!�B���\�=i"�V�X�3��y����ϊ�fݟ�Z��5�[q��8F���4��]�����n�/�j������}�������3��}B��t{{z�%77�g�#=#C��yB������Δñ���R ���c�Z�t��M��Y^<N��%���+�-��"K�';Ep�'KQ����)��}}} �$��bƌR0Vyy��ꁱؗps�X��
��v��v��v��}�5[����%�7�:��T�X�bz�D��b�剐��˝�WV���b��l����Y���X%�T~�*����.��&�{4�	�[XX��.��'O�-������ �!�yj�x}���!��!��D��9�#	���3Ϊ�= ���*P��u�yr�YCff>���~�T�2�y���7����p�y��� vd�����m����@I uX�ُ �B���[ܘ�4}�k��Bx����a�qP����0�~��uQ#T���55C�^(��&w�]�F���ت�*�z�x���q���K�!$y�%�b�A�_����7_}mx�X�V��B�����78�䓥����26��A�sDfnG@�PU7T�CKn���S�=uC]�u:?�M��K�DBR�		�'�ֆ�?nHj�$�JJ�JO�ҊW��Ei���ʠw3��d�O���.Hf���|�̣7V,�g�Fcc#�������B!$���R���P�LV��l����:�j��X���خ'L9t�)���?�j�jK��<!�؛~���A���#���u�o~��.�6w����B!d�#L�/�e����г�S�O*�i��Z�j��z�z|�=�Lir�Ɗ����_h���
e��"����O�v�m�믿�֭!��s��,B�����_,u~���ݶS]1����ncs�\7��jð̌�RJ����21��u}XF�?�KJ�b+�$��o<!a��_�T`��U��R�R
VZ�J�R���&bbmr�:.Z�������X�G�)�"���;��{�-B����G���L⹋o����f$�Km��=m���{��}�'��ً��,('�T�������߼�;���Ĺ���0_o�N��]\7̟?_��\"�졌����9��#1�%/��*��]��*��v=�J���sn�mď��@!dt�j�q����1�p�Ȓ>&1א2Α����~w=�!��B!$�^YU�Y������ӌ�?k���ݟ�8wh,و0���
�Fݟ������q�d���x���?�	�/���Bh�@�;��n�Ν����5��G�!$�T�����g��$�D�މ������V�s�=q�e�a����b_2����XúF�p�>��u�y�Ex}U>��mIjA�;!a�b��ٵh�2�DO�� ^��E*�`�qh��.&�h���>A�c��eeeR���/���o����P�ݎ7�:nn.#b�lǘ��.>�����@B�/~/�sO��]����l6u$(A����|NN��X�H�ss�5�/-,�������A��&+�]�6{�8�쳥ߕh	R�k�}�6��/ȷ����ݥ����Q�-u*��2XҀ/���N!��k؍[������?������C������M�ZB!���㝍c1}���<��ݟ�5C�Ρ\I�ޤ)��v��Z;4���a�7��k� Zckjj�`�<��cx��'uCIm�M��5���D�_6��g���;M��"e��e�y"�ŹU�N��]��\��¯����x�s�?�x�v�i�Aj�0��2֎�A+���06�{������j��QZ��0,E�g�w;;;�m�^G����$
�	���68�[݈��6�E����)S�*M9��1}�J�� �b���"�w���<�#�����o�w�}B!����*���X�Ad�n�6����4������t�,�]�;t*������[)PBH*��+1��p���9�!'+>�m��>���x��/0�JL B!��d��o_eUbJ�*_��\/��Ú�����Q��J����^3�+�`�͛�����rV�^�;V��!���Y*Q�O�sO��Δ�?{�7)봉 �=�k~"��E8S��'��NxG������,��uuu��������P�&�>he����$�]�خ���h��\N]��Q�P^���1i�z`<6�&.X��DB�;!���!��P���eҶO�J�Or74���	������`&w�خ]��`lA4��k����;����~�BIM�u�hK|����v�
Tf�b9.�v3c�O�2I`0La�Kn&��%�t�oI\�B!�g���mϼ��}��LE��q1=ߏ����-A�@b
}�B!���.
*jQ���ݟ5چ�n(��69��O^�����m^�W�0��+����ӦMCss3n��V���{���BI=���̙3q����"f��P�M�:��9�)������:>�t}�����!���X�ވe����.4��Y����1�Ѯ��dCS���4���U�@%t
WJ�� �g�B�D�H,�vAA�ϟ�]v�w�y'z{{A!���A$!�|��8��ӣ�V0�c�/�v+���6��jH#L��e�J�ܮIa([�Z�A!�:���?!�BI.D�������k����oB�'�!�w���c���5C9�R�x����.HthV4�=�h;a�)���g��]w�B!��&���8��3q�	'HI�^;��h�ۣ��Y��vq(C��u��M��J��IjC�;!Q��7�4O@_�i[����1��ݕU`���خ$��_q�L�;
Vf��h_$c��%�<�l����z|�� �B��gҤI��K�/�E"@i�)^y���=����͠˰��X��vEC~Q1^Y���!�B!���瓕C��� w�2i;�[/T�e�A�P���ݻ���]`^3t{M�z�����ܵ��ء��X+�fdd`�ܹ�~��4����BI�5���^�w�1ej��#��ve�0h0VaX���55D�XJ��2��	����(��t�T��΍>�J�ʠ$�h�_3V���W�h=�ݎ�`ξPK(�h�Z=Vޮ�����#����.L!�2����g�ƹ瞋�c��M�
��d�onW�/�	T	^�J�ܞ���7׏ŀS�EVBH��ï��WaM�V؁�vn�!{oB!�B���_mØ=i"��}z�Y��s�A�PQ*���]M���ĺ���F�S�L��wߍ�n����*!�2���G}4�9��Z3{,����nX;t���ܕ���H/��E-�"����(�r��m98��=]��}�P%��=����j;`��q��Qb���+тU4�	�Ġ�����Yg��=��7�|3�.]
B!��*++q���c�̙���h��#�ˮ��	T���0-s���hjWTF��R�ҊTY#ׅl.CW?E*B"e��K"��U��O���>���6!�̙>�=����\� �B!��^Z
�\�~����^(�{���}�xMVZ���[�&w��X3�fPVqq1�����X�`:;;A!���GEE�T;<蠃bZ;Lֺb�s�5C��a4����v���ٚ�ݡ��.��-�����wB���0�r{�q��{�_����	+��W,Q�\�B�`�� �b���B�'�y�n��nx������駟��!���L�>]�&N�U�v;Y*�}�2�k����M�VZ��4"UzF�����NB"gI������㯧�(��>']�7|��
$����=m&�8P�zp�}��B!�2zx�5s�ƣ�s��ܮ0����X(T`T3L�������]��5C�c�r�a�a��ɸ�����G��B!$y�6m�ϟ������
C96�u�X�ۥE���v����uC��^���\PZ��Z��OH2C�;!1`�	�km1fV���G�/�+T)�X����*�ocf�G�S������c�:��c�mk�*,,���G��^��[�r�JB!$���˓:�s�1��Ȱ� ���3��}�JqJ�O+LE��ndl�jlצ/�jd���q�`Ֆ!B���O�+���K
r�ܵ'��;^�+�Ǖ>&:�`�v��c�������7�kA!�B=S�Km����R�vuxJ&5Cy[�n�ً4hǇ���j���c�ӊ���|�7����a��X�������^����B!�$/999�7o�Ν;*j�v�#�����I�0Ts������
Z7T���v��_R�۲��9��wBb��A7��4�Ǻ�P�LK�dT7�"�,�!-��[�*^�����V�w�����m���.���kLf �B���w�]t���#�Bݎձv��ܮL_���]ܺBk)��t��SjK�C�&��	��L�Y��x`��{0���U��8�������`8��vB!�BF7���++�pX�}[��w�ݍ�v�Pt��j���]6��ռf(�21����a,��233� ��~�M7��o�!�B���v�MJm�v�mm[;L��b��v���$��d�}��ڡCSK,(��F>/8��#D�Đ��a|�^���y�,�7Y��w;�E�V���pe�� ��#������X+ǆ;��]VV�k����n��6ttt�B!�E��;�8)}A�0�E���X;�S����|��~k�H���FwS�J�4�b�M����j��	�%�L�"Q����BmE	������q����/���w�3Cs;!�B!��������م����0�#-GM����]��#�� �k���j���~{<��x���裏J�!�B쏨��8��3�^;�C�0�������bn׆c�kn���i�s���ݡ4�k�?���5Et��Ę����6�;�Y!�aIh��>㻩@�<"z�L�i�Ie0�L�
g_�Ɔ3W�m�|���i��p��7��?!�B��;�/�S�L���=�m;Tf�B�<�06�{����V��C���v�oh�`f�֦��,N��4��,H�����/�K
��{^��]�X�矾�8L�)3Cs;!�B!�E������\����4�wS]%`��j���&w1Ә &w�z��#��ŲF���8�!�G�4���B!ľ�/����ԩS��Vʱv٧W/�ܮ�!Z7�;+���`,Q;����[�Ǣ�As;!F��NHh�4���ZԻ���a/V�H�0��&�����oe"�L�`�}���2�A�]SS�;�o����N��B!6!++KJm?�3���7*�P�&B��M_���e�{l��C�"�6�AޖƔ4��e4�O��]����c���SP_5KWm��g�*����ڇ9W>�!�B!$u��v�+��T�Hj�!!j�����Տh�1ɺ��13�ۥfm�z�k����v��<���<��s��E!�� R��Ν����7(((`�0����~��e���ˊ��}H�خ���&�k�۳���QW9�\ �C�;!q�N�V7����s��:-- W!�bUzz��T$�`ev>�}��g�H�3220k�,L�<Y2���� �BH��y������첋�Z��H沫xejn"R�-A*�K�خ4�MmW
U^�*��o�R�"$��Ի#�n̟;�p��;�IK���ڇ�hn'IBq~n��,�+ʕ���߉z�B!��TCt�:c�f���Y�ñ�V�UIT־$s�%����)w~�l��n�brW>�x��Ý�h����\r	���~��X�t)!��x����?�{ｷ�m�z$s٩vhnn��:?���±�en7Km׮�I�%�㱮�	B�94�G�\=��k1�w�Ȗ��n0�g��j�{@���T��+�9ceV���e��Xm�����nÿ��/)�}Æ �BH������ܨ
J�n���x�W���ւZ����n&R��۝f� �J���P�7�d���	I$���=����/��}�O��v~�#��(/��Lm� mO�҈Ң<\p�+ �����z��uk���z9���bD�f'�+jј�L�$�:���:nD���]�UuC�P����a���ѬZ�?Z��k���4�|���$}�B!�G���t�I8����l;Y��f���v��a@�P'+Z�v���]el�C�4�Cq�?f�i��Ųͼ�#�
4�g>]������1�K�V��so�T�(	V�ڧ|N�������x�t�A�2e
,X ����@!���"�E���?;찃nA�.T4粋@e����nfl7��(�7�;u�z�vS��'T9�UV��[x�F���ɝ�v�l��f���2�����~sHj1fL�&��uM�3]x��)eI˚�=�¼l��Ǣbl!Č�7!}|��$-A �$a�
���$מ|5Ñ���
�Rv~V��S�5�h�#�&:�;}�t)���~ !�B�ǎ;�(�EQ`W�z$�ڥ���on�3��r����C&�v�C����%.�[�&�in'�*4�� >]���'6���u�M�k���n�{��d���9�y"�7s+���WUU�n�A���N��B!1"??��vN8�)�!��T���(P	��:�-�۵b��0���
�ܮ�^p�6��/.���;!L�'.?逸���v����$���љ�B+��U�c�%�b��@l�0�?}�q82A��Yx��ˤjB���vc�P�l����C���m�������Ё5C��D'�T�Z1�Gc[��z�!<���200 B!������c��g�a�����XϺ�|�cjn�t{V�����B���v��}(Hr����jk���1��n�梟b
�$�ڝ���&�nmS�K�ұ��D��L5����cx�5�<VE�p�鍵��$��b9���%����ƫ���:�B!���~����Css���h�b5֚@%�7���h�ܮ5���*M��+4s�R�����6��/.B��X��G�m<M�4��ddBY�*K@R����j{�����_/?G\�8z Į�+��?�?�^��X���q;oq~���8�m!$�Y7�1�0ah���bR+�خ�y����T�B�Ь�>�=�v^^~���Jz�m�݆o���B�.�=W��ϟ?;�3k�qاgnW�hn7����B�"2��u|����]X�� }��4��@�mwbFCе,`_D�n(4����z��4��x�O�%3�zY�J3^b�Oz�a��zl4�e��|����kp�Aa��駟@!���)--řg��#�<R��_"ŨH�cul<�P[��Q����>��us�J����ʪ�<��ؚx��in'��4g�$KZ�������~1�p̔��x��_c�Oah争�RR��g�>'��>��򘟯j\���ɍU ��p�z���(�o�/���ڵHV���]><X��^��\3�[Z{��v�	��?�q)ͽ���B����"��HnO�����d1��5��p,X�ۍ��ۅ�]�v�1�7b1�턄�$����p`c#�ٛ�n"R���Y����S,	VдT$3�Ee"C�+�cO�(��`���>�:u*�y�<������!�B�#�ifϞ-��+++��(�Ĭ���MZ�[[�d��А3ts�7�!�l<�o����d@��ǌIì�m�s���y?����$�nC�{��'��!{o���L�1��܀��������HH���i|Q^6�~���.�Z�X1u���c0����1'!D�竇�gu���I�[g͌�t�Nc��f�u���F(F&��5�P�srr$}sƌR����B	��*�S��ߡ�����C;�
C��ݳ�nh���Z0�lj���1��܊y7�7`���6  ��IDATJ��		�	�o�9q`c�yY��Mn���/���(���p�*X)�aUL��(e��v��Ǔ���SO=ӦMÝwމ�>��B	ΤI�$q��?���E&�����*n%N�
?}A��hrWR.���%s{i^l�
�RB�}X�܇�B	dJ�x��dmG7���ǘ?w��9�'�}�f��Ի $^���p�uO�ֳ���BK�df�K�g�#.y�u�������������X���޴�?�6!Dar߻�c�D��a:֊�*��Rw�����5C��i��%�fI�/�5�h_�)677�;��;�#�W�ZB!�X���g�q;�0_�h�
��v��rl4���E�kP7ԫj��c��C2��[o�pHeno�'4�4�b�js�WM�pt�nr���{Py�B�
K��)yd�B� �*.ES�J���HD-����&,X� �����ΰa�	!�=���p�	'��OFnnn�bS���`|�T�
7}!���#VI��+�@e��n`n/(����p��N!d ޶wj�I]D��c����b�q8f6m��#�}B��[_-����õ���3�X>��;7ཻ���}��]���A�:18�OR��;����d!#ã�]�(?Y#ۓ�����8?'�ǿ�eN�����!���j'~>�[[U�[�*�����_��������҇W3��q=Z5?���Hk�b������>������E!�c���q�QGa޼y())a�0
cC�*���Fv��ݻn�������B����wy]��Z؈OV��NH���N��X�:�Y�pl
4��IKzFt�[!PI�[�8k:�P^$�Ņ*�]$�h�B'n_"�|�|����Mʊ	>��V���>��C��^{�{��k��&]�B!�����q�9�H_���9�%@E2W,�+S�
��J�����skfpw5��cn��J�КIs;!��QC]�X�e��.'n��wp���t�u�,����� $^l����z	o/n�mgj�5+#}�����$�����<��	!���݉iuM��V�ܭ���[���ļV��SZ���x��Q���=ܹ�n;�r�h�q��a��������o�?��[_&�BR��N;I��=���w�vL$�ўst����c9M�������_҈���?!рwBl�k-Ø%%�/�8c1B+Z��+!TɷR�;4��(�<I�O���k�m��/�W^^����Gq.\�����BH*SSS��O?=얂V��i;Vǆ;�����v=�ʸ�ఁ�]ahw�'0	UJA*0��/���vB!A�p�tdg�_��-/I���/w�4r}��h�r�sk�噎K9���~#�ɀc���$ux����ﶵx����c}%����e����k1!$�_�Č�F���w�5!M}0�y٭^q�ӽM���\�>Ǻf+#{4k�����5��SC�u�]�$���z
�<�z{{A!������v�Ν����QW+�n'�̮��3����R�͍����4aX.}s��~�W3T������D�WTIA^ku��m^�C+R�tS|���`�� '2x��y�!b[\�$��K*��VE-�c�L��{��-�c�=FъBHʑ�����>Z2��*bT4戗y=���!Pi�ĭQ[���a�J_�
����t�핒��9B!IDiQ�8�@��d�t�Ʈ^\��[���왇�"&��(s�o~���KBCnv&��㑰W<�O<��g �CۚNr�#���Cp܁Sa7��l���<ZVw�B����.L�oDږ6�1�X�z�[9�ʷ�-����� i��U3�EM�i�B#=�Sp��/�^}�UB!�Jzz::� �u�Y���N��a����)f�C�����v�`��n�N�+h(����Q҄win'$���N�M�g�0f6�����4�P+�?=���`��Ifٖ�ޡJb��>+���1�����f��/�9�h5{�l�ﾒ���g��.�!����~�퇳�>�m���mw�)���"PYI_0n-8���-]��А~{� s�V���/�Z��r��&�b'2������b�mk�:�r\θ�Y��؅)M�q܁�5�ۍ�N< �}�#Vo��:����~�g9n��,��d&�!I���9�}�͑�.BH$��܅i�M�71���z>m��������w�C2�ۨfI]/Qi�Ѫ)Z����W\q<�@<���X�d	!��TA�N�<Y��瞾��c̶�9�N۱:��<�ui`8��vhP7�3�w}4��&vC��Y(�^ ��V��-n�4�uhp'����m66 �����d-�|ӗo�+�j�J9��p�Lc𥹏,�ANfHK��1e"�Z�R>�h�R���!y��1eee�?>9�,X� _~�e�/HB!�Iss3�͛�3f��9db!FEc;
RᎵ$PE��hpv���AD*3s�Y{���	x�%��vBIB�L���]p�϶���4���- ����}�sI���de��?����z<��XҲ�=�E�z)�7����/���U�_���j�P�#L�:#�7n�,��B��ʺ�\3T��#15�h�c]#�G�����>�}����s��G��͛A!��fJKK�n&�s233cR���^;T��=�r�PYC��ܽ�C�]���X�Z�+�vh�e��Y��]؄�2JH,�����V���؈�nu*���^m��R�2�<�-����9���4�4i[�#0�A����(M�z�&�h��c!Z	v�a�w�}X�h��^�]��B�h 77W�N<�Di}4�Q�n��Xk���/��4��i/�W:/��������eG<GQ~�s-�ƂRϟKJ�t�&�����f��NGq~N��->�<��q�����~BH��d���n���e����!�A�
���V��W<�B�N�\�j��ܢf<��>5C���QS4#:@w�q�9s��������B!����̚5���oQYYV�ʘdގ�X�$�-_�PZ�=!����F&wW`�˿m�ܮ��,��Z؀�V��NH�����$��v�dr��n�nsI�ֻW7���V�U���P%3xE+��HwW]̈T �/���}E�dH^G�J�G����x�	<��3���!�������?��v����&N�s�]�H��*P	�#������ghw�TA*=�ʻ�SV����BI���q᱿��غ�o~��؅��M�A�|��J���5��C�|�����9t/�t�n(/ɏ��C.������ŏ��KB�%��vb���/��
xA2�u��B�;@�	�3������4w��X#���h�>�7F� }��K�/^̀B!��)S�ଳ��ԩS��x���1G��
���@� s�b1Jm�^7�1����������m�U�#����NHL����$A�ܧ�5!ߛ� V)D#��s�VhVn�v�/R��*�1I!RAn;�Hpcx�G���i��M,E�pE�P�H��>�p��S\\�s�=�gϖ�^y��"�BIv�m7)uA�
���l�]ŭh
TJ��5��/L	�H)X�)�P�Jb��`(R9�SZ�in'���g��.�Ӹ���AIAnHǮٴg��<z �.\��h�.��Ղxx�#�ɘ�HQ���w��BF��rb��zT,Ð�O�kfD�o|uBU����@s�R��#5�H�|��&´NQo�N;�x ���*z�!�^��BH2��Ѐ3�8t���h����u��.�B��*�jr�P�~hT7ԫw}���v|V��j�rJ��~(n�n�f5`�j��	�54��D��}j�P���i=(��b�Y��R�
8�/V�}ij}������E+9�Ay>Y�2�����F[�B(�U]]���Jv�ax�G�t�h����X�8NN�Z+�D۫D!R�E��D�ȟ��s��>�?�g���.H��^�[<�D��'���D���}����.ĩN8�P�����1v5��{l$U4��"���]���/([��ܲ:��Bs;!ɀxI:��=���
t��し?�Ʈ^ؙ}v��#��$��>�޿��w� �E$;��ۅ d4�����=��+A0r8����#A�!�W�\��.�1��L�/$��@k���U�T$����C�Z[3��ӭ�i�~�0���h��beZ�U�v[�9c�<��x��'���B!$(,,����O<���q3��sL*��A±t��w���p,�Sܧ���'Z���4���n�0�f5b�Z��	�4��d|�r��6����w�_o��֭	Vj�J��{.$�b�����a0mME�4��D�`�|���B���m��3��1����.���R:�ʕ+�bJ���M�D ��x��盨�gee%�܂D�����D�_�����^��s��߼x�~��|s<1��x<���RI��3g���X�SV�$Z�J�\���*�G�֤��/(�*�"���@edr�(��[@In�7'��o���w�}Y��̎%9���_a��ɐ_R�0�����r)H�Ѻ��7n�[��ɍU ����u�7�kA!�����C�j@�s����EY7���U��݊���f���*g�X3�GGҫ��i�Q3�R�-AXVj�� xꩧ����L�-���+jW�$�痃�䰚x��?{�3?�D���'����Z<w��E<���{A�~����u;���ӭ�wF�T��?�C9'�t���,����G�/s$c�P��Hh�����6�{n����Pp�{��ݻ.X�Ո��NHܠ���$D��w߄	C�U�ҍbݳjlt�]D�/VYi=��If�"8Q� ;D+�,\)��^��+J�A�Jt��1Vƈ��������^���7oF$����d"H��X�|ip�/�evM��^~�I�}"����a*~�@	����>��g/��"=H�,//��8eeL�ŧXoG��`���=4�J-N	ûn��N{AS��������ڒ��:;7�W���yٸ��_a��-�������p�/&���L����)�u��}�#����2|x�� �B!��uC��G��ro��[U+T�b���
��|G�w����Y�P�'��=�v1:>5C�eY}<��a���Ə��.��f����ߏ�?�8j�����v]K��e����)�$U�"�Yև��g�= �ά�w�&K#�F9L� !� Eƀ ��c��:,go���y��ߵ�������%$`�D"#,��Q�a$MN=�߼��vWUߪ�U]�]=s��ݷ�	i��3���|����y�ݞ�����y�3���gϐ���>������_,������Ax|:sƲw�tΘG�b1�#4y�#��nޡ�34�cY���;>�y�v�v~ΟG[im@�����; 
ou20u.5%v$+y�A�"�X�Tҝ�m��9)R�����u�,�m��73�w)Zeb�xNX���)̦� (AJg	�-[F�\r	��������^   cٺp�m�QSS�˕8�3'j�V.�e��!P�50��w��v�H�s�&4ӳ���C"  ���K\��'��|Lrc�u�vSTش��:{���     ��~� ��ϡ��v	�C`	�'�&Gf��ͻ?'���=y����A����y]x�a�`����Us.\(v�~���?��?hÆ   ��w�!��}��������w�;�xoi����^}C�b��w�����v>JJK��,z� �� ��9|  m����I�����ɭP� ������1yS!�'+�Pb�z0-TY�i�j�AtO#�*"�؊0w�����k����ٮq�4i}��n����>tO��   @��}�٢u�N��D~�E]�
��_�*mp�T�w}�*njl�cj�h_07/�ĩ�p�lo7T|���fzak�v�   0����I�vPT��o����_�B     �0hm��������V脡��%���td'���I��ŗg���I{�|}����u6��WO0�׺��5����Yg�E��v=�������v��E   @.ijj��~����}H�d��5��^�]��:����ڵ�����w|v�+v|��>�+��׻���vx� ��(p6�Q���tZ�>�7ni$+rnb0�d$�96��P%5�D�}�A	�ԸݭM�i�J^'W"T.�������|={�l��W�B�^{���x�	q�   	�9�S�8�x��y����Zwl,�߃Z�j]V�r��4�+�TT�D�T5��!P  �-��������"�    Phl;����t�����c��(n'�&��ٲ'��a%y� <C�.�#���ǌZaP�aО`<�0甕����_OW\q=���b�{�   &t��7Ӳe˨��"0_0�9Q�ú��;�� ��o���<CS1������v|������}
��w@�@��Q���!�M���ۨ��;%X%��av��!Zɛ�&��@��"��L
W��Ny���=����+�����R���wz����sM�st�͟?�����n��F��/~A�>��B�   �s���-��B�^z��g��8�gM�_;�˵@e�䶂CC���N������-%ʹ~v�  �{^۰���Koo#     Px���g�&�ES�Po��.A6���)�n��M����̕����9:�Q�UUU	�pɒ%��ϰ���   � ?~<�p����|�&L��w��n�{�����af!�|��o��cs{�;4z��r�ʚZzz�D:܋�O �	� �t���d����1V)�Jf7�&�*�,����0r��̐le0�K�DU�7!B�*2l=(E+qXW��������.�慠)]��N��~���v�Z��L���
   ~�3g��_s�5TZZ�wqJgN�Z�s��vkc;#�(�@��w�*0�jD�ri_�in磤��6΢�n  ������{;�o F�     �{��؞	t���j?dnq���v^��1lϐ�BR�M�!?����F�#�u�=�:�aÏ}�ct�W����/���   ������.]*v|�2e�oP5�+��Ϛ(z������z����_�{�v��q�o8��n	���]��k�O�G��Rw�  � ��#�CB��|V1u9l�SJ�J>U50XĪ���!-z��B���Zd3C�փ2�n�I�*�<�>�G)X?�lD"���l_�~|~��w��{ٍ�|�������{�9��OJ6l���   @&�u�������@5nܸ��t��:��c���N���!���d�}H��])R�)���Jz�s*���ւ   ���Z�yE���!��7ѥ�M     ���HЃ;�i���>|`���4�[��v�aJ)@��f^�������x�f��J����/H�/�{��v���ɓ鮻�%&����C��	   ��7����3g�1?���XT��^��*�
���C��v�b,�ops{��zzh[5�ǐy 
 ��(CV�j��R�j۟��V�
2���Sc�g��'�V����I�����dн(��`k�OZ�J�v���֚0��q����O/��"��g?�u��!�   ��1{�l�馛��k�����@�(�X!X������}����a7���ڕ������z�P=�F�  @nx�͍t�9Ǚƾ}�s�o��u��t��TY^�{o�j�@# ��8oQ3͙RGQb�C�f�V �0���RA�4O�����&w2��Dꂬ�3�w�Щ�]��m(V5�g�ce���Rϗ��u����0�����вe�D��w�����    '�/������[o���F1���w�Cw��z�hl���5�����lo��<�V���PT[ � �0
J��M�tM��n�m
��T%�Pe|�jeQ�L�r��$�M����:螺�H��i�A���U���pu�Ma�v�x���y���:��9�C�/���~�󟋠;   �_#�ΝK7�|�خ��l�Y��5�
Pn������@e#N�TZ��#�P,��j^�k_0	S���	u������?D   @���V�c��c���������HQ孍������+7PmU9m�w�n�?��vw0�9�q*M�PM;��-{Qԩ_E���{�W6l�� H>����'ŷcye�s�p �X|�sΦ2�z�,�;�CY�e���X�q7�0l'��ar�������E�]��q�b7�c9{�E�|�a>��r�!z��ͺ��&���{EPq���j�*4�  Ȁ��%K��-��B---b,߾`PsF�wh�����s�oh��5�C'��T��볭wh�۳�p{�,Z�ZL�� D���]�ZJ�7�۶'GD*�p�jb�he0�V	�h%稄��he�g44(�����71�д�w(���Vˏ]�ȁ�����f������;�<Z�f�򗿤�k�  ��	�o��F�=m.��\�S~�D��^P<3���sq�8�"LǍ�v{��lO70��TN��,P�Ll���WR�  �c�b�ﮠ{Z+��쥨���ʹ����մ�`;�	�n��t���.����{�8���7���u��S�`-��>@_��TWS!ƞ|�}��?�W�Г��b���3	  �:�Y������H�m��~��K�Р�94�{����ӵ�G�;4x�F���Xv���K�Я��տ+������P�j�������u�]G��կ��#   ��B.��b���F1��`�ε�~��wh�[�錾��;��u�۝��<ϩ��*Z��|��&Z�Z Qw F9��]��Ltds�&�(S�R�V��ɌS�h�67����i�J�I����U
s#CR�J�ܓcىPQ��%Z鼷�:�1>�>�l�����/ӏ�c��nC  �ZX��馛�ꫯ[�#خ�J�=�kxy�tNjw�┎@e�[��*_[*Ī��3iek)�  �7�KО�N*$�z�F?��L_���Th������T���������ڻ�(J�������7�]���诮]L���c�;���6   �Yݚ�����l�}CRܭ�!ix�:�?z�1�^�lpWy�EER�J�9cY_g�	F�S�:ǯ���8o�<�������鷿�-�X���  0����GߛP�=@��F�Wh}���˱����ή�z�X����/�-�R��|�&z�;VUp`����9���{���@f+CJp"��A�2��^Z����ײ����V�sqV�J�L���32��GΊ�وJ~B���^�/�k�9'�1>�:�,:��3E����^z�   �>�s��hٲeB�*---�`{Ps��:}&^�
��"N��)՘]��N�J��kn-�jl7�/�7��/ �    �b��zR��Ҭ�	4i|U���6NQ�7M�D`lû �  j��2Dg�n�����34�ۍ�!Q�6d|n
�+<Ñ+����*�X���<��3$ˎ�F���'�+O��5��	r��؜9s�_�"]������GA�  � ����[n_�(��~׍f��)Ԟ<���y����\|Cǀ�����%�����fzc�  �� �^���6SmA��Dj���<%@����S[�O+�w��aE\sD��&�p��z�~��ԫ"u3C�!� '?"QP�R�B�1t��O�=����裏&o   4�9���N�k����;�<�<*�v�X���A\#8��x�'���s7qJG�rk^H���*׭!w�n��fz�5F      ���go8�>q�  ��Wv��MtL�.�����к�gH��a"Q�k�g#�/,J��l��EZ��]���#�u�=h0bcc#}��_��n��~��ϰ���   �.jkki�ҥ�kƌbl4��:s��Z_;y��\��7�;?���*��Z�e���ȣ]���7䣤����E��BN	����; c���ґ�YtZ�~���5܍7qJ�:�$yc�z0}SSb�ҍd�~FJ�ۇojR�U����|�%�+y�ea��γ}m}��~�����ur=v�	'����Z�z5-_��zzz  @a������t�u��駟�2�������?A^+_��\�v
�[��T�J����ۍ"U`�B�b�U4��m�     0�Yz�B��_@   �y�@���f�i5���������#�x�5�=C�|�ݟ3�C�Gv}&C؝�B�%ړ�s��)f�����
cl֬Y�/|�>�я��;��$   �͔)S��o�����&MJ��`��u��;T�3�C�o�j�R���-�X�;>;�+*+�厩���! � � �1v����xZ;uwq��Ū��e��ܭaw�ΐ�TXE�l�g���� ��a��r�|�555�=��C7�|3=��Ct�����Ç	  @�)//�+������Z:��c�X6����B�G]�J�s�W����~�(NY����S����]C��mmW�Uee��nl6���      �v�m�J�v�U�qf��.���?���~�'���  @�Iz�S��iG���=p�34�cI_(��=��S�}���g����g��!:
�aT=�l�e;���@w�y��~�a��ر�   ���"�~�UWQUUUV�`�cA�mޡS�=y^�7t�݊���3��*�P{�gEȽ�v<=�"�E��Bw � G���Ȯ	t��R�:r�F�J���xe�S*�N)��T٭��f�V�I���i�A��nYEFK���������#X�R�]5�?�����b�
q�۷�   D�	&Q�n�:L.��|��s!Fe{k�]>f
T��q�0e��D)�9c�]%R%�)s��1�n'P�D*Ŗ�����*z�H��D�     ��NmU9���7PUE���/���y��   $a���i��q�uhr��7$����3���3�2����C�Zʱ�~�zh�&v�a.C����jkkEȝw}��'���w�y�   D��`�����˨��,R�v�X>��w(����*�����C��5}Cۀ�C1��� �Ll���WR_,N ��w �(��qz`K-m�I�m;m�t���|������	?;��,\��˸��5�.���f�$R�yUD��E�ǠE�\�XaΉ�X]]�q�t뭷�3�<C<� ���   �̜9S�Y��;��`�j,jV>-��faJ-R)�)�ւ:"�N�BR�ro_�����G��:zb�x��G#"      c���+�y�$�y�~�����   31�������Ӷ��3t
�KR���g�����Aw;�aw�_h��#��W?/�к��z�`��A�_��rQJ��������^˘   ���ŋ�ݞ�;�<*r�Z\H�v��F�wh*Ĳx�N��V����w}6��ߐ�Y�BU���;�p{U�lZ�ZBC�� ��@��1�P�H|�PK#ڪ����2%L�+kK�5�lq7^S��.�S����T�LR�"�6���D+�"��5�uL%2�r���%K�Х�^*�U�V��;ߠ  ���~:-]��.��@��-Dq�Ϛ0-'a*y^j��UN�v>�l�[
�k_��ZP!R�L�NnG�C�      ܶ��t��6�<H�ߏ   5�>�ZJW�k��6�gHd���8���-��7���z�V���g�hqWy���#�a���l�??����(�ڭa;�8����$�ׯ��+W�O<A}}}   ?TUU��_N�\s�hng����sN>����5���;T��nޡN1V,������n�n�a,6H����r��� � �M	:sv��n?��'��S�!�Zc��(X���N��aڂP�ߥY��7m����KA�Ma�ڝB�ټ��5��p%[�n��~�V�^M�ʘ   ���8����)��"����]��`�Μ\�Q��n�c�t�)�XR����3�4��{j_P�T|��~-oM�^      ����4��n��u^�@�>����7@   �y�5A��i���-40���<Ì��P<��X$�d!�9�.w�6����BU���3�B*�>Z<� �������ԧ>%B���oh���   7L�:U�q�u������X!�Uc��+��V{�f1n�u���q��^��?���]�q��;��ή�za
4(dp ^��c�4����;ykcp
��JK���%
��Ķ��vO�SE�-M��H�F^#H�)**�T��xcc#}�3���o�]��W�X!B�� @0444�UW]%�S��2w������U�Xe+LY���T"�5؞l_��T��*q�Q�2�T�D��k���VT   
�����Ʃ"l��{;	  �7�JK�??-U�s�����Oһ��   =����6S3�Hz��pWd|�η��l���ܭޡq��/d�*���'�n���D"rO�n{�WO.J�v?~�)S��[o�o���z�)���M���B  ���?\č��!VTT��Us�ձ���wh���<{�n��V1��o�۳�oh�K�JiSb6��}�  �� ��ҡ�t��6����Z�"�p���Y�R53$��m?(�*�-�t�!L�VA	LaP��r%<e�����n��f�馛��_��{LX,�  �n=��E�a
S^�FQ�ҙ�����I�J��)��v���8e����8e��l�)�p��H�Uk|.�y;��   
�������A�3&�����3��/   }n[r
-l��:��76�O�:  ���}�tx�L:}����I{~�9N�k�Y��靟e���oh�Sa��P�ݓX�B3~<à<E?��Y��:Q�2��lִ9t��믋b��~!  ��q���/�=�z�b�P}B�1x�f�P����!�Zۭ���?h����U�5��p=��D��� �  {;���މtUcu����lE+"�5f��i�A;�*%TY[��J���>��I�6ZR�
S�
S����uY�\�x�8>��O��O?M+W��;v   g&L�@K�,�q�'Ƽ�Mv�Q��$`}�0e0���m��*�����!�ւv�v-����^j�B�;n  P8����ޒ
�3��i˞C�z�  �GC]��=m�t��"��  @���Ct�w2]>������Nޡ�7�ls�b��w(���Gq<.�T9��7Lb���~<�|�ؽ�w���-�q>N;�4q�ٳ��x�	Z�j�B  ���3�Ȼ=�s�v�uQ����LQu�����C�b,�p{zh�2,7�06|���L�L��UM��C  � Ƞ?�����ʖ94pp��V���`e�KLAw���20f�*-V%��Fa+��z�D+�s�\�6�w���Κ5���/��n��z饗D�}͚5�&  @�c�9Fl!�����Z1�Ka���(�S:s������Eu�=S�r�V�)Ԯ�gn-��������^[WO���~��  j*�9S2Ư9�8�  @��	�����C=  �?]qz`s]�2�znOjM���k1i�0����[܍c�~!#�B5~<�0<E�9^��(����O�N��v�������W^y~!  8PZZJg�u���.���21�����Q��|y�V��8�W�e��y;�0�p{U�,Z�ZJC	��; @၀; @I"QD�[�>��B�G�؋O��͏b,� �s�`e�~�M�������)�ȩ�A"����:S!���&�bQ>�'��ݮ��l�{��ضm=�����Sww7 �X�ۮyA��~��b,�n<�"V��)?k�U�0e��[
f�U6��q��������F06"R��)�Hen�BԠ]�}D�z@Tq   
���U����$   ��������J   �g(QD�Z�.in�����mX]q������r#���\�%���B��;���.?^��:�zN��t�]cܸqt�E�c����/|�G���   �ĉE)MMMbl,���c�
�g{m��a�g�P�w��s�o��}�ۥ��RbR��'�^ &� yjs�N��Ds����xK���<4�,u��x�$�`E���lg�؉V2�.Ī�J-T�E���E�ms�2'�u~�������s�ҧ?�i���?N�>�,=��S��/���  0��υ��~饗
a���.5n7_w|4�X�d����B�,C���P�U����Z۝�\[��T�*R���,tQ=*   ���	������4i|��   w��XC   �����贙-4�k�3��z9�^a���K��n��_h���8l��{~.�5+|.�к1�9Qs���������|���Nz�'D1�믿.tO  k��R.���~�������?/׈�X���(x��1c1V����ש��v�B,�%���Ụ��	 0:A� �ʺ=1:2q}�z���P*��pã����JK3�d����`'Z��܇�;v/2������z�7�:�S�!���B��������E���;v���{z��h˖-�  �Δ)S�K.��8��!4y����KQ+�k8	S��N[
�(�P�s��lav�m���#���)o�77�   (d�j*m�-�;�֬�J   �cp�{�8�>  ��vRӤ���r/����>����>�C���'hW�%}C�?(��I0��d%���3$�5��������;������A�׽\�����.]*���Vv���~G{��!  ����3fВ%K��.?�#���g;�+�P5^a���F�ޡͮ�:�X:�X;>��~�r�gKН�9��o:m:�p; �� Zl;����lvuڟb��˛���2׹���d�����*PYǄXemf��������@U�U�!�0�|�ڽ�QAW:�gϦ;n��vZ�~������A  P���Wn[��+�.�ն�xԃ�(	XN�HR���{5'aJ�C�vBU��v��{EU��5�v�G�  @�3������Ʃ�    �ȳ�P�ګ���tPg����d������N~�[����Tv7�c�1�1r؝�,Y
Y���vS�m�ٮ�2Gw�Ϻl�7��:�����'>�	Z�f��
��y���#  -p���Σ�.���>�l�'2��f�>�~b.�����C9�����<�ۭ;@�c����S{k�p/�C F;� ���ӊ��te�l��,8��W� ��Y�<�I
T雰�p%�(5�N�b�0ejrigP7��U��]���u6k���y�\�97�q~<��q�]wѓO>)ī��zK�4 @���c,��/�X�-ps����t-��|�X����z�S�=}^ue��n��`��ĩt�=f��ۥX�p���J�l����!   FU�e��o�N      �z����j����znW������]����m��r,�]�=�/�mr7{�d)ʒב�e/4���{{}P����'G����z�~�a���,�� @�a��k��ɩq���/��;�C�B,Sk��7t�[��:����3i��R��k4 c� ����V��9���{������F�op4*���&*砻Q�RWv�r,�����vc3C�HeE%Z!b=G���՘����������Z�v������O�S�  �7����/��-Z$Ƃ
�5�`�j,J��k�Y��R"���$Ly����H��Ӑf�=%N)ĪXl�J��ҊM�qC�  0z()��1�㛧      ��P��V�]��L��[\u);���?4z��6�d�=��j�z�ZM�#�w+<5m�ks�cQ��|�^�r�>��'���_/�6�b,�<� i��شi�D�����Ɲք5�O���B��\#�:x��J���]�����w�
����l��=ao]3=ފR, �� |��5M�K'U�����͏!��'�nlp7
W���t�]�Π��Aw��3�U�v��@%���Gy��U�ʇ ��P��`�G���~��1��9s&�|�ʹl�2z�����_֖-[ ^ �F}}=�s�9"�~�g��B�Ϛl�%/׈�X��)�9VAʩyAi~��M�����TZ��ǘ!��=�n���5|�}Z[�<z�u����   �H���na�gM�ڪr���'      
�g�т�f:�tw�+C�r	�Km*���BØ�U����|B����0�r#hJ�S{����a���<���˧7�e��k�^�x��c��=��Co��&=��s���SGG�B @d��a�=ĳ�>[|-e��5��`|Pa����Q���X�R,��c���J?�l\��g��[	 0�@� ��-�c��g2]1��:H��(��q����Z%%z!w;�J�7~F�ʮ�A#O5�J��9�\�k���ݵ��裏���.��~�iq:t�t�{��Ӹ=f.�luuu�Ķq��Q��?s��(���F���|�ٳx¿�|mߙ��;������������O�o�*_a�׃/İ{P��䣝H�y���v��v�@5����@e��.���*Z�;�6�@  `t��7`{�����>��{�]     ��x�@��UM����Sw���F%�C�;?'�ڗ[�]b�	�x�~���&�>���\�e�Kyi�%��.���������;�T�=�����g��uz>��nz��W�g����z������ �.���"����̻�3Q��S�Z���;��z�r<��w(��Cc��T�e��<��3<C�)��'�s&ҁnx� �Ep dEw��\EW�̢����7G�J��~�C63��gW�b�*��t7�U���
T4r6�6w�5^��W>ǂ��͸�5���x���O�^~�ez���u��aG��^�����G��?����
l���@���5&_���������H}S�/��{�s,,����Z�?���Yg�E^xa�$����)*�|�q
���;4/$��n�v�p���=����IS�U�5���   @�t�8o��OO��H��j     �z�j[-]�\C�������n1V���*Ŋ��ܝB��]�����5׵��B�ϊ�ڝ�#$E��|�����P{�A� ���]�iMUU�(�������z͚5�7d�T�竜)�A�~�3�?�|�3���U����Οk�j1Vex|�N8A4�_|�Ţ��ɧ8�<�\��������X�;>�l<CyTO�In.��8�R �*� �fh�&���bZ<��&�lARS+C�x���7X�6w'���8���t�D���e���Tm�f�ʊ�+��8�m=ʂT>��l�u������#_�җh�ڵB�⦆ݻw  x���8��y%ۦ�s���0��X.,�%�e�T^[۝�)�p{����оP9y��T<|_�q   ��:�r��)�w������	     �B#'Z�ZD�47S���~�g��j<�*�A�r,�������^�v���3����:?c~�������:��p�>�!q�ݻ��{�9Q����;����)���D����a���;��r*��LA��ۛ��;��?{��>����$dS{CC���a�<�B��TF��?��;{�<G`��ҥX�ޡ�g����5���0�A� k����sia�^���$������p|���$b��4�����I��4��a'X���w�-�XP��(����
N�B��@�t�E(�-�]w�Eo���hk���@;w�$  ����^����nk��&hQ�������cVa�(X�ϻ4/$���*�慴Penmw�L��������k[���9� !  dä�U5��W�8��:�W�AX���Y�J      "��<D�4����"L��z��9nis����_�|m��|n*�2�m��G9�o�=L0j��h��O�N˖-������W_aw���3 �0�P��'�L�w��O�:U���#��&����B�{�}���&c�`��R���+<C�+����f�IooŎ�  � ����)�BKf�Pס�����A������,Z�O�f�3�-�w'�*����@2�>��n
���X�*3��t��1��~��;��~�ɟ�惷%\�n���ք� ����?O,^�8���P��5a�[A[Q��E(�,C�r:T[;;�S:�vlE�240TU��+�� * @�|��K����V>�v�?�=������8���dO[���8���v�*����t�gD���     �"���5���ɇ���H�+4iZ���ӥX��{�d�Wt����N^a��,��������_��l�u����9�^y��8|������A�= ]xw��;�Ǻ�:1�0��(�Uc�����=T���P�4�b���w����G��I������� �w @�t��i��
������l��,��U�=����.�IQ*y#�����Nb�Q�2�U�Fw�6�4a�V:׉�Xs��?.Z�H��smٲE�����khk `�_W�9���Ρ��N:)��'���ӹB��Y��u���A�.���J�R�S���N��T�v?���=C��<��:��b�  �����64\VZB?��5�PWC?Z�
勪�2��/^�nw����ᯩ��'�{w/u�7yB5��篥��%ű�	     (L�uѪ��tes���4k]
�0ᢁ��ܭ-�	�Prw
��С͝F��$��}�{�s�c�����xPk��'M�DW]u�8:;;EН��_y�:x�r- `l�;=s����N����Z1���������Y�K����\���s�c�����z��:�v�p��7Lۇ���Xv>��nϩs�AW?��D4��  Hp ���7�i�&:�t7��o�4�����%螾Y��G��C�NbU�1�>����^T�׋�h�� �5��sMMM���멽�]���x��h�޽� ETUU	1�SN���ٳS���ӝ��S�
K�ʅ�%q�\�t��	T���t�=)B9�Ucn߳Ml��C  A��@;]������V�X[�q������/��S�D�8���o��~�w���cf��yfm+}��W����::oQ]{�q���H_��<����#      
�X�hUk1-��L�z�S����_h�o)K�F��3wv
���B��Z���Q���6w�o�v�r�����_�ܰƃ^c=?~�x������Z�[o�Eo��(�z���0�������;<��Sš�ӳ����ڽ�G)خ˕�h�/�2<D]�0p��l�Z����Q<|_v���^iE)  � ���FM��#m�&v�f'�*�6W���������GnO���*�`e���n���hejN�Ƃ��x>��b^x�8>���Ѻu����_ֻ�+�� 
)H�y�"�Ώ�snk��/�*j"V���U���ۍ�Jv���bU��M������������;�Z� � ������k��;s�N�����]E����N�H�����2��v��o��os�1����|�N�?���Or���ϡ����H      2k��h��9t��6���P��R�~n��sFx+tO$��ݟ�~�])�|�� c}-�B�6w/^�D��F�-~aP^��<�Z�(��O}�S�m�6Z�v-���˴f���(�������>��o��3Π���>��:�+�p4�ݳ��S��m�g�`{Bx��p��wK���`���V�UYSK�v������ jp �N[O��o��+Z�i�m[��ʦ�����xOV#��F,}Cg���Tb��R��8�-f����읂��T��_�)(�*�k�\���������M-b���'?I������녀�s�N�z @~�mO:�$:�䓅0�`��@)��$X����`���5Ԯ�|T�ܩqA
SI�*�nn��SB���o-�
��s5�]U�яp;  \tB�W����>���u����4&���h�j�9O�m��!�>����O|�z�[�SYi��<�~��k��/�7m�{�      (dvw���:������2���XV��i�紦��W����X	C9����F��X�%B��0}�j���zr�`�B�^<�(��Aڭ���y~lllǵ�^K���"��ꫯ�cϞ=�
(��3��,wz�R,޽�x�i�۵�<��UO��D�0{����+���+4�=�T���z�LZ����� �A� ��"z���3����v0�M�6��6���4�`�lv����N!��V'��]�2�V�`D+�X����B��r-D��g�vڴit�e�����Ɔ?����/P{{; r��F9��cE���N���]�q���s٬3��x�D�0�)��$R)����TV�ʮy!S�J�S1�s�F�*����� PRI}#-oM��  p�����%��G���Y�5�#߼��������|��v4���Rey�����6�6�������]�8����~�՛�/��:C��      ¦?��K���f*��F���T���چ�-~aiJKK��l�:����Z��C�(}� ݥ���F)���ot��;������z��Z�^r�%��y���b7h>x7莎���o���Zb���X�w�)������F=خ˥w�
���ܼC�p��w��	:��v�_��B����! �� 9�]��{�lZ\�F]���6C��I�rmf�d;��Xelg�[�����G�ж �㪱 �\	Oa	Wٌ�Fu��Z����ؘnl�y뭷��7��wny��G��0�1Gu���?�xѴ0a��0)��A�R~��R��27jaw��$�D*�}�O��^�����TR���n-�$T95��ظ�2�V�H�[	  r��[�C�G�i�Ǿ}����ц��}��$�Χ�����n̏V�Bg;�.;��y�gM��߽����rq�      @����!j��H�*�QoOOJ��BU1�S�=c��%��~�gy���·�$+	?&�K���Q��	����͸���u��y~�?�8���z�����;"��~!7��+ w��0K����X�>��w�P�jf��J���;T�ٝ�C�b���;4������>bEe��J�A 聀;  ����v�ч�k�����U���VN�����[R�R�3X�4ދ�ܭ�u� Lb'V�q
�) u��ׇ5���ds��Z��������O�tg!K�{zz ��w�_[,X@'�x"-\��-ZDS�L1�ѹNX�s%Xy�VX�V�D�`���WW���0
U:���im��V�*B9�/8�c�T3����SC�{n �����I���}�r��o����� �_����]�� =�������q��-�7~�     0�t(F��hɬ�lۧU��S��\#}��a�����0����������?�ҬD�����w�=Ho�mn��:�ֹlϏ7Nj����[������+�П��g����{B� m9��E;;�b�z�TWW�:�?�v>��aB�Q�[ǒ��o����om7z��z�N;>�Q[?��QA](| x w @^JЪ���-4sh�h��ݭ���X��i3�3E+�6wsC�J��υ`���he�E+�^��^ǂ�r�>�qݏ'�s^��9o��m��{�8���>v�����oБ#G �	��ܮ��v�N9�jhhH�"Ю3'���ӹ(S^�FU�"�[
�*�p�}k{�,L�B��ւvq�V�y����&Z�iH܋ @��	���ہ����w��|��W�;ν���i۾���O�E      �:��|S]��L��[3�Es�
嘲��R����7�osOͱ��y�c��w	?U�?&d@^��q\5� {���B������4i]v�e�`<H6lHy�z����_: @
��͛��a�0<�(��a��a]#*c:ޡ|t��!v;���ώ��P{Vޡ�3��"�_��&Z�ʾ!�C �7p �7v�h[�L�`Jui������Ūx�/v���������U���t�J�݋��p����习��̩��?9��?8­�7n�w�}W�X;v쀈��'����������4G�Z�:U�*
!�(�S��,N97/�m+����.NŅ�}����A��
VUц�i�n+��{�� �0�R���77�Ǿ�[��A����?XM?���2�7��rj��F���� ��~   ����-C�2��U���n۠�]���X´t<���p��۷��s'�P�ڶ�����K���9�����1��~��;��:�����B��X�4ݹ �=C.� ��?hg�����C<�3����\'�9�����c<�>���;��B��s��=�y�	G�P�3b�,~�7�P����#��;|�o*�ߊ�v �?p ��C�|k-i��ءm��vyC6�XVVf+V%_������ܓ�U�A�*6�uC�P��h�$S���$Z���B��>��1��s^�5���\�D9r�޽{E�}ӦMb�µk׊�w���h����	nV�����:��ϟ/�k�q�������~<�"�~�]�j+R��m���F�Jݼ`mn7�T:�
�]k��
N�N��^N��  Q$
!w�ہ�����o�@_\v��qe%�󿽉.��Oh��C@.��'/��xǁ(p畧��s    ��M�b�����h�@=vfcY�2�`��?LXK�F|Ä�3T�b�}Cݐ;?:��<|��i$=D�G��̧����|��s����9��Yg�%���W���rA�cmݺ>!3�3f�@;{��%.Z�����Lst�����?��'�͘��wȸ�����q��[۝��=x��b,CȽf�tzt[�"� �� �H�H�c�q:~j3�+�E�}��m�f�k[�ʦ����`���n��vB�HXnr����c2+�/�t ^���8�����^G~�>}�t����c�"�Y,d�����5�+��*477�;�*��p�B����(���DA��&a��ܨ�Svw7�ʋ@�l��1�P�Y�r��乢�"��B���|�  D�|��n�|�7���&�ҳ:��ÿ��e����)��# ��o��p<��f������:z(_p���n������m��8   
��X�Vn,�s����m4�~��k�p*�2y��R����&=���Z}ô?ȸ����������%c�G!�����5t��e���ds͠��ͱ���q7h^��X��G�m�z��E�B���s!�1�C'�|2͝;Wڛ��R���<��e;'�P���\����Gu���g�ޡ����;��ͭ��v�����<D�w8�G�S'��8 @6 � ������i�dv/u�kl��)�*���]���(XI!J�s�tD+��&Ib��|�ڽL~E'/�����:�y�9~�q8���������l�B�7o�;v��u�����!f��!E(�X��@;?�P{]]]�\�k5o�V���̍�8e��bT�Y�2ۍ��@�C�k�K�Bu�xz����mC� P8�#�p;��G|��WS��z:�i��\����7��_�_�Y�����H��k���;^y���3���Aˆ���c� ޽�w_MW�c� �y��z�    P���=F�&̡3�SW��b���_��&d)�˧�܍���oh�
U��/t��9y��1ae"�3A�~^����E��нNkt��g��|6s����,�:�����`���;���*�BY���� D��������(�S����z��s���X5�0W>�j<�P>�O�v�v7��/��=��l��ޡN{�kk{�Dz�`�9� � "Gg������M�Tܱ����f��rÖ�ق��<1"Z鵹;ݽ�ܭm�#��X%1��j�V���:�s^�g3'�y��բ�	��m�6����w�߾}�8@Pȿ�3g���|p��[ZZ���B9�˵���*w���
��G��a��0%���mE*�Pe��┍0elc��<��\D�8 ��C�ܗ�#4i|�ɓol�ۿ�p;�FOߠ���'��N��q�A�sNh�o}�
��& �e(���|�A��.�>w�DZ����-_���mړ������~�77�Y��Α��w"x   �v�Ѫ��ty�x8�ͶKu8�-d�]���cx�����KPU�e�j��l8�X�i/1��{>`X���|�lר�yY���9v�sهY�h�8$��c�ΝbWhnzokk�� �5'NeX��3�+r��w)0�7�;/�/��Q�úF�>cvޡ������;�ʰ��v����C�_��;7y.�ܔ���p @p � �,On��I���� �tv�������F��N�2�2�#���9�n݂�)��[����d��3E*+A�VA�97�q����9?烜���e.�d;���0�mooA�]�v��w��k~�o|� ��f͚�
��s>i��ɦ��|��j^�
V�
�{/�`���^�����N�]'�Ώ�!s[�J�r���i+A�0ŏ|��V�H��  2����?�ӎ��{Ć?g�����ϩ�w��;Bw~����[����>�O��v��~� ���{C]5=�n��{9=��5�iڤZ���?L���A�   ���D��o9N��B�b;D���b,���Z�&ݓ~���ݝB�����ih-];�%&�j3��{e;��sA��fN6�x�]ٌ-aM��A.ǒ!�7m�D}}}@�������T���#��C~��GM�h���	�Y���_3��# ��lwkm7���7�v�ͥ�Z�ћ�  n � �4��h{�$��i��ṑ�N��7��F���Ħ�At7
TR���
W��+����t�=
A���1�e��9����|�s��e;�_�Oǟ|���0���!�����~!l�s~<p� ��c�{2a��3g͞=[ls��]��?01i�$-�@�}������y<��v�/q�I�򶥠�0�(PY�t��s[�ʰ�`m�4zrW%�C� 0:xo�q U�_���u߳����u]L�7綾��J d�NȽ���~�w�����Q��'�
�c9f�n�9y���ہ�	���_���̫�ӏ}�   ���m��IM�ζ���T�a�3LX=ô�!v��{�7��C��;@�#�j#���lƃ^�v��Z��A�Q��2���б�!�����#�����^ܳ5ܼ>o�<��i�ܹ�G��bMM�i�W1b�sƊ�`�jL��T�Ct;����3?�",{�Щ���)j۵���S�]Ut�7F  � "��P�l-��ͣ����'�u��
U���V�DR����A�d;����V��*^Y,w�trnX�A�	z���{���y��~�s�ٺ}!���:tHY|߷o�ٳG��y��#�^x����z!2qco������)S���ܶ�'��u]PAu/����Y���uM�E,�cA�S<]G����m+(��:�l������������n   �%��E:�e:]q��y����O]A|���� v ٣r/-)����4�~<}��?�1,>����on��U�sn*�Ǖ�U���(���  ��C=qZ���>��B�[i�����y�����d)�!����Y�R�b�&w�r�0{�D�;@����1*�`T��0��x�~����ӵTs�ί�����:JF8��^ {���޽;�C4��yx���o�7�?� ������`%�0����<�0���?�u>������!:b%��Ot��Y]�e�f�㳝whjl7z����Vx� �pA� P0��;H�6�MC�spW�H5�f�����-M�j���Πr�G��SU~��޷!�v,�a��Fu��Z?�u���<��~�ۭ)++��S�����z���t��Ajkk��9��Y���w�t��wd�iڴi��ֹ���;��Չ����?W��g��a͏J�=��A��Z�]>�����)��(J�ۇ�x�V�A	T�p{M�$z��x�s�    ��Ɍ�h��zq4N�D��^#<���Φ�4c����������ڄ������G�;'Аyqq]z�QTVZb;�w-��^��  ���S�c4kB#�9�u��,�Rx�v>��3Lq�!=�d)����n~��3T�����=ƨݳ�n6�OX�>o7Gw^�>�j>{M�����:���> {���ݻW��G.�b���=A~��w8��>"��`��"�y������y�0����+��Ϛ\��^�flO>�Ɯ�B'�P'��KU�%w}6z�N�v���� r	� ���/F���:kv5적�e�}�g�{��!�����1)J%���`�ngP�18�ݕBU©��y�5��m��k�^�ϵ������l��5�n����<����Ǐ���f�:�����]Z|�@<������9"��2$��d�L�Ϛ[�u��,6qX]���o�ǡu��5�x�l?����R�ҙ3������`��u��	Tn"U�@������H��J����8e#T�aG���bӐ0�    <k+iѼ��q*5�����@G�j���2�׼纳�S��0X����W�D`l���Կ<0|�8d��ΜsB�nnG�   ��l��ʎ	����۶�6�;5��=C���g�tO��N~�Sݭ�@�[2�a����{�l�u>��΅q^wN6����o��Ǫ����w��A��d����â��[4�Ỻ��	�߭��V��9�.K���ȏf�9����:�|a�/�@���\����G��h'���96>�f�]5��;��<�f��Ss;��E�i�fx� �܁�; � yi� M��AM��C��*KC�j�A��3� 9�B�jB{��-�n��B��qB&�Aw�k����ky=�e���~���ӽ���:��]�~ܸqB a��	���? ��w�X�������uww�G����k�:��|c����9��0:�` �F|��cT�F~]YY)>��dh]պn�~A~�a�Z��B�}�V�
�g
PjQJ>�Sv�J�rn^H
S*��CFN┛X�!NY������j�M��CB�}    @���b��=Wӵ���Ǖ�Љ-�)Nh�No��5�[p��g���x�r�n���n   ��}J"A��&��f:�b?�vw�c<C�b,'��tO�~�ݟ����/t���'�w������Y��u��չ��g3G5/��v��ָ�eo������'�eX���k.������9��x/�h��g͞����G���ȏ�{��<�����񱅱&�"��hy�N�vU������7Tc�J���T!w��m[ە��A����?�N�M�	�!  � � (X��i��J����J;��@���T��M��*^��dh-ns���:�U�@�
���)e;���݃���x�k���|6s���4�n������u�ð�,�� ��F��xX������/������M����O/�S��y�K�����y�?^kC:��s����5, �Z~�ya�7^���Q���WH�U���(۽�.X*'q�*R����[:	S��*q��|h(F�&ϥ՛�?Ʊ   |[�ݿ�2�p{�����;.�~�D��-�rG�    *�;�-��芦��{`��˩���3t�GJ0JD)���w6��N>�*�Ϊ��P��ݑbш՘�����l��s/k�:��|�s���^��~׸�ӽ�g:Y���8 /��dA?�k~Ώ|�\~d����c흃���a�{�Mx޺^���s��s\Iϐ��9B��X�Cz�\�%K�x�]���	
��
�Gr^ء�B��St
���vav��خ
�����_���Yz���X���1��<�Vo.���  @�A� P�<�%F�&̥3�PW�!�wK3�]��Ѹ��%i��*Z���V�*�vϾ�!-RY�a݃���������a�Q��:�i���u:�u���VX���d#@�AX�\�o.��|�)��t.�aS�q�`�v�✟��P�N�1���ܮl�c\y�(�K�6"�   ���	մ���PY�8��N�H[�"0��w��v`d�������T���c?  ��Ѫ�Et��y4�v%���EXr�D_���_(���tC�� �vhh���C!V����~�{ϵ_����=�����\'�yNs�Yc���5t��H���~�?���,̒�w���G>�H���",�\"˲�9�3ң���#9Yv�A~>x�_��~�k��a�ٽ�j�C��a{�z�v�o�s���D/�X1�o����������(m�u�� �� �Q���!Z�QC7M����6���h�r�n;h/Z�W���Z�6�w#|���N�=�k��o.��9�v}���z=��~�;����~��|�sE��l�YH�U���ۜ��=�v��W��M�2�q�l���L�J'�.�C��z�Lzb�8�@�   �B�ނ��q�0��W��v`徧�   `�=��Z>�.��O�v9�����_8����<Y����ٮ�]wh~��;�ɡ+M�Aw/ss�hw���z�A�����<�s��;�q[�{/��sm;d��s#z��Q���X�^��B��z}~���?̗��9�n|�!���zkn���Y��n��M��zb{9u � �/� F�D�~s�fMh�3'�Sב6s3�%��7oeeeC�i�*!�hemrWW��(P��|lCn�]g��k��o��}�nN�Ts���Y��^�^��{E�\�[A�W�Av���t��C�ʧ���j����.�Sn���v�慌-]�����l.�m�Z�    >�w��{�>v������c�\��n   �W:�㴢��Θ5���v���Tm�C�P�z^<Ä��=�3T7�K�Q��8�Hw>(mOct�/rnX�A�	{��|6s��S��3�m��:������~�R�+a}��\7J>b<��j�:��`��[L���j��3[�ݛ�UM�w�;>������ho�\z�!  " � u�l����j:�q�uo���&��Q�hu/f�J�ɽ���n|���]�!����	'���0ƣp���l�d3�i��|�5٬ӹ���e�^����r)\fם�*Z��l�j�nw�2B�6�v��v�(e	�Ũ�~�nk1����
   䚿���hׁv:�e:�n�N?��k �!��������i��ρ#]�W�� �B�    �yeg�*˦Ӓ�C�{p{�Gh|���.)����EX����T��̇�3����aw�9��\d����	Y+MN��=7��ר�yY���9���;�n��:��^���A�g�ȇ��{��N>������=_H�a��&}>��1؞��p清٭ޡ:Ю*Ʋ�=�ۍ��n;>?������ �� �Q��[c4�f6�;��:���*cC|D���Mv�R�J(E���;?�5��s�{��=)^�2�G;��>�n��\�=��a���F���@D�=���7�^"?�G�E��ȅ��{��F>E+V��úFX�v��}۝�!��l�n�i_�[VV��{S�Ϣya� D��2��������c��/��o�F�O���+� �Nl����?|�     �L�`�V��I�[��x/���f��������_(�C�h�'ˮ�7Xl��EYf��vW=�|C"��{&�Aw>g�����ָ��习�g3'�yNs�滭qZ��V�:~��{:a�>��f�>�h�s��c��\����j�����{k{�?��5�C���iO���7  Z��  ��5D˻�����г�L��!��屙�D4�g
V��uI|$��ʐzW�38
V���vB�݃��xPkt��g��|�s���^��nk�Y��ϵ�y��N�F�������&XEM��f��`��5�n=�_���ڮlO=7���ۇ��� U�ϥG�� Z� yd��)��_���*ʨP�?w.��O�Ow�!�w��        D�������tYc���n,�Rce��ʂ,�����]����ZK���aAw�\����x���r��Z��A�Q�j���uNk�\��5�z���+?4���{�0��ss1�a���6�*��mm��S�e-Ʋ��9�ھ���� �	� �1��7TϢ��Pg�>��A���k����^j���A�*IXR��kfP�3�V�\܅'U&�=���e�'~�=�k�\'�k��r���{�N6��:��f��z/���ڣ�0E�|	Wa�VA�Kt�fm��|ە��,����TZ���g���,���}�[��h���  ��ʳ�-�p���E-���>I�|�!z�        ���H���8���K�ͽ����!����Y�Xb�g���k�	3=ôo(�B�2,�mН�a�L��ۍ�������g�%�Y��:N��v���u:ku���Zپ�X"�?�l�1(1����^+W�b �v�q���^)V\x�q�p��_��Z<C���մmp��!r �肀; `�p�;N�7U�y��4�{���������f'�J�?�+u�]������&X����aw
/�n7D ^�:�^��9/k��׽F6��u���:��^����^�eX>*"ZP���x]����X�r���į��v�P�Qx��T[	*ũ�{��vǐ��qA!P�{����zs�bq�� Ѡ���F���w3��ï�������!       }��ѻ�tyc�zns�
u��Lb���$]�e�:�3L���v��_�]�u� ���h��K�z�n�}�l<� ��:�
�=
�\��پG�Av/��C���^���3�>�ڽ��z�X�?O��q��v�R,�r����x̰�3�C @�A� 0����!�X9�.�5H=v��*v763ȃ�(�6��X%�b�kc��]�=�Ҡ����0{F��p�K�=��nܫ��GPMU���a�SA	S^ĉ0Ũ��γ%��G6�-4�j�	V��t�l�	��*;a�*Nŕ�v��v[q�F���0���D�Z��   Z������Ӥ�U4�/U���:c�\��7K��       ���K�6��Σ���Qow��+4���w�]��c�6�!�۔c�����g�{�]!���;e�s� ���:����e{^wN6����o�Fw��z/���=@�N����/�@���B���v�]�7��ΥXv�v��K:�a�?T��Z|Ī�Z���@��; � �$�{�rc	�4}5�ޞ��f�J��n|���`If轘�܋�����@e|W�e��[�=��������ݸW�����`������09��QD����$,!�,0&���:\��e�1��p}1~��t16� ,�BB�&�
	�6�<;;3;������]�U�=�=��<�U����ݙ�>���mC{�Tq����S��+�4� �$�!�%�̨k,�h���v�Z���^��.3���/(��v��JmW	T�k���v|f_��qS�"���f�'��/F7�ԝ����o|�m��c�A!�B!�3��<~����;֠8u K��Z�,���^����X���:_FY/�%e���F�F�;GU\)�B]/n�1�qI�������5�o�Nܵ��f��e~3��c�������v0����f�X���d�g��G�0�4��8{&��{�\��CBHgA�;!dE���~����vL"w�``���T�ҋUA�{:dr�Y�p:�:��,�=���5�W�"�AP��*\�i�=�fN����㌉3N5V6^7G5�d��:Q�L��Dҟs���E��`պ��ϯʟ����{N�خ�D&��P��-x�)_Q���n N9�������8s��j��BړO�� ��S��������΍��q�'F������_�'�� !�B!�t�"p��"6�]�������i�(	�2�f2�]�3�w�齱��I��$�����V���϶��c��/�c:W7�f��k���F��c&��V����n2�]j���f�	e�4���Ac�>��ZS��}>%�]�%�X��G&��;gFpxw�҉��NY����mc�q��4f�Ψ�ڑъU^�{Ɠ��ن0��`"V��M��u��sx�!�'\�m�=�tN�}���#��X��y��6kخ��sڝV�ZI<'���Zi|��*�9I	SBc�����]%L٤.�M�E��]"N9cu�v��� ��p��"|ew���A!��'�~ ��ǿz?>��W��'oю����~�Ÿ��u���*��\&�Bl�����ç�y�����k^�}=~����U95��>t��D!]��s��!<c�*�^:���Ey0VM�Z�e&�t5+S�vk���B](�������jT�BY{+눦�M��yQ�u�G]�v=�X�x��\��&�D]ӆ�6�7�f|Nq׌��(ɱI�[�����L�6�a�z�O�����vQ]�|U�����QR۳==X߁��:�v��	!��R���B�Ƴ.ê���U����D���g�s3�T��p�VoA(>ĦvS�;R�4wS���7�pՌ���ү[?�:��َU���3�k�F���>g����%�Z�$Z��tc�!h��`9q�s�3�#,T��)qJfrڋ�R��$/8�v���~`)�!���053�_�����%xٳ.3���{:��e���Oczn�B�3<Ћ[�������+�?åx�{n�<�'ֺOܺ���g��lZ�
����@!�3��`�}�p��<.�:�Ɗft��ce�C���&��L�T7��B�|5�XFwu V���ͪ��J2�j��q�����ج���V�>�z^�k���۩��R�n��z��nin��u�X�ݞU�C[c{AQ?Z�	w���	�	!�����،7/	E+��@� �5����U�av�&��7��z�mA�2�����o��bV�;�NQ�+*-���*[�i9RLװY/���@+���ψ:��(�q�(XE]���v�0�0�{�f���-�>A��Id�6�����}xl�����yBi>K������ޣg�~�ќg_�_y�����I�>r�B���?�Gs�CO6��{�Kq���:뽏c����J
=!�����b	�}<�K���%}'17;�B�����Za�������3鴴f(JxW�
EFw��V�Z���֕�������؊Za��	[��['�I<�i��g�f��m�'Q4�jS��/���}���ZTG,�$al��ݭB��EiZ��~hR7��XC�8�[����3!�����B��/TD�+7����1��]h��%�"����^7�ׅ�tM�R�V^c�hB����]dr�}BCu�@kJ���B�l�8k���g�jl��9�sMְ]+��q�򱵻8���׮��J����^��w�2��)��=���$�|[

��u$qJ��༎XۉO�w��e� ��N�����[����f�o����5���'p��y#���������$C�?2\�͘�_�_�[xp�QҎ\�k#����+J������G��p�__{�x�SwT�3�_�[�ɡS ��P/��]�ŵO����P?N,͢�x����<��!���<z2����q�I�`i�X��.�cej;?�ꆞݟӁDw�Za��.��ꄲ�Za�SW�5�Wi���^��(곙�?꘸�����k���I=�ShU-2�s��_N3��85����Z?��mRs;�glW݅��ޠ,�k]Qu�u�R��:ar+�����3!�����B<p,��ӫq�4J����(�Fw��r��	T�d�h%JbPA�JezwE�PbC���	W&�����(P%adoq�V0�)Z-F��Yݡ��rW�)ZQ��k�	S�6��]fn�S�Rja�����-�S����<Vo���8��vBYN>�����s���#�}���#��_�w�ӝ��/��q^�����^�K�m���;�ǻ?t�Y$"���;7�s�y=�{*�/.������
��ןǱ33�v.޼���_�+/�To���]x�-�$g�������w�?u�Va���<�S�gnw���V^/���>��B�\�E���El^��M���ٓ�zB�X���탱j;=W±j��tc��t:S�:uÒ�(6��0�;���vqHVR��f��ev��3&�8��(�esL皬e���Y�$����^��6c;����CQ��=G1������R�v(���2�ڄb�r9�N�÷N��n&�B��	!D�+Z�l�s7�p���Ƌ������
ƂU�^��^��i��u��n&Zɶ#T��+S@�
&4�W^�s��[)^�ε�Or�l��zQ�U�1���o�NԵ���f���Z�ώ��r�VI	[� Xٴ���ʟ!a�&q!hn׉RraJ����D���v���T�v�Y5�������P��%��*���=x�;?�y�k�qrT;>�I�O��\r�:�����|��veۺq����I�~��w�'�~�����g���.ϼ|;���^�_z��v��W\���66<�_�ux���H�3�׃���ո��m�����������ٲv�?�7��6B�|O�q�� ��t1��8�/�IC�t�X^c��v�A!]������j�06�7�%e����4�CP+����^�.��$k��#��X�x��\�5l֋�~7��zc��[QG\�b�1�T?tk��ks���6�#z�5��4�Cݎ�E���m���8ݷw�uj�Ԛ	!��b��|�}<�K��ē�`���P�*8i��v�A���v�Ӂ4w��=�ۊ�6����.<"Wbӻ;O'8-gC�s��o�N�q����9����M։�f���T���-�p�ѪU�vݘVVI�	�Q�k� 垅�v�E)���.Om��.Ȅ)�8���ٞ,�l�m�
�ϖ���n<��D%%���z-��u��'Yy�����ƅ&��#�tJї!�DO6#l���w���1z����7����W�˷����Ư���R��N�E�=�����w~�B�������$nڱũXZ
�b	v���EuB�>�螮��ݟӵ���^<µC��=���I�0��@Tt�hM�^�lC{�Zb��Q�Q�wl�9�y�kخu�($Y�l�e�S+��Q�$eV7���N�6�]������v���X��a����vO����܊/���B��	!ĒGN��hjϽhٹ�X\\�T2���hUOe���}�L���c�V1���/�������/��fn���k�g;V5^5G7�d���k&��v��WR�k� e;>I��J�T?c�"���njn���4��S�����;���;�z�:Ѓ��o� ��n�1���|����YO�a4��/����z��=�ĩss �BV����s���Re�V��<\�]�����Ç��n��y�D�8	B!�A��������u�9}�������2��Q0�~UIt���+��42io������U�CY���ae-T+����ܠS�qj����1����	uu�(�E�<��6kE]7�hJ�Ѭ�90�'Y4�I5BU_�����ިz��5C��uĠ�=�`,��a��S��}dr�ur�v3���r���B"P*�pϾ�6���K�?}H��P7�[�V��Zz{��^3��ū���o V��V��(��c|�E,��=(^uj�m�16�Dc���g3_�F���z^7ӌ�A�5�m�o�e2�S+���L�
�	�="�J��nl7���2S�ij�t;A�0���02��yfw���!���[����_��o|���k��\�k#���7�����!��R����#�|��?����~�>�G��h����w|0����7]�?닐I���;��|��q���#���!�t�g
�m�Wm܅��0;��f�Z��ce�i�3��au�g]�Pot7��j���ݩ�ðD&wO���6�����Ю����7g��X����t�mױ]ׄv�Z��fR�n���v|��u��P?tk���`��gh�T���!6s�ga�Г�^Lj�g��}pdGrk�=Nb;k������s�|��vN��U��03uFlt���]Ѫ��P۽}��N�Bp+B_�{����Xw�_�	Xq������+���C��W��:&�$Ǜ�3�o���zI<�i����s�md��*C�ɘv��)���ڤ����8��R�X��*a�4yAgn����ف�𕽎с���iʿk���_��#��_}>���v��uc��{_�W���x��iB!�NoO��x�;�c��������ct
�����/�o��2�h~�_�y5���7�>p!�t����j<�����Vw�ݣ��{��i��d�p�P���EuBU��^3T�
h3Ǽ^���v�c��j|7�k�N�5�~v�ӌ�3Κ�TGl�����=�z��0Kan��
��v������r�3��w{��:�k1y>��<��!��Dhp'���s6��SCx��1L,��¢��.2�{�L���@��$�;/�3&_�J���"C�N�Bɟ�Jw�
Yu��T���iN�{����3&�8�X�xݜ8�Lֈ�^�g�t���R�J��n:n%V��=���@�����f�S!c���]+T�Rڝ1����ԉm��~ W`�!�t:��>�9z���:6ܯ�qr_��o�k��_�Оc �B�����[^���%�o���o���½������;/��'�7��j����{�B��B�T�zrp��qs��C�l����X�za:�������&F�p@�,KV?@#�]P/t��Z��T/����K���u�f�u��(u�8u�n�ju-4��E]c���PC�:7������m�b�j���y;>7�v(Ih��<Wo�=�{q�N_!d�B�;!�$D�����ѓY����P:w��� 2����#Ni��Gu���6���kpw�+q��_��
`�v���J�R�VH�&5x�j|���,P�R�JZ��*�A��K������%Z�����v��=�2����>w����+J�
Tbc{8q�&�����Z�	�8ևS{��N!��7ڋ�����xu%�U��� >�'�����G���� �B���l�����MO�X:��Ǐ���/�S����s�߾�Ȥ������N��/���@!�{9s�������ɝ�j�<�O��E&wQ8�*KT/,�ϕ��t�����[4��YP/��~X�!.s�0�z���g[�z��:a3j���;�+I�[mog��Z�Y��u�V���?	û��n��^4��°LM��@�(�v���X��G���,+���I<<;��vB�� �����0�B	w�.a�+����ų��"U&S9g<��x�3�{��G���+)�{��v抅�F���]eh�ۅ�D�B�>���;w9��Q�u�G]G�Vܱ&s���͏�V��mh�a��ĳ$?��ku�hWpҍi�`e���Kk�S6N�r�('��D���*H�)�HezxS�[	��\.�щI<p~�w;�v��	!��w�,^t�?���r<����}�Ļ^������g@!�t�����x9n��	�1������),,u���N��գ��.ߎ�/݆o?r �B���g
�cWoZ������ka��>���f������F�{�V743��v�.Z�e��RJR/���F�$��~լ�8���c2O5�f���xF'ӊ�c�hE-�Sk�]Q?�=}����=j��ol��G����5�����ކ��w�s�gBq���B�Ĺ�">�;���;p��,f�G��Ne����e�����3��(d���sc+Bw�´O�*
�)�x�No��D�RP��Լ�R�W��̵헍1W�R��:G5�t��ZQ׍B;�ϣ���!�ڝ(Z-�`����~��T"s{]�
�SPS��TC��T%�0��.��m`0�=�8�D"U��ў��s�#L��N!�ι���O>������M/�F;~��0>����uo�B!�»�p3���'J�S���S8~v���~�۸l�z��Y�)ǽ�Ƨ��N!+�����`z7^���#����vۚ��ѽ�F!�c�����eY~�{��,�}�xh]mPD�^��Wͪ&mx�;�d�j��\�5l׊�R%ɯU�k��jh׍i����X`��α�F�
�>c�[O�R;���~�w2&/¿�-"_����M!̀wBi2����Wo��2'1w�|������t����zPbt�$4�[����긆ѽ0��ī��p�%O�{I��,�������(╮�*۔�V�2��ۮc���NHkX.�-����n;����ɘV	V"�{4�W�i��SAs{�^'D�M������h�T�ąb��n+N��$i�nOo/��[��}��S!d%�/��y�?ށ���{���d���;6N`��!���!��l���9o����}��-���x�;1>2 3��B!+�|�koý�p��"rg��Fa��1�v�c��F�U���Z�LwOůF�V��k��M0�m���(�Q��'�u�n��|ӵ�X��iv�1���6�یo'�{�L�?������ZX?Ԙۣ�c�R����n�2c{QQCtk��`,Y�й/��X�	w����"!�����BZ�}Gr�~j�ܶ�G�����j[f���*��=]��F�t�yX���Waӻ(�A$T��#�w\I��P���jv�6���Q�����5]'�I>��h�����6�����_�����e�vq�^���Ku�)���7��D)o_P�%/�D*�[���u(���8��~�B��|�'F��W>K;vx��wB!+�o�`/��G�mL�-�o>{/����@!��]*⋻�#��0{������R��Za�0+����]�tZ�%��hlv��/F��^��Kv�@{ۖ��n�gL�q��Q�����ͷY'���,�Y�]j���en��b��[Y?�ĊR7�����}��'ê�-�۵��ڡ3ndb�sv�/Կ��B���N!-�TJ����]���
�U�!��]�*�
W��z��ճ7��*<�fw�V�A��3���UB��ZD+�`����yY��~]��[�J׿�U3����1���k���I=��i���ĳ���ܢUR�V;�ڽ�2��J��\��E����]����N�!>U���2c�I
���^_�]�z3�u�'vS�"�Re~1g4��� �BV����~�#w~oճ0ĤvB!����^\�v'�<p��S(z�5à���p4�t��^pj�Հ,��銮��
�y�T�p,�к@,i��фe�Bxj���)I��m��Or��8��(�ustsM盬g][��l���|���m�v3���4�~轎U?���jMj�~S�8KV;t昄byw{V�
��à�]XC�axt��V�+{���B�C�;!�,sK�J:�X�V<ws�gU^�z������D�L�$_Oi(��kUE��V���oBC
�t�`��+b��U�6�@)�����&�T�cf�X��~�x�Jן�@�t�B3tsT�L暮e���Zi$�5ie���$+�q�Ni��*W>*<���.�l����H6��*I�ab���.��y�L��}S�ط��!������.U�)�����R��?!��Ng��"�}�_v!�������(��m�K�1a���s=��S3decc5v��xj�ձ��u�X&�wY�[#,���B�{_�U�FX��k���4��g�4��̍2?�:6k��F/�c:W7�t�(��褠��y&��V��U�_��iW?\�ꉡ1�uCy�P����j����Xn1�ecn7�r���!Ln�W:�����ބ�hp'��e��B�۝��n��O�g�b�#RE��9����h��oE�Mh(8�����P��"VY���L�$43�'mv�2�t�8���c2O5�f���xF7�
1+�gD]c9L�-�`e*J�*A*hh���P:a*(R�D)�����S۽T����ctb��M�ѽN:/�)B!�z�w�
�m_/��*���2>��A!���`v~	�B�	�Й�<c�zL.���B=Kdv���[� �]U��Za����Ou�c�±��Bw��Ю������Ix/٦����n�/c:��u�f�Mkw6�I�WjPV3>�kv[(�ɘV�ڽ׉�k��u��9�ebp��ښ�m������4�_�W�+�vH!Q���Bڀc3|v&�ͫv��0w�2�=�1��ݽ�����y�"LW��p�	�ݽ�U�DwU{5L��aP�j$�7�W�%6�&5z0����c3N4�f]��U�L暬a�V�g$��?F�;I~��L_���J1�dL�M� �d�.yAdjW����5�&N�S��V�R�������V��}��=B!�KO6���W�K�I�8�Z������}B!�{��+!�;
�7��ѽ'��ݖB��,..�j���,whC�{#�V3�
����ݠ3��kvO�����p�p��i�P�elx70��k������7g��X�x��<���kخ��ڝV�%�1�f�r�e�QL��Zb�@�(�X*C��nX�����s{�f�����n�U��Ln��SX�Q�]C!$
4�BHqx:_>��5�W�������*����4��E,�V�+Sߎ0lv�OtW	XJs���
V��╍��;V$^U�,�@e*:%�����k��g�f�n��f<ힾ`;�U�v�1I��E����.PA/N��(}ꂙ0��m#�M\T6�	����^qjpx����N���B�d����m/�O_�K:��vB!�{�U��B�=�B	w�-a�w#��������=�0��k�L��Za�Z�s�a��.�Z����ٽ��:}ڀ,Ϙ�x�+�7�;$evO�?��q��I�Wͳ��[#�zI<k���ץյ�f��P,ﵸ~Ni�^�������bi���X��[p��fN��C!��	!��}�P>�����������>�L�G.V�CbU��6����t(��/Z�����u�v�X���̠.�/X�E�� ։U+ĩVSq����⬳�fv�q�����W��\��R�I&�TP�2M\���(#a�.H�)�(�^�Sn�+:��^c{� �$������_^�K�chn'�B��|�wB!�[*������V<gS�g�w����J��*�]�Up�f�J��thY��,ѽh]/��9z��F(���>f�f��S�Mj�ɼ��۬��3��V��#+ʼn��^��~hS;����Xn��&KW/�1���׳r�y��v;Fw�$������Bژ����Fq��Il�I��L#�0�{��A�J.V5��΋wg�\��
P�T���%Kso�W:s��_���	V��aa��A�j�Ѹ���������7Y'κ6����Y4�s[�j9L�E�*J���qE���)[�{0�]lj
S��V����8��J0�䅠0U(���ߏ�ѭ�}����	!��y�n�/�|����vB!�����!���L���)lَ��-b���J U�&�0��±d5Co{�����T�Y�P��Ov�6��4Yh���kVI��^��_˶'���qꋪ�Q׋󌨴����?�V�m�tf(V�OߵI��=�j�qꇪڡ��4���É�ạ���&˙;�z�=ч�;����B��wB� �}(W�sWoZ����1;=-��I�"�J���	Wn:C8��MhHi��Tw[�J�ր�f� ����$*�)iq���6�DY7�g��!t%��8k,w���R��Ȧv�E)�X�JYP%.xSt�viZ���^�T*qJ(X�b�����o ��-���"���!����ů��:i?��B�ʀ	�B���L���b��.<m�fN����u@�]��j�DwQ�Pov�����B_}���)y�!�.��m��b�_߷	�J2�*�8�X�xٜ8�L�ۮg��I=H3?��Ċ2�SB��5�h�C��)&]?��E�<�M�f5Dub{�;>;s�'7�N��n�	!����N!�}G�c�z�jlϜ���s�4�um;B�m��>�nr��W��y�������TwSs{���L��aqJ���k��J����Q�����7Y'�I=�[i���U3��c�ѥ,4�����Ȧv4)��Qڂ���T$�= J��)m�T�j��p���iJ �bƛ_t-���gJ�in�l~꒭+z��r��?B!f,,�A!�4�}g����v���Dw�.вCU3,k�<��y���^ب����UcP�'���uB�k�:�{wl�.X[�cE�6��+��g�n~����mB;�e-w]3����n;���?=��{+S{m����t����^�%��k����}5Ī�ݴf%�bl_��?;�}{��{4�BH����B:���}��0�]}S�9w�BOU�*��v|��4w��cvW�=�n:C]��$4�5)��?��4��F�
�W�������L���֬�i/�*��׼�t2�ɚI=��h����s�-}�fl���{[S{Q�T�R���L�!J'L�M�6�TE�����il'��W��T�ɛ�/���y�s.�+���y�������σ/�=��O��� ~|��z�O@r��BH�9|�P>�ؼj�>��4�g�XYA0��fX�/hk��`,�ٽQ/�	E�B띠�/T�N��ژ݃aX���k�����Ǌ3�t��ZQִa�M孠[�l�%Y4�|(����#��S?���Mj�E;>G	�
cy�����ؾ�1��?3BH����B:���� Fp�q��¬ct�d�[J��u�����Mh���S�i�v��*lz�W֢UL�����,�ݡ�w�ؤǫ���׭e���Y�$�u��^3��6��&0$���^�)�����J�����lA��]������.L��s�@�F����E�4�B���=�/��X��I70>2����yx��n!.�_��닰k�d���w��%>5Bځ�S���cgf0��Դ��d3 �BZ���|��ݯ�\ąSG�N��B��]op�c��I0�,�]�t�/z�Phv�^���(�����V��p�8�t�mױY3�����&����U�3t-�ދ�[ej��AX��D�nϚ��vE0�kl�ޙA���B��	!��g��T�(��*�]w]��3C{�Y�L��^��Fw��]gt�%ZE0��Xa�_�
��t4S�R�Mj��<���kجw�n�BVψ��r�Vq��{��]�� � ��(%J[�Q��R=e!dl�R:a�(��+F)�)�	!����W��?��e��=����[p�3Ǧ5�p��eR�K��3��e��n�j������7��rL�&��7������~�F��A|�?��󝸰�k�s�{Y�#��Z�F�6�ڎk'��Fwg��[�=fwS�{�Z��N���mw�v�]��R3��vh���:8�U��V�	��M暮u�$��h�ע��XQ�td(Vm�I�7&����n����kl����#�B�L��v{.T�;�z#���P]#��.�5�_�i�{�p��)�=�D��#T��EB���^7�=�fFw��]gtOJ��	Wrӻ^�RWĒ��+��g��Q׋�~�a�oW�,ɏ���U�dbT��&��)�Y$L!,P�B��R���onۃm&��+JI���8�����kq����B"s͓��÷�
�=�V��I7�fl�wR������7r�{��I��ן����عq�=�G��h�3��4!�����t�jtێ�O,`���ݟ� -��]ft��ܫ5�zm�`Z/T�dk�&�l���fA}��s4xO�*C{��k���%�c2O5�f�5�zN�Ҫ�rbE���X�{��]gf��Uw�N����i��e�=ۆb9׾�����88�	�9ُ�4�BH[@�;!�t!���>�I��q��fOEڛ����>m(Z5�_R���.Ou/
�դ���e��^;�J�t���U�oU��w[K4.���9q�η]/��QiW3�	�����n��M� 7e�'FI����v��]�� Ml�l%hcp�R���U�8�I�y(W��i�!��˶�ǿ��5�����N��S�x��)BH'����'�!���>W(=X3��m(�p�0��4wQ8VV��n�tu�碸^�	�Y�-?�M�nOY'�uBQ}��0��k��Ú_+�p,��&kDY/�sH�_�Vb��Y�P��g�P,�k�I�eFwۺ��~�6��Ų�r��'7�;�{pl��Ec;!��4�BH��ӹ�ы�c;+[.�9Ry���U������L �Amp�EFw�x%��fv{�*������9��%�9���cM�ę��e�(k7�٭`9Ŷ$��*#��$��{��=x��`.F�V�w#S���]kj�Ra�z�12�?��
t��w�)
քB��k�$>�?�����4��n��o�:�s ���	�BڅSs|q70ҷ7lR3G���X�Jñ,w�6��
���ڢ��]it��5C�w�6C���Vخ�X��6kجw�n����$�oE-��k��dvQ�����6�G���ljl�
����d��l=�[��i�;�۹�3!��4�B�
��А���필�⹪p��nC(Hq���%��kG!�nW�9[6��īD��oM��gub��oKoxwƸ�q�)���sT�L�۬eͤ��-4��mu���<��*�)x��'�IX��ݳV���%��L*�ąVۃ�T�ޙ;�z���NZ;�X�B�m�8>�'��ի���4��n��؃��u?!��ѓ���BH{1�X�����ܰ%�U��1��n0�%�����Xz��xG�X&�`[��_3t��n��
�}���5���g2�d۵��oK+L��V�l�@��s���.Kiw�6f��M}Poj��뇲 ����8�C���?Џ��|� 0��vBighp'�����0Է�ڒBj�(B��.�l�A�*$RL﮹=,`�ܛkvwϦ���3*��-���]8J!dU׷���ʠ�o��͚I?�]i�����Zad7����6�%Oi	Qq�)[c�wKA�%�B�$Ol	T6┱0%Mj�
S�ԁɍ��>��@!�$������^W9�p~O����E|ꞇ@������i�&�b��H!��#Ky��}dRk�S[2X�S�;?�L&[Im/xM�
���t:��!��U0���.�#���}ú2˨Vب��;3K5�t��Zq׎B��ϣ���#���6��Ƌk�Qj��P�����y�P�'6����v��(6��LﶡXEo2��v�0��142�ٵ��@��HS;!�t4�B�
dn��;v�Л]��l͠g��/�V�+�P��sD���-hxw�&�6����H<��*�>~�{H�*�S�e�jbCt���?xWH��0�����5]'�I<o%ь�I��/�'Q[�v�lml�_t
�ۘ�U�vS��q��:S{lc�H�*�����̃BI���A��ǯ�$�����B!^F�@!��3����{:�8�ܰ�����(d{�fv��=_3�g"ݥfw�`,U�0z@��͘P��5�W)j��tw�{g�c���ͷY'���zv+Y�z�rbE�ۑ�Xh�
��q�Q�������2��$�+���`��WM�8&q�\��f(!�t4�B�
�Ih�ko���mO۸���c��I��[����Q����I:C���¦wo:�_�R�uVbIn_������W���V��qL�9&�Tsmְ]3��t:���xN�5�kf���ڃg[�*�������5���{]�
T­���R�c���(�zW��X8Y��A!����	�0<�9�/��;_w#��e���1����vB!�����Svl !��)<p,�0��n�O����'�L��@�����`,}8����R��lk����q��=�����a��c���7Y'κI?�[h��w�V�bk��1I�����Q���ݞm���FvuP�M�0N0V�X���:<va̡���	!�ӡ��BH�MH
���>b��.\9���3G��吕l;4��W�6_2�"��'ZU��)�\�����(����`�m
ux���F��P]����bD\Aj%
PqI�k���(fvQ�J���k�ܳNhR������]-N����%�(��n+L9���$��qW%q��vB�^tݓ�O��
t���V��	!�+:�?���^S��zA!�t��!`��N\3�G~�(�&wY�6+X7��c�$uÔ~hS��C�b�Ѩf(��g��=�i]�O�±L��曮eݤ��δ�6���X&s��Նv�b��.�/F�ǩ°T�X���1�;=[�5D��{��F���>���s �ҹ��N!�Ǿ����h�6<cK
��cXXXP�ӆ�h%Mo�T)���#V�,u������ ﶇΆ����+dU�*q*���%Jp���-`y�)[A����4[�j�p%����P�v�%IV�L41��ۓ2������K>!��KZ(9�Yj�h���@0�;�6&6����س����@!�DO6�w��ft����3��B��u�n��.���ĺ�a��/� B!��9|�P>R�݂�7�'qan��ӳ. +b0V�:F0��f���k�q�����u��|g�ذ�]M�.hj�O"K5�t�n�(�%���H;b�η�#�k��6+C{m�V�b9��&5�j-�����I�j�1�����&|�H��P�B�thp'�"��b	w�.!�Z���҃���9w6dtO7S��4��vW��W�_̒	W�k���!�p�4��g��G�

Yr�Jnz�!(�J��#J%)�,�Y�]�$?;V&@U�۪��4BTm��=Ч�T�]֧�䂔{�
P��D�*�*]b�N�*Z�T}����&�{$���NZ;�)B�D^�`�1tnr;��B���'�)�����!_(���G�x���#��t���%B!���Rw�2�5�r�zl�;���'�v��6fw�v�n/ˬfh��N(4�W/��@����\�W8Vu��Ȋ�n�u��bU���ۣ�U�X��ø�X��p�Q7�٣��,7����l�
��cx�N�'��9*_�!�t4�BQR(�p�A�D8������C�1{�DE�		V5�Ig��m7h-\	D�T$�{X�
�''\i��:�{@�r�t�"ӻ_����-U�C*Ԟ�0���b2O�f~^�I""��Dl
�Uۍ�����>�H%��������.3��)�/(L	)ߘ�Z^*�@%�T&�|>�щI�(M�s(w�JEB�\.Z?�n�5��Js;!���=�6N��%7\*�[���ʹL��x޵OԎ���kB!�E��>��#y܇Al�؅+'1�HE��x��@,�]�ͮ��R�z���ݮf���~]���u5�(�X���	v5�v	�2}F҈>�N�?._ V�O��`}Ѥ���хb�ꋒ�$C�d�2C�I0�p�g���_[l�m���*��;�f~pn?9�ݞ	!�����B�1��!`��N<}CٹX�_���t��]gxo�W�����6��d��^,`9D1�[ޫ7���M��P��$Tɍ��5S����L��щi�%|EKè�i�'2���M���kk
~�)x61�R:a*(H	��KQ��$fv�*$Li�|�g����p���0E!��w9��������4�B!�8��o���U4�?��n0�����o����q�}�`�5!�ҩ�;�/�ڎ�6Q:���v�B�.жuC]0V��(Ʋ����8�w�}�&tv�Hk��;<}�p,����F(C��$��&k%�~3hW3{�?�$�����p{�Ϥ�(5�{��bk�"c{5C�ݻ˳��=�3���^������ݞ�ñ$��j�{}�}�ݞ�s4�3��BV4�B���\��v�#\�+7f���OW�U��$��L�:�*hzO����]���䞄�]kx�VB!�}�h'8��(43�˷5ԭ�Ώb����� ծ�R+��5������r�{���׆��(���ꐛ���T8��+N�)�6�:qJij7L_p�9I?ëVa&;�of�P�"��n��؃�����]����Ӡ��B��1���_|�����'K�u���5?}��-?�5|9�%�燾
B!�p�_��7��j�6�TJ�env����B^3��=s�5C�"Z���������%�7��&�d�f��	�
���K��D6�{�k���X�`,�:���.1�;s���D�j��ݞ�q��<���BV4�B�Lc;�~lىk�*)�d�u�J(b	�+YJ�R�&4H��A�k|O����M�a1�!	�*$by�)Q�J��Yhl[l	Z2�Vc���6�W�Q�Gp�A|j&I[*���/#�t}F�g��Z��
Q2q*	C{�^$FE5�{�R@�
'��|��ȸncn%.�)�(�����þ�a�Y�F��!�t;������!�z:O�Z��q��!�b�cr��?�>����g�I�q�hr��\����a"�|����?B!��������Uy����l6[��j���mS�Cm)O���V�Ɗ��Jw��ܻ����>�ñ<�m�p,d�>��]_wl���8G'��b`�����k�a�����{mSOl^(BuC��]\K���D�����S7��h��*C���.�!gL>_���A��F�w��9�D�bB�J��*��Bڒc3|q��l�u[2X�������f�v�p��.2��S�S�kٖ�jӻ_��9؈X�kibC�F�2�E/�������;#��ޤ�O�hl��O:T��X��]�/�E��Jl�]��'�垛'N���p{��.�����L�R��m�*�@U�D┛�>84���GҘ�˴vBYi?K�8!�����x��?�����O���o��z��/�d�C=��������!��88W()�d6K녢�a�-X3�_7�c����p0V�P���R�{� �{�3���r�Di���F�>	^�n��xm�L�䠬f�@u_�����^�7m�~\�5EUm�=C�̃��;=��%͎϶YZS�4+���1��L��E,�v�BBY���N!$Qr����1)�`��	<u|KSǰ��'3��	vF�t`{BW̒W)��]$b��+�	���n{:{�A��v-Jx]����M8͡*8�����G�7C�5��x;C�h�8󛏍9]=_��L4���^_!���{�2��LM��k[C�J�
����!C{@��T޴���]gl׉UAQJjj�;��\���q�Q����vB!�BY)8&�7��3���{9�w�������4���8z��`���9���?����BV�z���q\1�C~�H�^(�ZV'�ޛ���v�n���B_�Ц^h_+���	�7�6�����z^�Ɍ�*�L�Y�ݩaH�x�J�r�����Ƅ�����͌���tufv������C�t�Cq0V�nhalW��U�DmZ���2����3�4&6��s���!��L!��B�ƞӹ�Aov3�٘�ƞY̜9^IiH��+���+`iīHF���� �\KhxoM��Lī$�J�;�bV��v��F@ਜ਼�K�Q��1�D��2'l���,���.�W{UQ�g�ƈ�ebS�^y]�Wؽ׆fv]�I���]��`bh�R�T��v���I[���j|�hg�0��B!�BV2�|o��O�C��7_��UC����_��O�BY��;�/)�n�������?7��ct��fw�u"�X���XI�ܓ4�k�)�p,�4Kb|��냺ڠ�o��wN���l����cb0���~=q=0�@,��=0�& +JQW+���	�2������K%�UIhl�����k���v��a�����<:>����~���3�B	C�;!����T~r�A��H?֏��ի�Ν���d2Y��}���uaʻ-������n*b9$ep׉Y��ꍱ�]�X�{�7���<�T,2����S�D�Jm�H`=��1V6��05��j�6�*1�='ip�nl��BT�2�{��8�v]�H��R�4��f3���G���#Lk'�B!���1�����������\�t3_��Q�z�C �BV:�KEܵ׹�Ήո|"����X\X��b���@]]P[7ݽF���XqC���Z�c	�M±t�º�����6hRT���z�x��-�h�g$]�F�0,�q��P=Ѡ^(�K����u3C���X��v_���v�nϽ}��ۈG���N���\B�C�;!���r|���g����tmO]���c��s>����=p֙�e�+:�E���=lx��M�+�������,�����{��%}J1�+V��6�������X�3Ë��ϗ����<{q�[�)<_7^g^�iE�ڽi����4�!��]��P��瀹]jl7��+��$�di�θщI�(��;�
ȝv�nL[ �B!��<犝8��?Z�{>yQ�����۴I�́S����7B!�Ϟ���B&�Wn����Y̞=�\.�4��5�[�C�B�N�㻿�'���[���e���u�޸>hXԙ����Ў�|
�Aͩ)FC����m°��e���������D�qk��5����A#�8˭�k�>C���]�ebl�����58Q���;�|�X?$���wB!��#'��#���\�9�u�)�?{&�� ��gK��䨋X�{J%b,�x�>��w0���c��2!+�}�-�iڼ��pl��Peon����U�iV��e�AqI�f|_k3�tF��9I��q��Sz��+PM�r#�IR�L�2��Fv�UOiS�C�H��}��G�9�E)B!�B!z�$���J�|���&��x��?��� �B��B)����q�1>��l �g0;=m����n�h�0��(�=x��
�ꄭHvW���x���*�{���*k�A�g�iM�δn:����x�?.��A�`a�@��u̍���i_�v�@,�0dj�E�DO�дVh\O���C��XX��<���}�ѝ�CB!v��N!d�Y(����~������W�$L_8�s��@��3��|	2�{�6��	�2�{c�_��wHB��1�{���4��{�i�XFm�>����k|�%�vEfN��4����6���BT���>��mL�"A�onOX��U�v���'����3ۏ�����)B!�B!v8&�_�����w�Ͼb��������� �B�S�Eܵ׹Ǯ��x�x��cX\X0�jB�P�%2��j��ڢU�0Z-���NhZ��_���>�z����f�h75�{��R��x�:m�]V}V�������^(�������c��~B3��.�%}R{�ڡ��.2�g2iLl�޹~<pĭ@!�D�wB!mž�|�pD���5���W���u��(�]`z�	X"C�Ѷ�³�ɽ��nfh��٣XqD*��]3&t]m�ߋڂ�y�8o{P3�2n�	
?Q���L�CO�hh��MƘ�EcTb��.6�{�%�(U=�)�e-T�"S�̮��&���|�����0��p�S�W��vB!�B!�XX��������ϼ|;:����wp�� �B���3��B_v��1����={�R�Ig��P,U���쮫z�}ie�P`v��e��t8V�s�ڠ��%m�z�uH���g��]�I�`���	������%;����E3����b�ñԻ=G�!
��5Co�X,T��kq"?��<�������!!�����N!�mqūLj#._����,LG.�'5$`r���Hh���f���=$b�c�X|Xܒ�Y�8۴��f���Mfz�{��k��Dka*e=�:JA8Z%<Iƕ$}Z㺤-��`"@��L�D3�W?S!J6޿e�����F��%7��(YH�Ҙ��BV��qc��#%�NAQ�B!�BH�8&�_z����^����-_=~�4>u�C �BH|�%|㠣Gb��"\�1���fΞ���LC�du����Ʋ�	Znld%���Y٦�Z�a�j�"��M�b����z�st�D��i]QSS��ez��%����P,��]���~���]bv^5�����#��^�	!�$O�*��BV�����@��Vov3�٘ņ��p�x�[:m`vX*K�������^,^5�MM�^�ɤ/h���9�����鬒�#�v�O �Ȅ-�8� �K�z�|eo�`�#듭ob^�]�R����1���Yڂ+DU�eb��ܮ�:0�P%2�������R8���:��B!��9{~�f06��k���s�!�4������A!���b	�T��A���5�W�)̝���
�I�2�{û�v(�JL��Z�����p��k��5CemPV+Ԙ�C�:��F(��ψZS����(�X���<�qB�Lj�&uBU_��<Klb7���&�X6;=��&5D�`,Q�0��chx���w5�?�������"!��fA�{��ߛ�P_z����`_������\�Hta1�Ky��|a@Yٔ��JRC/������13u�&�(�+�uPĊ�����,���6��U�2�L�T}n����cԆwXlU�:Gi�{-����D&Ř�X���s\S���FOQ�=cJ�f3��O%>����T"��>lf�R��F���.3�Wۋ�k�06��S21�����TE��S�1�jz'���4�Q�"�B�
���<��g��C����}���9�w������ �B!���L�q�^�j6����\8�s3�d�Z�{��.	Ȓ��m�����^�Jk���wY8����6���-x-��֢�d����΍�U�1X�3�dV����nږLQ����ܓ�2����fv�`,���P������3Y�;ꦴ3���dʯ��z0��S��ɦ�ߓ��|�r�/������Bd����8�q׍b��1l����ym�m�`Fz�ۓ1Zk~)���05���.�������=>�ss� ���¹���Ϲ���(�\��dzsS'+oڼ��:c{��+`��eFw~�{��4�7D�ƽJ�r�&bAK$d,��JT+�u�{Y��=4�:�z�c{��Z2n����Q���T�k��LV�ڃFv�����AA�.D�M�k� ����*��=dbטۇFW!�7���bߡ<��&E)B!��\���}����u�n��3���{+��i7>x�����1��=GςB!��Oʇs���ۀ�GQ�;���B�d&wI@���nS+L+j��0,Q8V��Nh��uAXfAY��m_��&��v��}��,��RT���P��b3��k3��OnX����5E(�d��j{�P,�Z�i��6kphZ���������<!�S��V��[�c�Xճ�xxǇ�*;�:�&��?���-bf~	'��^��Ss8vv�N����J�5i4�7�գ�t�.�:�'n�EkG1T��q��V��I�'B�S�������#�ǁӘ[�BH��$5�S1��c��"\�!���pa����aKez�km�fw��]ix�	RRӻG��Z~�J�.��4����"aKvW�j���� �Ldb�����zc{�J*@�Ũ��]����mJjl�'-D1�+�T�vs��q\��N�p�kf�kFB!���ǧ*!�����B!�BH��ȕ�t�j-vMfp�x��Ә�'��-1�'�<���~�{�>TL��B�cnxW��eF��L�Q�u}��&��FUC�jf�5�vhcf�^�r����ݿvx��`��[7����:�A�0r�0B0V0�}`p��I��Ã�r�g9��Y?$��?��4��i�n��;7���k� [~�51�_9�����E�?y������O��Cgq��,H2��� ��\�s��x��x-6�-�������Z[9�L{�M�{�����x���c����犸�`�|Ջ��<mcz/`~�$r��\��������e#\)M�A㻯-�Ԡ2�;��-��Zntw��}ɧ.�ڣ��M�4�f��EmI	Vb�r%ik���E&v�}H|��I�>1�#^I��Q���hWR���:�j�bj��X
�:��"!�B!�B!��nd��B�p�Vc�u�t����fΝ���D�0��=�V3�7���&�c�j�~3��6(�O>�=ʽM�M�9�z`�9I�
u�Qj����Ѽrj�mk��6QV��.6�B��E�n�I��M�����A~`5;׃=�r����޾���B�_�;׏ᚋ���'��%[&�ͤ��c�ɦq�Ʊ��]Ti;7������>v��>Y�'Ѡ�="�ϸd#�}�f<m���?�v�y��~���O��B���1|���+�<��M���f����ރ��^�e���l蹀�󧰰� �D���he*V����߰�Ml�S����CFw�hezV]G���n;&)L�,՘VT�s�O�Yeh�Nac�8�AlbW'���Cfw�%�d��&���0����(��;[�3��K������#�B!�B!���88](��*l^5��Lѷ4���)��]V#���5���FwQ�P��r�8ؘ�eFwy�����F���]�n��J���e�Q녪>��=x���fv���Ԏ�Y=hf��	C�C} ��NhSC4Ik�������\���f����	!�=q~�:��_�Y�n���~�+cC}���͕��}���S���W<���/��C���������W_�k/^߶�v��=��+�V���\������cG��2!��Y̗�f�Lj3��&���y�,Ma��tE�Ɉ�(���R��1��S��	�"1Kjl�E�;�yU�
l/4�7�+W!�J�fs	Y�>յm�I�͘����U�Lĩ`[T3�x����8�(QJgb��GQ6���M�Q*�!2�����A�����|?�?Z��ch/�B!�B!�B!���|�p���.�(a�0��sN�{�W+�d���~��=��=X?T�E�w��]w ^�{�Ψ^(���񪳹�=ʽ�M�n��
�������+*���X�Zb��$KQGT��XI��uDU8�&���M`6�
��u�\s;!��/'�*��7]�kW��p^{9	���k/x
9xw|�𾘣�C������Q�F��o#=x�5�+��G������W<�oBȊ�P~S���|�p�ƱfhOY��dzΝ��RQiv�z�L�*�*���4�*Y���^�����yϦ}b��:(0�����6��L��^ӹ�^�'�V���mz#�(�]-Fy�.�ٽ"Z}�A�)	�{��+:9��Iu��ڇW�B�w�g��Jǝ��!�B!�B!���5���zGq����. 7��	:���n��nW+Tރ�((+�����ʕE}���n�e[lg�{Ts��OdX�]����EuD��]V��{�EE�Pdh������^�4�G�
�S{OoW�ƙ��;Z��)�kƝ�	!��D}�%��s�n�;��w��t���)�&+�{�Sq��������S3 bhpW�y�0^���xo���p��1��%W�-�
�� >��Ǹ!dEqj��{�9W���n�e��:����i,�ϋ��&"�+,Y
X�fw����R��bUX��o\��^iX@<Ѫ:_צ���ٴ��%GC3*)�K�6ս͵�,j��nh��Ae��(���b�F�j��=���
��'ë&1��C'S8q��ω���;��B!�B!�B!�dn��	:�Lj�o'���iy����R��^/����~ӻ�(2��{�x��r��nۧ��c���hr�5��k��uD}Qox����=u@O�0\W��Ek��M�jC���!c���><2���$����cy�O9_9��B:���,n�|3^q��e�0����,^��x�;��ޓ��w�໏�xr�����~�<���Za!��e��ċ�������o<���EB�Jb!�w$���)�X�K��T���y�N�Ep{Ba��J�
W&��M���]D�@JCX�
��������
R���8�uc��>8^5.ܯc���jI3��l7����'��Į>����u��&4�������dr��^*����(Jc8t��!��(b�!�B!�B!��8����NUt{��=�f����N���Y^?T�	E���
�ҙ�m녺Zbr�j��>���qofn�^�c���uA�����v���j�g�Za�����nXO���02>���*��dG��;<s�gBHg�ߛ�Kj'^y�0:؋���⪝k+Ǐ�Ň��#ܷ�H�=l�Ư�t	�u٦��� *�=���]x�5�+� |��af>BYi�J)��5���1\�6�-9���a��4���-�"V*lv��X�"�0�]��0�#�'4�{���
V���н�����o��)�_{��[��6��ɡ��c�}zs{p��ϟ�P���E'wl��afكb����1���-�p��t�Ts{P��R!J�_KX���l8�A<|*�c��t�#�B!�B!�BZ�w'�ޭx�,��/ �0;3c��nb|�mM�~�{�@�@�PT�E)�vY�구.������}��ă�*-�1��R�킱Bf��C�aX�Zb����n['�bnW�ڣ�bUR�GGP����><x���s���=!���ɦ+)�y�16ԇ�Γ�L�}ox>p�t�#���thpGuk�W�pq����!�z2x�3�����"|���/|w
E�@Y��犸�H����Ć'�IcM���Oaaa!$b�j��R�r�����njt�U���av���'j������@�L[���^�n��Za����?V&h����{��]|��j��5m!�/@����$�uƚ�m��&"�N��m'�����c�ό���,=�C���b!�B!�B!��.�-���CNM�|�ƚ��x�Dk��͜�
e!X���, +n V4��:ˬV(	��d낦aX"�{cL�O��oS��Z���X��`��?.z0���kV����cIk��:���hr���I�ۍ�6�X�=�P��N��a��B��랴o��˱qb��S���_�����c��7�� Ǧ�RY�w���چ7?�)X�¶6�ed�����W_�����%B!����ί�Lj#��&��9�g0;=U~#�lQ�7���Fw�uRF���U@�
���Mg�P�B�=`x��i�aa˗����}��{Y[m��R)�ar#{h����+�"Su���~�5���New��⓻���.����o��m��Q�^1����v�����02:�|�(����y�ܿ'G�JR�$�B!�B!�BH3��
��غ*�'���
�?{��Vy���-Y�{e/�w	a��B��R�h���Bi��Z��(�m)�z[n�C�-���=BȀ �vl�{H���#ǉlK�lI�����p�y�<r�ǒ�<_�N��6���=R���s�0Q�=��a*k�Z��Za�����q��kzI�����>������m}�������-Y5���K-���| Űz��'X?���3��(�.=�S)�����@�-�5��X[j��U���84�.p�7VΗ��}[2�LL,����Vy��-����p/�ˑkV.�����_��/>F��~������� @����M5AeS��b6�ej�Y�z"∶K{�>	:�޻&�����8N|��P��米�]�w�1�%'�R�K\�=Q�=�~��{�?�y��TnK]|��m-�<����=ں��S��O4%��
��������CކZ�=��dS_A�>�������J��}A�l��Hî�|        ;��ʦ��<N�XdTN��M���(C?a���Á�jtҚ��WO~����6~�Y�Gؽ�}
����#�<̞��`*wMdOt�h���������� �I��Y?�c=�`�}��}�r�����h
��z�!�ܹ�yd��&�C�ѭ( LF��\2I�|�L�[M��X-&�`�4�̜��'ߕ�>���d���_W-�,�8Sl~PC}O�7V�O,��?�����Z  ����XR6��.&�(��o��ިx��k��`GG�2���{'�'��5	5�
��{�<�u�����Uj�/���}�u�%>N~��(N�;�S{!ѭ�g��	O�	N{�;R
��?�`:�:�P{�ɦ��u������6U�Ď�;5�`{J����d�	���"ǭ�s�&`���#���hg2
       �C�?$���ȍQ���i͗�E&)w��i����غJ°{_A�T�x��t�v��N��=�x}��5Ã�ۺ_\�=�5������L"�D�n���7A��h������{��P(+>��|1q��ۺ� ��Z�&�Ǉ�5X;LV���46���(��ФU���E2�,W08�
\򳋎��^�&w��}	��j�#*���ɷV-�%SKCW�˭_X&ϼ�]���z�� �\8j����ʦ�uާ�e�7,NiK������L,�O\%���#���D�P'�Tڄ��;�Mb%�wݯ�4�m}8��<���a����6$���&	��ݒ�-�� nB�`{��	���N��C뉂�]������M�ɩ�����ړLJu�7~S?�����䖪6�l�I���;D�       ���-���t���nv��"��r��n����ؚC�Za�uB��c��^�U�]��m��cG���ܧP$+�~��$X/�uҽhV���}��ِ� V�A϶�����>
`�O� �ą���[G�8��놩Vp�V�s�p����k���ϑ�啈�#�|��:$~���[����+�R�Z��sg.�(&�-��)[+�P7b��w�,��&Ў�"�b�x�>:O~���ew]�  RV�a�e_P��3���K��$��)��l�����@J!�>����hKGeU*�}�':Nm����7$������{�(ڐ@*�U�>��I��G�8?\Ov�;��T'���5	��]�ɪ�ǉ�����s�N�9s�M�٭i3�5a	�G�w��        }S+��[�wcg.���2��$��a��[���A�@�����궦�O[:6�@�����?q��T���w�jH�=�h�u�h�ۺ�F��|��b*{=����-�:a��Þ��Yr�y�3�dO�I6XCT��`���X��5�d�a����"������~ ��������K��:L�|���/�H���^�󫟑�=����q�  goKX��#�=�+�W+4�XOD◈�EZ[�c���Ǉ��	��tO%���p[϶����{����J������$>,��~��{��֨��gx=���SZ'���s�)Q�`&�������or����
��O@�:��l���A���f�؝�Xe���E6�F����rO��        ����n�wu�5��\�\s@��Vikn��a�8V�����5О��a����W[l�y�Gہ����zvo�}��:LL)���`K��R*����~`1A[*k��Ǚ\7Li1��a�}|��۝.�i����&�l��HxE� �lS�s���K�4/G��Q�8u���/?�m��r(:��96�\w��tZ� �����s���{~���ܦ�A; ��#"kBʦ�Y��@J��2�k�B�Z�U|�M
�zOd%���U���ڵ��0� {���P�Γ���x�~�0�޳-Qp=�q�!���2A��-��3Ğ`"�@���`{�I���(�{�r{$bsKc�&�Չ��H]׳�D        Ȍ�MaeS�L��rZs���:;�c�����=��X���n8��{϶���Ֆh�_[��Άnߓ�`|�����H�z��5%.���8�uî�@�S9J�=�:b�������b����Εc��̲�6*�{��� �I����g���$H��sF���\��W���M5�l���㐛�_�42G�E���ɘ"���ț� h�{�wwl+u�d�� ֐�"��I{[���='�MZ�0qeL�&C�':�~0�}���>���ݓ��S���٦U����DP݂��ݖ �?��m�ǤTgev�8\�Z��.V�i3ʦڰt4v=/��'\       ������I-�U"��L�X:�j_K��B݋cůfr�0հ{_����6���:a���E�k�}���n��-��YOLV+�zb� {�uD�8�^��s�>h��D*k�����g��X O}����r�����}�P��^�\nx�5ٰc�Jɀ��R���eR��㘙���m����� ���л*'��9Jd|��@���EZ[Z�OX�q�k�*���@'�DR
��w<�}m��'k�z�dP��j��| !�T���4���V�9ի��`{l��"��Dm.iYeg�ȶ���뺞��PY        7��!eS��J�	�cE��h�֖��k����ɂ�����ZO�*�ߞ�8�����O�8�y��D��_�k�];��8پ�x0����!�!�8V�:a�`{���0�ͮVf�H؜s`���D뺾g���/f�Q��j��0o� ;<9V��EG�-��)/n�#��C.�>ut������
�k�������w�Ij�} Ȭ_$�uR��c+��f)���i�9�_{�t�}�'�����$U�aw��m=�Ed����z':O֖�m��k�j0���㡆�S��u/}OLI���&�������X�bW���M�}&���ڦ��:��       ���{q,{l�u˄\Á�Xa_����ű$y�} �CY3Lp�/�>�uC-���\3T�s�0�x�놉�h�'��k]1ɚa�0{4fw�s�Ø#u�|T�����îc�@*,f����r��rAvY���9G��O�#ϼ�]�T�}��b��%����?�����`�/j
þP$��D[B�H�����$�٘k1�s�c��b�x�E^�2��wc��򋋏�o�ϋR��. ��j��;���g���+��:L2�m�gT���X�>	�����&�?ލ�&�zNf�:1�j�]$��{|{W[��z�w�$��S�$���b��g[*�Pݎ{���%���'�"�BOj���p����X�!`�]MQٵ/�ܧ��BUv         U�/,��M�Y�e-�q�F)sE�m
�9엠�E|����k�n�a�u�������s�輿v-�c�0�x�����}�t�0ٕ��%v�#��9�1�]2:�)l��v�lkI[���5]� ��`(Ԝ�.X*s'�p���Ե�C�M�F_G�)��i���Ñhk8m����f��e2��V��e1�^�-�؛�t�-����Q�
�Y�@lf�<��'2��$x
N.���[*V�I�����^Ӳs_�����ۑp䅊����`����~��B����1N�uA�ǱpR��Xy���Qy�S~��c��������@��	�F���ؙ�V��r�%2!�$Ŏ�䘂b��%�K{kKlr�8�J=��Ez��y�&2��+�*2�r{�dRIo�?����q���T�DS*ǉ&�����Y	'��`��s�ɖ#a�MڣV��ewsT������5��_�  @���f)�Zēc��(&���:BQ�D��-${�����\�IJs-��1��j�����3��QeklI�2F[����$ϥ���ƨIlfe���1�T�hD���J��+t'�-!c��5,{��z^G �ε"��F��3��3Gl�(�����r�Ar�!�E��h�֖�ߓ�5\7�-�%�>\��q�%kK����~��d�d�4���a?k�Z�Jh�����՝��i[��g��ui�uug�� Zʱ��'%3����^��TYߺ��5�v[G�s�����W5��k��iv����eq�˶hl�kJi��":��
r�isc��~i�g�D�}��B�Ig�v�:��{��4�^nl������?Pq�_�=��QC��=��:֖�6*7�h��q��!�}��ƽ�Km�O  �C�?"�Vu��_M����%ϡNj�@9��C␀D���oo�`G��dS�Ė���`�I���$�K����Ie/7qߖ�8�y��$�H��z��������������6��<��T�ۺ&�ԉOu��bWC�v�P~=m���%*����O*� p�Pm�Rf��csd��L(��M��/4�4?����]>yw[��k
�cb�Mf�ct�C&���a;?uя_X�V���>ٰ�M*�z2I���9�������:�#�u��=,Uu�����]�2FuC}�W_;g��|U_S���4M���M���{�{}Mc  �pT>�+[W�=�9,E21�(��%��(�߄|���;|Ov%h��&���*�5��{W[�}�����o�;��O��DfВ��`O�n�3���z�t_7�/�>�`{��]�="6{�؝959�C,�4Iu��*����� �f��|�R݅�wֶ�+����:�hln��m�:w������5[��������;:<�麸�k?~��	n�~&�.9y��ay�Oe���i��c?,6���_�>�ll�����:��]�bo&�����\w���Jr�S�sOS�rH�����O/:J���il� �����Ķ����\)r�b��|GD����s4(��_:�>e�Ht�>./�W���z�w{�}?Ǳ]��dmɨ��J
�&��(�j�=�C��>���{lf�Y����v�m������7J�Zͬ9,ц��� �P�Vi?~�W���B����2�"�S\���/VV���MM���V	�S��s;L�9����<�^�8��X0����B�to����Y^��"� �٠V����in)e�Ʈ��h�+�]��\������8y��J��剽�{���������}�8���1ڬ�׷Į�  0��������<b5��:MR�4H�-"nSPLa���������h8�OR+Y�=��¤�����%�'�s�4+�/�uÞ�IlOe��W��}��)����Y�]=�Z-bw�%juJG�� V�2l�7���������D ���(7��T�N(=��������-���ʵ�g��|�9o*;u�����]��o���\<�<o\�v���|���������hX�$�*p�-,�=����-��{��>W�����Vn�b�{��L�����<{t��{�'ϵ[��m[�V�gG�տ{A:�\� U�m��v�y��~�*O���(�Y��\�������K$�!Ae����'��WzIp��T�����R�}�yl�����N��z�������;����j?p[�@��sױ�b��!&�U���$�|}���R���ְ4w��rS��/8�* 0y�r��|9z�[L&��Q��6���,-�g�i�g�7I��[F�68cQ�,����1��Z�ybi����ѿ���|�3!�e��ϗ�f���h2���m͑����(c���{Fx̲R���t�����������m͑���{=�   ��@HdgSXٺZ�P�+�Y���;D�֨�L�� |���������',��J�]�n�(����}�ǵ8��(�������
�S�'YK�3ܞ�PVך�2 �*�&�C"&���f�M��Xu��T�F$ج��nuv	��ިos�Y�P�R�կC-D�~[��5Ϳ
O���sO�śF�E���7��7��R�����
֌*pٳ�5�W��֪����7>�h�nMۀ�'�*?��H�:mY�j�}��?����֋o�fm��؍��|D�=����<���w��c\���M�'7�s�\��W� �@~�W�O�{�~��Z�ڿu�s� � n���AxsD,�Nx��	H4�p�#V�A�Iz�c��G���e{�����v���Q��rOi��B
�L&�����&��l����%(Fi��C�%��ף�Ҕ(�^  #��(r��\�ܑb#4�2���y��	s�����{���a2�y^9{I�8l��r���FY�4_N�㕇^��De�/-���^}�s�
�$�u���\����z�_{d��-��T����9�PN��'���1
  yj�}[}H�uk�*�匝yl)v�(� KT즰X�1FC	$���U�Pq��*���|[l�ߓ����?���n8���Ű��\W���v1[�b4�$b4(���a�}��T�FzT`�" 7~f�?wL�?���O�}�qe�7_���c�]y�ewAEE�ֱO�p昂oL,��$�9��?�X������Q��ap���S����ml��q���v�~お��2��|ٚ��������R�����KNp;�_a^2�T.��l՞bR  U�IDAT��o �d|eKtKׄ�Aꤗ�n��(9��8,"sT����e�I�e� !�F�$K(�����Z�H��S�����&��'�dT��������:p�ߍ��4��h4vN"){��"�Y��D&�o�l��F	��V��HkG$Zo�+�KT��}5��  @jFX��2J�cpJ����e���fy`]-^5V�(c�D&�f�xʰ�V����9|�K��g���Y�֒���JeBq���w���1:�S�S�h{��j�<O�e2�����R�Π��9��?�U�/�{=  �ԫ7w����V��-�@�Z +_�ԵA�%*9��������DC!	���!	�u���������.}ȒԊb%]74 ��d�0��^!�~�{����:6�Lb�Z�d���d��5F	�Y:�Fi�%h�F�{U׶�J�	sr� ����c���Ӳ���pD���v��*�z�k2�TT�	������=uݬ1��5�����בc3��,�+�\'u-�'�<,�W��#��f�q����������W��,�؏.?}��;��w?4il^ޣGL+�k4d6�f����Y��� `��&��O���o��}��GtZ�b7D-:�Ĩ�=�ay�r`6E�}T�qT��m2t_ 7�)n�)�-6�Y����j#Q����n�	D�����*����JiD%��զ�Պ��`������9��*  ��Q������J�vM;�#�K�r��{��! ���r�)%�"�&Nr�-珑_>U%�j:C�h�S.;����9b�+�A�ە1�s��ZX2�%_9����9r�2FK����=u�Q  ��t�J�._ �}��f6����wYE&�r7�)[�Se%,�HH�:Z4��Q#�	c�C��D"j�,�
ս��������MZ+yQ,��X�hP`�cՍfuo���iPW,1�%��R�`E�W���z�f���kT�:±J��Q F��e�r��Yy�U���}Z{ፗ�~R�����[��-����/��5��^�5�kE�T��$V�=���.�~��1r���v�U��f͏�X��Bn���O�ݼ�y��œJ�W�vf��q�|�to�l�^�>  ��I�@H�_��J�<  �0s�\���B1�mהZ	��猒�=Q%[��Ou=:z�;�T/�	���r������+뷷	�e�^��\��"?8g���齲aG�`�N��/W�{������u��'���J�   @��Ԇ�R�����/������j�� j&M-������n�Rh3�����u����{��tDcű�����I�u @������%b5g��Ac[G��-{�k߾��+�#���k/>�o�����Z\�d�S��/��2[~��2�����|s�>f�����w��{��Na7^��V�����J=zF��Sf^����?�X.���#$     `�:��9�<Az8�&��Y���G+	�����Y��3Jc���F�}0N]�+������j��o�Q&�=UE�}��X�'�[V H��(�]].?}�R6�&�  �G�Օ�$���<  �u���Ii^NF����n���.?}��n���n��w=~�Q�K�+�w�2�ث�LR~�6��6w��(מ}xF?	�����͵����ޖ�������P��7c�K&wT�K�<m���ѷ     O'��n� 5�����r��{dgm� uK��	�g��d��N+�}�
��l�[�=�p{�Y����2���=|Xh����%ܞ�؇����?��5��    ��X�t�,>�4c�����~�o�{��W�q�e��x�/~f����O)���ǽ���yW�T7�Ȱ	�_r�,�T���cE�QymK���G���U����Z�=|����>����	�c2�'�+on�+�����B     @w�'8��	2#�j�Uɾ��]��ZX*&����	�g�U�,S��N�k檍��6�.�2F3F_}�2F��S����#~���Lqؔ����1��c�    ��_⑋O�����^��{ss���\���0�_��^�����{��Q�ح�u;mf���Er�}/H$*�5,��'˪��3�X���?�����/^u��`��**��k[���gf�>ݘ�����>_�o�'�-T�    `�(p�	efA��"��Dn{�J�:�|���(W�R�,��qٍ����Ç�H8� ��n��~V�F�h&ysLr�2Foyd��q�@}����hf�Lrթ%r�c��Q     �1f�A�]�H�fcFﭏ����޲�ƫW7���O�􆻞�˱3�-�ͱ���f�+�5˦��/m��}�]�!���yY$ml�<�ޮ�o�l՟RQaPK��q��<����/�Ŕ��s;,r効r�C�     .�l��o��� 1�r�q�<�nC� �?S,E^�O��&����������]|b�x��0}�CV,̕���kg���IŒ��>f�͑��y���6	     @&�=�0�\����zus���M'-؟U�n��̧����,�U���b�#ݏw��3�M�RY�&z��Ys�	U�J���4���oϩ#����Kg|7t��'����9�58v�(Y6�\^�\)     @ߖNu��1i�_C>T���q���ަ�v(�4�s�H���y�ڇ�R��6{\�,��ͦ�K
�Տ�d_sP�ۢI����=k���[ۤ�5$      �4��%7-��F��v���z���[������}r�/�8}t~A:�f1�7�\ ߺ�E]^-X��	%�X	�t�^��{������$t�WV���������aI�'�v�\y��j�X�    @�,f��wLZ�Ր��$k�̗���t�^��e�ʐH�l2�9G���O�tgT���
��jQ��Q�g�=�W���8���a3��er�?�      ���r�X-齒_(�����^t����n����_=31o�;�hT:k��"�̜1���]�7��_v�l1ӻ���-���=�n���M�>�xɪ?D�z��E��Lc%�"�C�9z�<��     ��Y�s�zji�8n�G�|�^�[)��I.]`d�.[d������LuIYcT�8�%��j�����;j�[
=A�9�-��V'�MTq     �qԌr�?�(���Vn�ݝ�n�_�U�6�]��D���m����t>�%'ϖ�7W�(�nW!�M/�E�K�������[�w�U��Su�e�����5+N�=�����ч����.Ս�     �E�Gp��\�>��OY�'��Op���z�V�?��\��3T�w��<�>���ϓ{�Y#��ܮX�/����i�kWl     �`6�+'�J��<�ޮ'�s��_�䑊��ѿxx��j�6�<ד��)��uY�Z�w�j�%�M�Ks{ ���=�n���Wr�WV�2灿���`�w�i�Ƴ�l�/�0Sn��     �e�8']u昙y��:	���qE6�Xb����.q�k���L.�Ǫ�C?��?��V|^GU�F9�<��z=Y6�->�O!�(     �֙K&��BWZ�ō��\��g
��k��{�|��f�<������(�_��&��}����8o��.H�K �g��~ɍ_=�i��|�����?�u��Z������1���[dgm�      �8j�[�/.�Q�ˑw?m0F��d2��).���fcT���,��71�:jz�
Ba�6�,���>j      �8�f��1S��o}\��f�IG��Uۿ{�Cǜ�`ҫ�.�)���V��������f�A�_>-���n��?U|���Cr�+>����-\8�xR:�W/���g�M�.     @�F����Q+dp�x
cT�'��^���魆��9��{L���:F	�     -�Z:Ir�����}�����/�����=���W�����^�r��{�FcZ�����/}$Ս�����p���o�m�;�����h�}���
�;���t���r_��5,|    �J���3s�C R�5K��"Пi�X%�p8*#YY�Ur�i)��!�>�+��CT���ig���e��@���1
     ��Vo?{ٔ������n�:��k���L-���3k��3��t�o6uVq��S��*�Nʭ9rr���iln�ްL��[����p��:b�c6���FeP�}���co     Ⱦ�	Q�U��,�^��4e$�>�1�WV�A&���J��d�G���c5����j:d$�6�1�W���ʷ�      �)ǉ''-��c��`ϝ7^��Y�f^���(�^W9{|Aq:�?y�X���7ICk��Hup_2�L����w0��l�}�O�:k�@S?����s��?~v������	s�����$��}     �ktA�&:1t����H��)LߥT1t�k�H��)`����B���:�o��(w     0T�W�� �[�?��O�B��G֮O����U�� ߭�e����x���ߛ%�tp?{Y�~X^�p�k7}����E۶_�Z��iS�rs��[����#&���(      ���-�*ϳ�>.�=�Q}+��C2�Q}+g�2Fu��Q     ��e3FIY�3-}7��#�ZO�ŭ_[��{�S�^�h�7����%��O/~$�`X�I7�1�.�3�(-}�k��>�ٶR�6��w=v��f�Q��OY8^~��&	E�     ���C�Mϊ�|
�<zV�e��\�W7�&Y��7�(     ���'���W���W��K�6߽茫'<���3��jݷ7�*G�(���g�[��Y���(Cz�~es��~���5�����O�=��7��^v��}�lr��rya�     ��j��vh����x��nM�$�0��7;���Q�c�    ��*�ˑy�S�zkUS��iW	�n�u�N)���b6i���E�	���&��8lZ�޼���{��N��w�=�roe�7G�S�#�    @���<�T=#�<ƨ�1F�1�s�g|Dlf^G�,��Q     0D+Mc*R�yo[�y7V"�������?�����9z��}ϝP$c�ܲ��E�E�%SKc%��F�]�	2�o�f����.���hJ���R��     �y&����H�h$��g|HF�<�6�ǨQ�뛌#�9�;3�!     `�\�	��S�����n�t�_�}�o����*w*w?g����&�]ܗ���~7l���K�m�\���wA�ǡ��R�ԏ�9J�              @�f�-�b�C�~C�����r� �~���5����玝5�D��>n��p�YLr��Ҵ��aU㵂�����ۧ�ᯏ�8o�Z��>v6w              ��:vVz
R��i�֛.?�eA�U5/j��r�̚^�ot�K&����U��Y�/>�TV�M;�ko�l�YѼ/piC�M�ˮ�e�O��R��               ��`9zf���F�Q����JAV��������o/;k�QZ�}�2^Fn�}JIZ��pO�����zUc��<s��1�iٯQy�=\3g�               �K�R�qh���u�n���
�foSۗ���Gv���E���_�$�p_���{e}k����K�U����E"����q'�              0 �KOA�O�#Ȫ�/[�u��޶`R�-��\�+n�Ե�%Ӳp�X�b���ټ��?����kk������WP�e�'��Ѡ^�B               Џ��4�S���1��n羦{L*�E�>��B���BQ���M,Ҽ�H4*��?����5��-�t;,�O�|T�(               H�b6ʌ�����yW���\zrP�u��c~^�⿩�m7i���	E#/�>sl��}~�����+׼.�����큫=9V����W@�              ��F��B�Z�����.�s���������勵�w�X�?��,ܵ�Ko�izB�W�m�ؿ>Z<�d����W(����                �t��Q����5dvu����se���}�*pI��&��IY�y�Mk��mw	t����e�m�=K�              Nf�!s����}����x����H�Ӧi��c
��͕�IY�O.�ռϪ�����8�M����wF�ѫ��f}���:m�Ԗ�O�               '�˴���k�xJ�+������?�x���N.󎜀��R��}�i�X�;7_�f��^�)t۵�w|�G�o�               ��[�؛�i��pD�C�	t�������@�>'�x$ӲpO�_v_��]�YۺyL�{��}N*%�              �������������^]#Н����y�]�����Z�}t�K�>�Z��
t����we�i�}L�[               �X:�{�[��ҍW�\���7�I�>�\b6%�H�d-�^���Ls{ r�Uk7	t��C�Uv�j�gi�S               �Xin��}���o	t���W_�qi՟� R�uHe}�dJV�n�E�6m����"Э͵/�a�Z4�@HZ^t              e��nD_�V}k�ne�Y�]��>��騼]���+ЭG*��t�+��6��TǑ� �
               z(�uh�_4����u�j��(��Z�Y��٢�Y	��95�8��l�ZCk�nt��k՟�l��Y�:B              ���]vM��k�n�ֹ���F�Tv�ײ�|���?Y	��s�������ZS{�Ne�Y�]�ɱp              H��qfw_��I�k�`�?Z��qh���KV��4TpB�t�#ޫu��U��               ��qٵ&����]�RݱQ�>=9# ��[4�3,F.w�s�`�Q�>3��              ���i����m��p�]�k�T�����bҬO�H��n��	��k��D���b6
               ��������6��u��ŤY�֖��w_�p75�8��oW	t-kp���              �dNC�2
�
t��=9V��٤}���Ǔ,���!u��]�uZ����              0�Y����Qi�^{ Rv���d� uV�&�+�G�Qy��"�@ע�日03��              ������e8,݋D�a-�3G@�=�hڟ�`���ϭ�zU�@��&s��}B���              B!m�*�����dԬz�*�~,�%+�t�%;��ReG�]��F)к�P8*               �.�����l�t�n5���/0��4|"�d6��-�2�!�3�              0�� ��h���0�u�=
K&e%���4�S�6t�l2�jݧ?��X              �ґ׵��N��٭&����:2���J����C�>QC�@�,�W�>�1�               �����C5��Y�6�)G�kW���|�Q�﹪�= ����{�/�y�v�q�@לV�x����              �p��H�ۮY^�%O�k��2��l	�tT�v;m3��粕iݧ��              ���B�Z܋s�Tp�9�ըy�}DTp���׼O��:N�k��G���:b��               @o��>�P�]|3�f6\��?Ϲ�k���f��u��8ʤ�ܫ�%���`Ь���P�[�����<�ͤe�{�               ��#k��1-Wv�u*7�6I�>�6�K&e%�
Gd_�_����T��W�[g�X�<$�S�w�A�4�2��              0��#k�[�V��V�u��.J�����J��jp�ZL���,���	tǛc[�u���Tp              H�*Y�����N��wO�G��Z������ɤ�ܷ�m���5�3/��y!�K�^�QZ����I               �X:���=��
_d��4�s{M�D��Q��W7k�gi~���TTD���)׺�O�j?�               {�Z�#-C�E^��{w<|ԏ�X��@W�<��Z�������Z�=�Ie��V�o��"�@7"eO��vL4j�g(��ʋ.               �D;+pO��i��N痔w�]���u��(jޟ�ܫ�$��Ԙ���tX͆����*��#Ѝ|��\���T�aQC�               Hnke����\�r��|�g��+v{��W?�����?�O����)�ؾ,�uel��8��ܰ}�               �ow��i�Oд�)��q�z�Sqթ�/�
,߱����E��=�iY��6��<�>cL��u��˗�YWq�GN*��j��Ɲ�              ��}��N�>������r�_][�>O�>7ﮗP8"��Հ�;�e����Y�q�M����rx� �
\����`�              �SY�&u-~)p�5�w|��!��<vش1y�Z��1�HEV��|R-���Q���肜˅��.6:����V�{�              @����FN�7V�>���+S�����H�U��Gf�Q�~���F�!��_P6望�c4�W�o�7���}�\�|g��z��<�U�~��Z-               H�Ukp����q�nR?'Ȫ)e��h�g{GH6���UjXY뀻�j6���V9\+Ț	�����7�              �L��F�"F����_��슇��T���⷏^<���Ժ�w?��P8"ِ����[�ʅ��м��
WW��⊵�����7��8wb�8��m�e�v
�              ����U�=Nۢ�%�9����?yD�jAV�_xK:�}uK�dK��W5���[�ִ�B���r��F9�P�qFy�04����ō�Y�4              �p���4��f�/���"�͊
����??mt^����"Qyi���^ظG�?n���ΟXt��~�̥����A�\�cK�M(������`�               ``^�X)W��'F���-t;֏}���5mT��i(H����X��l�E�}݆�i	���X�xj�^*Ș�ŞߙMF��mjȻ��               ���/�?�����5�{���oV�[wS���!AF�p��g��_�����!��up�^�,�w���1����tZ��߻㉛tř�i��;�`��������ww�.y               ����;;�p_�u~�Ύ���iWQ5����4Too���H6�"���[��p�uڌ�s�R�Ҫb�:������aQ=��v     �
t.�8@8V !=�S� cT�ᨘ��Q�
�G�U_B��QcT���      ŋ�*���êy�GN/�B�=��Rq��i���{+�MG��zo�t��0����Z���Sf��nѼ�#��λ���ι���	�ƹ����u���v�Ɏ�f     ٣��p��L�M�|Bo�@X\v�@���s�E7S����0*N��z���a     �����;e���5����z�T��滿}t�i������ �nf�}����i��Q+�/�R|Oźu�X�<$�ܵ���e�K?����     �����l�S{�2���t���pl��::���U?���A!��B     @O�񩜹tR,_��������'��KV�+H��Ş��KZ&�6��'[+%�tpW����e�Ii�����{�]�(�'	4UQ5N���:��7��oC���q�     ��m
�7���^�4e��i
��B�/�
m�4Q�V��y�_�ڨi�uT}�/t�j�q�     @���ʫ[�d��r��VC�GM/��;�z�o?���M������������>=��eucg���٣���1�F�������w/:���ɛ���f�]��������%�    @�U�er�]�O{�U)cT&	tjoC��t{�1:w�@�*2�U�d�h�@�*y�     y䥏�pW��X��E9+��w~���������zԲ��U^�R%z�����?�cg��t<��B�N+����}��7u퇂!���ǿ|����꿱�C���v     ���N����k�̝�P��Nƨ�c����<z���9     ��;�)[��W����L(s�����o~a�y�!���~���ʟ���ғnW���%�GAj�ܷV6ʋ���13G���|��4g|ɋ�֕W,_��p���w?4i��Qw��ƴ=Ɵ^�P���      }ؼ�'Ч���Ե2ݵicT���^M0s�.�@���ò��p�&��u��5��Z     �����&�ŗ�N[���u�w?�č��|D0$Kf�Z7���IW����ʳ����]�]��o��f��*����1�EMV���J���ΙP�v�ב�1T�◧��&     @?��tH�?,N�I�/�;5����> ��V��lQ�hD�_���)(���R��EvG���P��4��{��l��.      ZZ��V���F�O*NK�V�I��S�'�o�U�ճ^�O���#��.I�c�����$�.�۫����w�	�Ƥ�1�L-����y��z�`@ήx�z�伍Sʼ�t>���� ��    �5����mrܬ��� ��Q���[���#���k�����Ey}y�1��׿��EN��+���    @:��_����%M5�%�e71��?߿���7_z�'����'+N^0�2C��A�m�Ͳ��]�'�����̮�N��/��If�{�%�$���Z�RPauW_�(�e�(AX\��R�f@B�&�!!!���3��{�eqeW�����|>��ɄDN����s���N��䷸w/n�!�{��]w׵g|��/o������޻ޒ��.r�g�    ����r�{b�V4��U6�����eq�?�|��w���9��2x͓���k�YK���������1�,7�   ��7�xx��]J=r`�nF�xƅ�����Olޖs��������-���e����X��7���MO,�/~dB��#���#������~�}�o钛�v�C�i����RR�:    �ۂ�ձzs]�`Cv*�S�J�o���+�9?�$H��Wʣ��)xͪ�s袵51vX� O�\u�H_�d]m,]_����܌6x   ZHk,��mh��5�L�t��I���Vuo�+n=�#���}��M���_�/Nd���i�w�a�z��9�������^s����/����]�w}h�!�=������U1���,   �k��#�xnk|��!A��6c?0{{�FSgl�'"�����o4�٭qƉÂ��E��������k�7�������3
   ��l)���_��-z�	;�ܥ�ˊ��v�^�������W��gԕ�J�[tu{]CS\vϜHQҁ{���h�q��ע�.,(�c��K�o�gط��c�7�t��5ŏ�=d�Н[�\���{^
    mO/����C�m�Yۢ��1x�9˫l�NĴ������ы�*c���u��m��e���!x��+�w�-m��9e���k=   в����x��#b��-z��#��+-.\��7�'�⛧��༫�������'݊Zn���{x^��Z)J:pϼ�dc<0ky|���m��t��g��WN���5���t����9����ߥ��v0�5�w�}s�W   iklj�k������l�h�;f����\���s>3*
Zt�	o���)&O��o��0�~xC���Q-���7WY��<eF��lF����Y'�4�mh{Uc���   Z^��ϯ��|��_}���JK���b�%�}��'?���.�����-�niK�m�[�/�T%�g.�oN8fp���>t��}_Z�q��_r�a�q��,�N�Ko;�	C��ثU�\�zuC�3si    �C�!�مq��=�����6EM}S�-]_��߯e������ͱ��.��gɺ�xtnY|h��A۸�����&^Y]����&�
��Ol��Z��   @�X�jk>z>刱-~�A}J�>v�n^y��~��/�N����~Ȅ�6n�?ti�m�M��۞����HU��˪�����?x��_�>�>|@�Ž������z�U�	���ר/�V�*{Y*j��S^�o�   ڏ����=�[�]�����s�*�7wӓ�c܈��yP��u���2��=xs�?�17��cx��u�X\�.��]���=,7���ַ�gT����   К�~��8`��3�����Q\p�!�]8t���}jޚC���Ś�d���;������&�k���l�����=���q�S�Ƨ�*�ػ����w������m���M�ԥS�ǘ��)}��(},�dߚ����Y�a[U    �KeMS\z�8�Sãk�V�N��k�G7o���9.�g}��QQRlF[˦���Z�������O?=*���ֲ~{}\u���ew
��=���E�f����RW=hF  ��W��?��\\��E���-~�lcy֬�[�v�eS?����0+:����sď{���/-���-�Ե��=����޻�=F�k��u-��g����=��'����sN?����ιjʷ�}�����l�uVw�X��Y   @��pMu����q��C����m�h���Xu��+�/�cM|��Q�B�WQ�ܶ&�#o��Mٌ���8��B���:�<:eMTՙѷk�������;��vB��V�LY���    �-��X���R��	���9���wh�3{]{��Uˎ�ZG^L}�巎�uP�;&�2�K+~����6~>yF4�����U��]r�����}8�����Z'��?p�}9����W~�3?ѡVf��?o�g���M9`��ݺ����Wn�=	�   �}{fAE�*���� �{*�j��o[���wf����F�o=D�ق�k��?���_T�;3wEU\���8��!aD[NenF9%7�[�wf֒ʸ����Z߂^�Hhul*3�   @ۺ���1nD�8�]Z휽J�
�>p��,6픳.���=퓷F2iRsA�.w_vĄ�_��[[�܍M�񳛟�Me5����=�q{u���/��U��/,(��a���U���z��t����w��+)�����Tڭ��+���6~zӳ�   �����GUMS|��C��Uߒ�6no�����[����3+��ා%���m{Uc\x��X��6xw��R��M����B3��e[��{]�ь�[��-�=�6���RdFw�����gwu    H�o�����=F�k��޷��C��2�O���pS���v��h�~|����?f�e�ٹg[�������e���hw�{f֒��܃����m�s�SRt�������i��«��׿��[N9�1ڑ�\O�L��3�������7��o,�   ����̲��8��!ѫ�k�c�_U��{]> �ɶd��ϫ�[�����ۣIZ��6~}׺ذ�����W+s3�&N?vH�iFw�W��įsϣ����\\��ڌ��aFw��k^{��R�   HG���ᙸ��#c`��z��n��O~����w���+�U~�?�8e^�3�]s��F�y�����ui�[#�?kE�:}q�'����)ϼ����O6�Mο��>���۫7W�:�ڻ�0o��o];�I��?�������}G���=���'�����B�]�9   ��g�����+�G��#K�w��9b�-q��[�_�cd��nX_���8pt������{h�����M��hHw�,t��������W3�^d3z߬mqӴ��hFw����s��+��G��w.޽lF�z~[�2}s�6�    ����i�}0ztk�츴[a���Ě�/�1���K�V}��o��|$������C��d��i�?�����_�������C�����ٟaĀ��s�W3�K����u���=��O���4���`��SG��y��;�{ri�{��������v�   �Md�G~��8b|�����ޥ���SK���5�l�%�j����1.�cm�[����^����6�fk}\���l+>;^yuc\t�k3��#�����|cm\�Ȧ��x�]Eοm�k3��A�8�.,]���G7��I�O   �e��ܛ���}�(,h��{qa:~���m�����^�������M:픊H�/������~:vdߏ�4�W�o����~|������M�~����9Ν<#~�����1����2�OI���<<���V�xmٽ��T�{޷?�R[�y~r��c�.>s�Q�6���H��O.�   @Ǘm$}r^y���2>��8j�>ѣ������T�?�%f,��iY�r�9oeU|d�>q́}�o�v��i�X��>�xnkL�_n�p+�ft����h�9����`�mX��.?��s3jD[^6��������7�޿O�*1�oe���Z�^�   h?f,Z�:3~p��(h�U�E�]c�]��?(�����[��zK�%s��^wˤS�Z���o��>jpi���:��?��`A�6�C��zsE|��iQY��Q������)~|������20R���>=s�ɹ/O�ȴ�K7�-ް��ʆ���=�S�Z��U��u�?�������c��>3��%q��s   �\*k�⶧�Ľ�o�����������J"����PW�3_��'�ŜUb�VV�������x`��8t����b��R3�W�cֲ��.Z�ͪh�u��7ŝ�m��gm�����#���q#<��������,��<ں�k�b�[���f�W~F��݌���܌f�M�����(   �>=���(*,�3N: R�{����}r_^yL}������[*��\^{c�u'�8iR����;O�߯w�{�7�σG�ӿ�kA�dcYu|��i�����90��ݨ�o̯�?�s��^;���SR�;�������#{�vsYu��+r���U���64>��[ɲ+�v����wү���)�ۣ���K���YR<�_��Q����M1h�kw�\��5;   �Ϋ��9zi{�ػ(�ک$�U����Fׂ�#��d�j�ax�ژ��*��9�g��,�}b^y��ۣk�siL��蘡�bH���ڵ��hb�ݚ�hM�[Q/���_�B���^�[�?���{e3:�4F�ftp��(L�3��]��f��U�9��3�m-�`��9e�����{���k}I�64{��\3�}/�����h6����    �w���<����	m8�^Ե˸���玣s?=��z�u{�����k˫�U��=__W0��8��OX�f��I����yt��.{�ҳ{�޽K�wЫd�~����Tm�^g^�d��Z�Y�Q�;QYS߻nZ��_�F�e�zv��s?͎CrǗ_��Sg��u�͵��Uu���CqQ��®��
���U'�N_����m$   �_l*����fGY��Y�6�OQ�v�%�Qڭcp���E�5�QV��+��� ;�m���M�ّ�.�ػ0z�׌��f�}�]�7eٳ�*w�U5�g��yi�R�O�\�?2ٌf���1g�17�5u���^�[��h겿��_.���>��{t/��E�;��g4{��^ݘ��   �4����O��/�URT�kD�~�/�cB�8��_�̜9QQS�\S��T���P���Xڭ����k�nE݋��~��ެ�\g^3-�ok�q{�������OǏO����MvEG���E�u�{�=2?��;    �LCSĚ�����R������z3J��]�y��e��ٝ!    ���"j���:(����zv/�;�U��c��/��];-6��DGС�L]}c�}�3�c������Ô���b�*          :��箊�۫���}J���1k��8��������U����v���5;�l����wtI��TU�򳛟���          Ӽ�[����_|��9�gк".��|4d�t�!������X��<~x�?D������T�nz&��/          :�l!��^�X���1q쐠�565���7?�0:��g�-�_������c�������5q��3;�-          xseUu�?L�:b�������.]���=���ٟfĬW7DG���̆mU��?��o{�.��UW�W=07�<�j4w�;          �6di�Q|ن���'�>�������q��g�����:E����o��o!��[g�t@���=x�o(��n���n          :�g��/���8��!{޻����W⏏�M�`u�	�_7c�8�w��7��/��0<xws�[�/������          �m��q��O��w��|l��ѽ(xw��My!����E��3�Z��o|&7,����Š�%�ۗmk���Y�          �O٢�;f,����������sD����7����-������:e����_Ys�m��9.N<tLt	��������yqg�ɦ�=P          x���?���8|��8��cx���{l���9�~[UtF�:p�T���e�Ή��[���ǰ�����g������          �D��}Ƣu��C��?`��ѽ(x�Ek�ťwώ9�7Gg���׭�T?���1aT���G���w�]Sss<�����cU��          �V}CS���¸{��ġ�㓇����X7=� zqE45G�'p���g\�d>p����~�0t�6�?�Ҫ������          v��꺸��1��%������k�v�|Y�eq��⑗V�S��7	oӬ%�ǘa}�S���#��]�#��m��^X�L_�U          ��m��q��s��̏��%N>lL�[�����Y�6t�����-,^�-οuf\u����~;űw���{DG�pͶ�kƒxtΪ|�          �%�Wo{jq�����o��q��]�	ãkZN]QS��]S�y5^]�=���o�������-�=pŇ����*)��h���|��Ћ+b���          �����«�Ǡ>%����kD��7ڣ��Ƙ�h}<��ʘ��ڨoh
ޚ��jjn���?����w�s��-Y�=� �6oM��j�[          ���۫���䏑z����>4&�4 R^�^^]�/�O��6���vz���{����,X�?2�����20��=x���֦�5[*c����Ҳ��ܢ����&          �=Y���/�{���8`���w�A���b�!���K��Y�>喘�bs�\�>������D�-�P�?n��8���j�=F��݆��Y �[�s���[+�յ�b���X��,��[��          t��������#ӣ[a�5 ����C{�N{EQa�?����|��tCY�ǅ����]A��%poA��"�����g�E]ch��گG�S���޻�(z�v�n�_ˮ*���®�����M�M��u��+<ʪjc{U]l����۫c���TV���         �3��m������e��*���JcH���׳[�)��K��WIq��-.,���.�=�uu]�k�����khʷ�Y�����WǺ���~[U��iy�VVW�+6��          `�jn���옻|sо�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          HBᆩgw	    h'.���v����HPCCC����ۃN/7�����"=��8㌱A�w�E}?��/"=r3:.��rϣ�rϣgGb���g�y�    h16�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��۵c   �A����Q-�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,,�ъ\�    IEND�B`�PK
     ˡ�Z����C   C   /   images/ba153158-cccd-4fb1-9320-38bebad1b7f9.png�PNG

   IHDR   d   4   |l��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��|yx����=[2�=dOHB6H���Ȧ�
����R��jk{�t���zi۷������R�*b�V@TY!@����=��d��=�L&$di����I~�[���g��9Ϡ�Y�����b�x�Ǉ���'NwC�R�j.�s��u�B��Z�?q�'-jJj��c��c¡�v9�v�w,��G�O{5:L�	}xߋ�mgI34�o��RB��h-��%C����v��:as�q5��Q89O�2{{Z|؟����,{r��
�:6B�U������B̞1}�������N���*�Z��Mya�������\.}2��Á��V��P+ZL�o5M`�����3�)++3(o۾� ={�ɖ�j,tOrL�_�:��E�]�����������S�qy��Mʰ:7�-Σ	��my.�cA�	Ĭ��Q�Oar�e^�3<C��Y�e��w���k�5|���Pw-��X�'V翐�����mGOgZ�.��e����@�� B�@t�Q�֪eR6��f�賸au)}~\���e��^\���RM�����FNz2�:��i'���G���E+�AH �F�9D��59�X��5;e��DJ�V*����8~z�ɷ&'�{%8P�����V6w@�V*���j4t<5!6�ʖ^�4t�	Wx\HU� c�MN����H��BhH04�h��h�Z��׏��v�jơ�N�t�`�0|=0,�H�����c0(*�I�t@���p{!���1==�s�0-k<�b���@Q@���fC���ӭ�8^݂/��Q�a�٥5�"96�/k���7O�}s[��*��,�AV豿��������7�"�X[�������i!��T�wAI㓑7m*V,�A�ށ�GK�i%���p��Ac������D�.h�k�W�I����~�(��f�c�iț<������zss�`�utuu�HI����k���U���� �m���Q�D������*�
n��Wb�j�3�
��	hii��`�
!�������T���a���������CxsW��c��'�e�A�ų"`�*Fŧ�jZpOON�����W"V>/y�%!xx��#8�h)���D{{;��܌��^!:�����0aRRRI�187%%a��|��{��8��.�O��9��zΚ��-�I6���+������������ݻ�u�V�<yR�Ɏ�d�J�PZHFF�.]�U�V!++	I����k�?�8�����e�U�5Rg�w7Y�ƣ��	�"'#���?�>���
M&�yY�F�҅�����~I��r~pЌ#G�࣏>�W_}%��K��S	�������E��zsss1.:wݴy�����wa{�����I�ya0R¼x��B,_�� X�"�oߎW_}� 5�e��F=:G��Y,�8q���X�~=��<��Cb=�����"�����r�Pغ�f^��һ1))ڀK�C����}&|Yg@u�Opc#X��S7��{�,CHX�X;�?�	��n���3�*��+��y}�x���
Q�w�yG@�я~���Lg*��X$��ފGڅ���9���T<YƳ�Q��Y"q�������q�F�8�d�PrK� MVE���dF?i�iP����_��_�w���ϟ�I�&�?P��ڇ�]k�83g-2���Rf���$���g)�C.L�g�ñ�%y�B4�9ߣvS�䖟X���X)q�l6�7���/��Ʉ Zg�&�ؙ��
^/���t�J�`��[��o�>��7��ʕ+����_~�k�-��q6&�&�f���ibFSS~������iub��� L�LG�����F&Ǉ�h���@{[�O���|�V�Eyy9x����X�b2H{��ף�孨��H�c0��`4ۄy�"#)
��:8u�A+ٍ͋9�0c�x�t�CK|>6"�m��n��¼t4wP\݊�-2�G�����߂x�n�Y8��r��100�g�y���D��`�൦f�#�,��(��C`��Bz��q���vY�^�Ǐ�cqs=� b���Խˡ7��%6ӛ
�(f\+��������i30uz��G1�?%��9-@�]\,�f��T)�ع��� �F#�q����Ǵi����v<��ð�Ւf���z�"��ff�AO���!� ���us�VbޔT��eAv2��}�
'cJZJj�x`�l�,vܺx�\s��E��?�Q���o]���q��>��h7��C��&�!o�L�Q�~v��1�x ���D\�R���܂S�J`"p���{N�����GJ�<~�BԾ����HLF��G*��U� <"2;v/~0xL��M$���?�ȄU�O9����Y�/Qdm�������(!�_�BX���������n�K�Y�y�t2o/lD���l�l[��SR����퇫�EI
rRĪq�dQZa0�SSq����Z�;<XK�ha�9d^��5��ƙ4�	���� Afdgaz�,YӅT�����dM�QQ(:p]�bM,K&9�/F��<ܽ��o�aG|�y�z�Ǎ��fbJN���mۆM�6[��=u
M�-�����u ��i���iBPp%N��I#<����7^}�>�P��^HB(������=�P0W�jw���G���0g��N
�UL{�	�����ാs&���6��d塺@Y���:|t����Š�!�E����)QX4o�ģS�Nᥗ^b�H����s|5�`��
�u�'H�3���%2��x!����=��)S� �<����`��F�u��s�a@8�'�����>�'6,(�C�I���IS'K��+X�J�H۬V�\32�
$���<AC~ۋd���q;�|��K��c�	|7�p�fcav�QL�B};�,Y�6�-���pk5h�6�bs�����(�m��RJ�0�,�&�<��M[(����u�`�,C���f�x1��^{}}}$�-��ř��ȝn�:���!�ޡШ��{Y�V���B��OwJLe��Ĉ�����3SQ�I�0À���ɈFf��{׮]�Y[8�O�1]bSvO+�&8�%��vv��7�L>�4-��$��T,�����g���Ѽ6��P޲���֓� ���LEc��fsbDPf+9R�$����Ҙ���51|o߀e�^!I:̜�-��4~�Ν�r)S��|!*~ː�@8]kHl!�TС$r��x�?b\$&Q��x�����vYI�����{��c�Q}���B�<2����l��ux|�NԖՊ���\��`�X�� �W�J@#Ka��Қ3o.N/����~]]�$Ry�iH
/BC����$^�)J���tW94'���G�+Z׬�����?���az�������n��p�.X��;�e����jQ���Z	�LKANB�֛I�J l�Q:%rғ��B�؟2�<A~�
[�m�B�g���_�j����3y���db$��u��=zT ���AV\��p�5��C�ʃ܌DZ_ �/��R\1��#צ䎥�u1��3� �:>�aוH�My�S�$�˗/��w���}>�bB4�����\��:O��:�؂�'Iʔ��-�27���ޞ^�EF�ű��H21���Zy?+ ��MYc�WjpHP"5!F��K�O�<)w`e.���\�^��5)\^���K�Gme����Sl���'FQ���k��R�@}ȣ��U\	�I����Sc�p�e�����5(�
����v��V�K<A.Nr�NK~;n\���Tx�еJD���ߜk��b�j��Q��� W
�m���?}����}��a �{�A�/TK=����%�`���ݗ��QA���6��5�`.E(����X	t�@J��[׉����!-�r�w�}�af5�!����u��Ā��:8V���rrhw�`YBۆ�����-�@��O�Juق��:���pY��D����|_�0z� p9}�Kz��{����0 V
B,,h�����5ea-%��;i�<h|��XK�W�9�:����؛�{����8씧8�\���������/!��'��i�)��}���X9q1��N�P_�jw�)��Ff�qXOLL���o0צ���M�R��C��;)	�Sk~'�D�tW��p|%��D����c6L}�UV�v��a�U�*�4�r��^�N�db�M.ޚ-�=Oo�	z>��D��ϻMNt�(�NEzz:"�]q,��%ם8��=�)����b�F��Q¦PKi�=�շ����p�qM�,\��O6�=h�����ڒ(q�0V�F~���+>�
	̸��� ��2q����;?��w�."8��}p�)��B��Yݨi�cf�4����P6�EEF���q��#�&�G�'�����)��mX`���K��]�b���={�\�Mϭ�0�J��݃�is)P~�+Ic�����L���66 ��U��O%�����
�`W�J����A��FC*�{x����%��l�����cٲeؿ��.q.\ ~����,#-3�Cp�|��٘��.�x�:�a�:�;l�-s� ;;��@Em#�\���"�c�� &6Nji����F�]u8y	�q|��[Ɍ�uaP���rD��$���5��g���Ȁ�hjmC��$uAëf����Pd�p����E*��z=v~�V�^��d)D�R3ӥc&�+Ŷ��S���N>��gS���r
g����K��j1c��Z��\Y<�&V�6���:,��EAA�Ν+JȊT^r
�/
���J�Z��ű�<W9X�آ��J��bs��Sb�L�V�^����1v��
mnz�Y�E��6�����Id��3�>� ~��_I�ݻ{�⑛7��Cu����}Z#�`4�IBg�Х�D����<!+e��Ipsб`��N���{�;G5�.u\l�$nڦ�����;3O�G��?���Ue����c�C�x).(�P�������ix,�_�B+[���>�2��6l/��-QC���C��6��wO#3+w�y����U�-��$�͞�#����W��9Fh�>6�4�Y��Ox���C�슷�<���B���Al�u�F�9E�1�s=�� V�E�z��'۱�D��?Gv��{��K�PY�I!.ܐ��s"t.~��G^/ˢ��hnh����~&ۣ�7>���hTg��(��M��N6l;���(�췿���5������o���� �����~�Q�P=�'�A���ȧ)~�q�z֬Y"ރG����U4g��gh���k��i�F������T7wK�W��C���h7+�����JCTL,�|�I���ٳG@9q�X����dS��!~|p:QT���&���>�(n��f�7����]�{U���O� ��=Ԅ�̃X{�R��*6皚i��۵ՕU�6#_�V���=C�Tu�:�(^�46����@��׿���.�����K���::v�ă�CT��6�GZ�	Q����'���'�s��[��C� k�	ύ[�g��rf|�?�{�R���?����,�RGk�loGVN��Wt�[T@�(���O���N6=�e0�������\<����l�C��<��[������,B\T8
��A^^�~�mq/���İ�(���>��01��p�0P�����8@ԸG,�����yO[�ڵk��v=^ܰ���"�Q�F��I��w
{,r���zS'QgàPU7�E�E�D�t��}=s/2T�%��9<\�4�����<��|V��ؽX�l)�������f�͛7����?�*O�b%u�Q�E����k��$����o�y��`��!�¥eЄ�l܁��]R�:{��e�u��y����4�ysfc�ĉX�n� ��[o�����4�Y1BQFm��I�֬Y�'�xBr�yԞ_�16��WFvC\�	"vc���[G��99�������ơ��$J %%�|�ь� -��c��/�)��{_ɽ7^����b)LO�Cp��˙<����ԐG�[��pn�.�c�op��u?�+;��R��A�%��_�T�O��9�6�K
%���?�Nז-[�^__/%��2È�[/��-K���1�PQQ����������B�������;��/��~�_����za�!.2f��p�NO�����X	yK��y�K���ݶ�Z��p�s�=���k����QUU%���lο^�e����[n�E�8qŃ�b�{}�gX��	6������l�A�����QZ���+"%5E��2[`Z����R<�dq��� צ�<����38�I�~v(�+[�q���ۊ:ƻ���Ĩ0vj�x^;opX<=Av��� ��w�fwbRJ�����A��]a,���a��M�J�U�g6�@9=��51ib��0�w�}����K����if%c�c�p	�����j���'��������_���a@������_5�l��48�x���+����9�v�t$%&H �5�_$���|�� ��t�xi%���>/�ɥ�(z[�ԉ)�@	[��9��e��_Cy��ٽ���k �}/r)��˚?Nb̠��[�җ������݂�da�5��?$#<<LX!���-eT]�<��4�ʚz|��m�~з�y�9��^8�zd�λ��b�hQ!8�a��`��|/=�X�D�{%��]�ES1wj2SE����el#�V}'J���T3�6a�+d��X��c�E�/˛�*\�m%Ƽ�dG��J�|qEjE�r�d���dF�]�p��ε���PX9�����wV���X89��i������Hى��N�fqb�lFGW�j�e7塚��<�Ϯ<��c�u�J�@g���>���|7?����#!2hgC����R<�X]�(Px��0<���r���F\�I�:y8o�d����g���`���@�����[�NKV#9�E��`�-=�PJ��`j��A%v�:�r<�	� .�W<�8�M\���fŹ1>�Lא�����o�i��&��A��V��e��w�8�#tDE��0�[o���n�[j��x��Mf�iSR���-�NLJ���k��yǩ�>:� uTh �Z4���`Ɗ���<K�y��w�ԩ��D����~��a㲒��v��>3M|P�r�eu e�
�����H*q��Eh������]]������J5���Պ�+gG��Iy#=6 �fD�q?]�U	8F�ێ���]|%YV*&�����h����[���/?����K�&N�uw,�ؿ|IMs�|�����������j��AZM�[[v{fg���{7��o �H�_��,�T(��v����C�!\��\�s�s,a0�w��3x�3�Yj�(R~�C��/������"|H;[��7����gz�� 3;X�_��܇c#?i��~�����m�o����H+I�3�B�:m"�v����T+�7�"W��T�Y�(��}��A2��6#5bQ���+�g�صٝ�-mM��]��ܜ�����`���5��&���ge��>����-eM=A��4{�+�D���9{&��Ӷ�4J��:<^���N;~��YAnS�pzݬ��%>�ʀ�NE�t���*��m�C�V���xlN�W��f����֣�)�u=1##�a
A[�N�?q�&�+f�5��A�/��z=Qĸ�o~c���m�OuSN��F�w˺"˟c�U����������[�m�[�Z��
u��m}�0�@�b�k_Y��)5d8y�Փ�w�=/�s��~l�R��dl$��q7�G�����M��/�&D�vI�T���Q��؊�E��	
E��A�۫�X���w2�f��3m����h$P��� H�4��e�+K�.yF�sq�6�i���kv��q5���qa�e�;m�>zW����/3tJ����UM�Uc��s����+�A�fqZ ���tKcZ� 5 |���MF���P���__�%��q��ߎK�r��o��Ʒ�\e�[@�����lS��?�    IEND�B`�PK
     ˡ�ZM8��! �! /   images/53de2a41-b288-4dfc-9a43-3e5c75810bf2.png�PNG

   IHDR  @  @   !��   gAMA  ���a   	pHYs    ��~�  ��IDATx�����l�u���}�~/g8C���H��%Z����l+J���@����Ć H [�-+	Y�ș9�}��/���U���3g��d)���F��ҽ/�ww�UkU         6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!        6�        �         `sH�        ��!    ��g~�[?��9�]���4m�R����g�a����.�E�A㻞�r	_�]�����?����p�M��j;�`[�?�3�������&|�ȟ����>�	o����#��Ǻk_p|����C>�Q������t�M�����  ��	    ������ßYRb�X��|>�w��ہ��6�y�	נ�5H�߆i�(V>?�[7���׼/_z����g�ß�����������\~���s��}h�K\��мZ�t��yh�Є�ed��B��nd���F4Kh��Xsy�q��Y(���ބ�n�{���c���܆�?��.��y���	���2�F��*�g�m����N3���͑���]�!|����ܥ>J����c��_|�ٛw����S�o[���㰴ehm���x���[�0��u��>?�!�����o�Ϳ?���W�Cx���6�q���N��_�/��K��軿�;�W  �/	    ������/�tӧWs��0�B|LS�&h��; oGj���{����
@+8��@�5 ;/�wHVފ���\��c����b�6�3������u��wuC,�n?���K���|�};pܼ�滵�Ek���K�������n�iI.|�1�ϗ����[?���휏[ۥ��v1�q�����c���v��zr����}��q���kB���¨��|�yMl����NɎ��Ң������g9]=��4�������R~P�Ѥp?��i<��ǘ�\׆��4M~�r��K����awݗ�g�3����㘏Q߄��Q�f����]�mL� �M9i�vܻ��7�mПK�]���51��3��o���5;n�=VҾ�}n�X���~s��8]�ol���K�&��|���4Z�ܕdO�:�Ӷ�C�aֱ>����mc��\ئ��9�-���3}/�]���g�o�_���0��z=�&���w>"��k��w�����_  ��   ���G���fwqn��M�vѢ7��ܹ��2>���5��RZX|�|�w|��G�?�����?�le�����[_��qݚ�[;�>K߿��=���o~����?9^�����������>��c��n����������s_./v�n��mN����p��>x_�㏿wۭ��\��y�g�����n���o�����9���n���|���et��(-\>��z�<??�_{x��H�B5>�?���3�_0&�豂gB\�KK�.���|5���І��]�����y'�7���]�R
�rZ#��?��-����]��ϋ�Ɨ��}wþ<\٦e��}���E��5	����+3�/O�,�?Fӕ�����l�&ty�N'ߗ�b�|T�@t7\��z�e�����g��ŷb��p[���ڜ�j�q��Z��\)�Y�f�W�{��e����7�I��v����Jc�%���Ǵcg�)&?tC�����K�}��0����O�d�t;>��تFb�}>z@�vؤ��%����>�
�wy���|�:Jj(���D�B���������&�����A-���������h������m"c��c��y:�J�&�_�|�|<��I����9/O��L���;]7؁�����qCjnx>>��`�6z�E��3us��|MђY��:�ۭ��Y�%��jbdI����e��F��]��<�	�p�դ���oz%0��]���̢2cz��sƼ�M�ʋY����M����1R>�u����ޒ�[
5ϳ,K��nL�r��������������q�O��������%ƻ��W?���?��{  �/	  6�?��o}m���UJ��G�����o���\è/Z��;hyym����n�ߢ��F7}#��_���W���o�������my����e�^���t��/���꾍m34�r���U7�C���F�����yK���°�̧q��Q�S�?k�Ì/�Ubr!�G������5�8��]�0��]8<��������v��qm�Җ��i|�b��{ �u�o>F�ͻ�g���jV�r�L�}���<������ӯ_��2[�͛Cy�c8��s>�����f���{���,�ە��o+�B|[m���ُE�zp�9'�4�R�������;v�x[�V��G�4��j����7��v��cu�r8�}s�a�Θ�n�����vFu�B]��>�\�4�����u����?���<���~y��1��G즂@��|��u�Y@SN��0�Ckw��]�D��/�T�x�{�X�M=ȷm���u�Yk U�����S��yY�%�=��K!��Ƙ>�)|%���bl�%ͭfiǷ#����ԆTIGZA���������r��7[�����"�U��S>����.gh�ώ�~�r`����x���P8������3�-�Z��u�g�/�s���������������{g�i�.\�]�?ׅI���o󔿧����߇�~|�3�����������Q����������t���k��&��&F��h�J"I��`��qVH<���c>�÷˯�C>Vyh�M��G��w^|;������l���O�<<?mV���;O0�����l}�"��r0]�|��Fl�i�J��T2�Zd��A�
}��j���/v�������J�M�d������]�M����uSy�1�q5_|[�z��MQ�LcjT�B��<����D��Ul��{��ksm޷x��b=oS�P��9��5�$���:�U����ץ%��To.��NcV���#�����|�^�J�v���b�咏�1�����m:.��K��D�f�r(�ו�`��1�qnc�z�?��4m_�6��%�a��zqF��~龪�d�%��D��p��v��y}�[�t~��t��ޔ.�������_���t�,ݿ��o�6-�  �H�  �S��?��f��/"�����M����ҙ_��7��)�����,6cx^�}�8�*j�h
�����ω`���-C���V��uԀ���x�[]i�r�\�\�/#�
L�7��wf^L��Y�����#������n������{���?����_�޿
?�sߴ��t	��6,Gz�T��&��[��(|��Cށ�i�mH�.�1������i�T��a��`*�a3b���h��������u�p-�x9��6Hy{&��ø�8����9�al��P�]rnGF���4�	�M_�q��t���}��k��[�m�&X��ְ��$����g{'pu\���>����N�b{j1���|�>��������#�y�&�<�?���|��N�C�\�����c�r�<�p�n�>�휏���t}[n�źt����˷ۚխY�?���aׇeN��|�?��ã��5��n�_>Yc�[o����`��nn�k_��6�_j�=X�rݘ�\��WI�z	j;��������Z<�c����g{�������s	7>��w\��}\�
"��m������y������vt*��h�֘�AI��|
�y)�v`ݾ�����Pk���_��b�Y]�-`�0��N�"h��N�3�o)@|9_,�����=~x���M��/O������W{u�x?���JM�k^z�Z�|�\��t��ֱ�{Q�@���6��Dv��^j��֕���!�����-q�X�������v��Q�V�4���R�#y-�V��K3,���֪v��el���:�x:_�,���&j|���Ƀ���Y2@�vm��%�垫��VB��:O��j��{�7q�ӫD��E�$�f�����v��6�W���a�w��:���Z �Z�c��S��hv��~e�I��Z%>�-Hs�F��o㲶�REL
ޮI9����|_R� ͓��MWR6�+��i�ƯS݋��R*� �JY�|���Z������p.姧�Z�Q�v������%����g�^�Yt�Ә����_��҆J�÷w)��~�=y��kL,��kk)/��ح6y;�Z��m�'����Ckc�{�*U �.��%���׾�T����m�l�4���I�5�b���	������v�e��V14_[r�mH��3�RA�+iRk��y��߶$?bI|4V�Qo�Q"U���D�^�:;_�%^�6O{��?��qԞ�M�78�_�q���c7��U�ޗ�n?�i��?��@ �� ��گ��7>���r��A�����y���V���Y�����u��5��6s�a.�m���*�\l�퓽k-�f��g��_�(��7xHj5�~������˟�[K�K	>��Fs}�%�lb�?�^V|{�����'v��P>���7 ��<xTQ��&Jt������K�����]��p3��]���{s=@2�۸l��;�����}�g��������o�O�����O~(	�`�f�]f�9ކǇ{���/�Y{߯EQ�Ɵ0�w�{�7�>��6�UF�y�T��[g�V+
���<��vw��c��O>�}H�x7�P`����Xn�cJ��Z�.gK�L%0l3���k����ɏa��5(�ڌi{�2F����vT���� UW�z1�?<�h��W{�<�/�J����fa+x|7܅�ُ�wao3������:�ޗ�[x�f������ѯ�����7����ix���������)<w�p.�xy^�c6���ҫ���)��Y�๪���)k,�Y[�,�rk>���UPO�c1�2#��>^�b����Ny,�ߌ��h)0� X>��Ǿ�6��Pg�O�k�[��m�*@��>7�Yb�[�^����K>�}~�)���i���Z9p��6^/�Ϩ����Q���u&���E�h,�є����n�f�kL��T��a�c��<�ˬ��w�;=q5���53�c��f�w��l�F��%t��>�z����O�ZS�P�l�Y+����鶆K�PP�q�OҐ��Q���xJ4L%�i�����������v� ~������^��l��1ߥe�6z
���9Vk�q�� {�Nmn�vޥ�ϏƂ���]v/~u�t�Ml,��=��Z���ї|���VR�Ă��\��\�l��хc��Ɠ��n���|�ȭ�U-`�B,��%�[i�﩮A����G��D�ۤd���
</q	�M��z��/?��%�J��<���m��T��y���>���Rg���^Rz��Z�$��u�N���vj�mh���S�=Y��௲V9��P˧y[D��?=���	�z~��Q:�z�1���
*�����ŕ'ʔĺ�b�{��@��mI�����}׀xS��]ZOÒZ˥��y.-�j�d�s�ז��O���x\,��]bsM�hOD��4||��xѸm_�]���}Β��}�]C������TZ�Y2�$ ��S��5�M��s)�c	G�oR��N�M���cji^&rl�Ǹ&$��%�����xV���y9F��[�)����c���:M�
G�������B��,~�l�k伜��r���7�VI���uL�����m�uZ�#�jۨ�P��,ߢt���]���<���u.�է��o��������  ���  �X���+�hb�0����_�0R�R��.�>�)������e�Es(-�;͎[g�����zJ�Y�j���՘?d�q�}W�W-7�2;Z�ͨ�MPt�*�e���UD���O�G���ҫ���iR�o�����\3�w����V�.y�Hl6�-n�m	:L�꺛Ȏ��L�Ċ���X�}/-��ژ����l{*��_KI��s����9nJ�mmӛ�� �>akо�j�oZQ(9�W�U,y�pլ�ן���ÿ�?�u��[߼�n�S�ۇ$��?��������t>�R��tQ�|��y�w�`KJ�׼O�ϲ�KM*�(h>_b�w{�ӳ=�׾����>�<H�DK_Z�h2����lKط���I5����n(AQ� X֤�E��͠�F�s��<ϓ�=�7�g��=�a����
�;�ww�7�>��O��P[ה��|l��ł4
�(wd�ҋ�8�B�ǅ�M�y9|?<��+��Z��1ܥ;��_�;���?�u?�<z;,U��>��1.���]Ƕ������.�-����u� ��NX��ű*�A���T�"D�D	(�Uog�?�=��G.������� �RZ@Y`1yЮ�5�㆒Ь�_J�YǨ�����i��r敀�^FUV�j��ݥ,����	��on�ާ�P:�XՄaˋ>O��4��lz%���cc�,u����7���hU-�Yݻ�ngc�X�'���*@�5O�X�Lq�Ly,w6���]�60������G��j����?�E�O��Z#N�gmۏ���뱎�U��׍~DI��M⢠���5̘�O�Nc���c���Yq�qη��m��͏�Dv?�.@��T0]��n^�JZY+,%��4�ڦ�R6J�,�T`��詜���6�U�O���ע'J�U!�j5� q>������\�`���Է���e\�ѷ�|�<aЄk@7\��ba9G_�$Y`��{�e� ������"U14�+0�,ث�QjJ"'��ק���PI�̍%m�m�|�|c�K�[���g��Ş��]o��^Gɷ�z���}b*��z]��WҤov��v	EK@��:�A���kE����n�JG��9���)47K5Ѡ�ZJ+U�d�%y�Z��*j�X�}�\���T��ߜ��_�XP�2�5oZ*xJ�̖�P.i����Kb^�}���N[%���W;��ު�I�Z�1�=�v!�O�n*�:�����[�d^�����46-i�{�*h�����wk����æ��ξKbAc�)�:%bK���r��F�!�Bk��R���#;����6�q�'���@�Y:{{1ێ���X�3������XZmٝ�Mȸ�k����'��D�^OU�֕k~)�Υ>��D���>���9(E��ɪ�����be���kK����\�[~o�m]�8��r��X�c^�|��| c����|�9�{�f@�  ��! ���o��q
9���a�?ۄ������=�cL�b��
:��K7������9��6���< <��p�8fmc�ٸ�tw�G��;�8�l��)`;X���$S.
L��2�"�S:y/#Lxpb�c�Im��D��?[+s�t����h�tg��m�~�V���?|w%��3��S�͈��t]�n�Ʌ��(Q띶�xl- �A��#<����?�*cm?Ηu�k ���\�c�J�\�cꇰӂ������v���.�w��){�ƺ/��i��[�`��-ֿ��Y�U��b"���������}o����yY� bxQUӗ��`����6��i5׶�;k6��>��`��*Y"������xجx% �{&=�}?\�$U@B�3�H�ci6�f
�Ƌ�(�|l���cj�*@9�l��&x2H�XR&��2������Tfs��Ms8<�m�R���{.�ۮU;����Ƈ���W6[V_�1|>-h���6�?.�r:Z%�+[Ge�kE�U^!�<��k������;�U���^z���)�c^����K_����sx�Ƀ�������M�}�9���mV�����h<X;@��][ry���c}fs��\�n�&�J�O�xՁ�����7��X���QECj�ć��zM*��R��|%�����JFy��T�,�1̵:Dۢ�b�NT�F����וi.ufuo�)kv�CV+!%U,�iI���
^�wmFr�ݞJ��s�\�'O���m�g�Y��x�/�<�lqKpv�ֺ�-�<��S��!�?��><<�-��:�s]�:��no�ݵ0���C���[1Y@3z�F�X�� ��-m,m��Y��՟���H�c6��MLe�|Ix�`�N ��"��+�Q�O���*{nj��� �*�{�8�K���vĔJ��hLc��e,-��T�tyRӪ&�Ʈ�F���g�[��n�M�aM�(�j[bɌ�g��3�����%�`˨�^!�I���-�)�s��n,��[�˵B�΄���$�7��U�u^U4/a�&�{�W�v�����qY��}��?��@yy~��)g�f%/�ڻ̞��XTbbL�b'z�'
������Qw�R͢g�l�k��fIk�(;}��rQ��tl��J�oӋǵ�E�ǂ�.��@jו�������~��I�'OnDO�z���D�Wo)�ە����U#��^��x�T�x��$��W$,u��X��4���_C��ٻ���MI����v^�=��=C�ץ���_b�{����wmo	K�)A���d\�?��Қ<jV�s{���I��*-��	��(��$�~
���&_GdZ��s���{'=N]��`]�e5�ٶ�o�z(�����b�e�٘����?6��M�/z,��KݎS�FPi�i�!�>|�{��Vm5�D�۪ƜN������p.U/%y]&��s{_�*����{���ǝ�hɣ)�C~��|��������4�ߧ ��	 ����|���6����~+�ǿ�?��~7|�p8|�|��b�ԛf}�UpU-����� ��y8��C�kð�[��t>Z���)��t/
�t��f�Z3�w6s]���|��Y�~(A{���&��{�n����D�:��]bR��i���JUi*+|��`)3
h��4����v��w~�苐*`n���,d������p��}!Y[� �Lv��þ�Ô�LA�y���Zt��'Y+��Tb��86K3yۘ����6.��6�t
�^})���Z���Vтb
�������bH�s�*U������E������,����I��>XrA�q��W}��X��d�G���kZ;���fh[�(��O�����Y�x2A3��c��:٨z�xx��<Σ����@j���v����@\��9� ��x	��o%���ڪ��5S]����%�߻��)m���4�^��������>�:�}���SY�x�$Jw��<��x��}��7���+)�vV�(�uK	\ٶuC~���V˖�!���a�{�i֒f��T[�����_���u?����p����O?	o�>�~��U�����~�������.���������]���X��{ȏ��~�v����ב�F��<�-�d�d�lU�d�XL��f������ҹR;-��
(k���2C��u;_ ն;
|έ�����|�<Y(����%0X&�nWa�#�"���И_l!��^M��%<4N�jR��Oޝm�mg7����k]�7�/>���=�'�<�������Z���$K���pjK��܀�mQ�.PnI�|n�y�6cc�1�'�V��D�rJ�(����S��tT��.���Y�B�)_oS�i݈��C�Z+��0�e��"�̚���O%)�
;��H���u�pcZ����K% ������{ւf��j�f�5!�T�԰2�r2�J�����>�\�[Bi�c��J�D��k�y��n�ԯ��*�&@�<v�|����� ԄF��{�lTU5�ѓ�Z��o|��1����V������sm1&{�'���J⦬bkIL�{��x�5���<�2*x?��K}K�Z�y�e�X�����xRtn�R5w]�=��Vҫ޻4>,��ʅ��s7۽�Z��{u��Pf������1lk��}��}̶��<;Zz��O,돴�Ƅ�{E.o:j �NÚ�J��-!Y�;��ol?,����&��ZkIO���+Knѯ�O�˽B���}��CR�_O����V-��J��I�e�T}۔J�h�1
�/�V�R�u~�Sң�}�z��^��RD���޳�-�S�MY�\�ٕ�B��V�M8��i�̓���%��z/�M�XK�.�ֆ+��Y�����T������k��Gu�����~�֔j�u}�z��܃˹�������s��A�OY�q�i�UQ���6�^)6�5WZk��$΍%t��G�rS����+��8�	��ڸl|�+���U�.�nh�
��˲���^N�<�ζ�~����W�˱�_�����^  ��  �������4�7ڴ|�?�B;�>���O_N�/���w���^�������1��R@��l�n��y�������A��e�(�4S�,��Y��ق�5ȣ�t��߾�B��JZ�Z3M'�e�$A�x��4o�l��(j��g�+^�Y������O��?�[AE�v��N瓵�Pбך�'�[�̣P�s���m}���hQQ��AW	��1g���x�L,�<<є٪AmiE�6,d����H[f�6%�l�e�y���|6�}Я��}aN��O���p�����P�f��\J,[�IA�Um�e�Y�.���]l&��,�c�`N��o{���&OK��d�������^�li=�ekl,��<�z��Y-X��9��􍍟�����Re�<*	p
ǧS8��8�p����>����q�ذv5�����C[*�)���k��Q+m�6�V������z�[P3x P��.6_�o��j��}� u�Y������SJ�,���������Y}� �Z�\,P�\IA͆��K �\z6��Ǟ��jK���?X2a�c@k�gk%�� �Ͷ�巇]x��U~̟�����cq9��+������<v^�:�����P?>_��d�ϡI�y�6��I%�x���h�u-�~�i������K>NW����q�Y޺.�}��L�����{����^���fi<��B������Sf;[�TgP{r�V6<oS�x�J�u4[��)�:��3���|��w���c��)*���J���aۇd�������O��Zef�D�����eA��(_�^��{��hAE[�<���\���Ǭ��MS|���mQ�԰��rB�9}�[����:-
�E���X��`,ke� ��|-y�y�-�X`(3�Ci+��We��RI"���B?��Kg	-��T*#b�ׅ�z�VV� p�Κ�*'ᵿ�����ƶE�WI:F�$\�"�{�*�TN��j&%�U���R�R�2!��E[I,��v�����{����UkU�i��KI�ߗ��3߃��uW��Zo���ϙU;��&����K��VTYh>�����K�8x��g*Au%�uO�X����S�җ��k�
��T����8��������KZC�h�{[���I)�3����8�[�8[P^�/TɥDX����Ӿ��R�-sIV��"���v+�ϵ�Si�7���"�s�Uu\|+K?%�t,J�'{����Zf�����Ū)��Ti�mik%S��k��Vmd�w��-���G[�) ��-���o�}I:ƚ�)�&���J�œX�BJ�����KI6E��N���m���4֦��u��ʏ{k-�B9~�/�
Q�Ŭ��t]�,����oׇ�&v7��yrw*��/� ���Ug��hk��9�%I_���sv>�ڡY+����k�v6y���VX�O(��ʘ����Z��x
��cص;{��'U9��>&��w�nb�K�����x���+�	� o��k��ۿ�7>��a��7�KE �ώ ��BM~�Ow右�����������+�g6M�{>�%�����6{��?��I6�?0�z�փ�ۅ�}�UCx|�h��g[0s�JP��,yU�Z@Y�I�ϋ�lW�U������p�͖��V}��������֏���XJ�ݮ��D(3�,��<P5�6K���J�
�;'_ 5�}��5CP�(����D��t�Y�fV��Xl� ����m,@�������}X�ʖ|�SX4��~W3�/%`�d�UFx������L��Lxk�u��??т�ɂ01�,�ɒ�R�{�����<��im&��7��bl�`a?���.�S8�R�>��~��6!�l�T`S(���Ɗ��z�K�����6��d�x�,hc�*ɦ��z^kc��W�Q��[���$*�o't��.Y��n�ąi�<>��^�u6j[��'٢͌�*C�[�C��7�"�2��JU�X�{HN���Z����~���a��{B��ڼuL����S�I��Y��x��۬h��cz��H��l	��t���?��O>��{%�vvm��ǫ�}�җ4��U��������,�g��q�?=���Ƕf����Cx��:��t<�O?�$|�����ҵbcQk���`�:3=,%�X�^-�,ll3�}���v\�`�o(�a�mJ��f�v�������&M�Q_"����Z=Uf�+0�`����|~,@��+myt޻��K]Pث&B�v)�	�!Q��R[}�`� '5A!��1�؂�u��<�z�}�X۷y�K�L63��Z��Y��W�w�����~�KPvj�����'k�T���,�����䋐��K���~�n�\��43\��y� ���U,�0��NK��5R�Q�3�SIF/��wiQ��^U`�����Ak�X�h-��T�Wk�,��^a2��ڵև�^v��z�J֪J�C��e�mW��-��U���ЖD��}��u>���4��[B^/{�3����d��>_kj�{���Y��|�ԫ��Q�V%,��?���Fm�RU�	�I������[[�E�$�-I*�Gx�c�/�R��|]
_��W{��h݄]>^�Ҫdom/S���k�A�{�Z[��#K�y��=_�zJ~����K��K�L�n��\(��I�jkAMb����{�e����� ��E���]��|�우uE,a-�b��km��|.���g��阴>1AI���EӖ�'�oQ�TMʺM\׭�Tp�D��%�e�J��|,��+��z:i�{@L~��*j��S�A�$K0��?}��22�����S=[����mnXǂ&XM����	վ\/�$��Me��ZEVO�U 5��VYE��TZq��,����8i}���ZSM�j�0�g"�'�<��׬��i�qѽL�/��Ӛr��e���x��,y�w�u��c)����*��0��_�*���t8z+�������]/k>6����d�N�/��/�xWŧ���{�������X�K�^�����_M���y7��G������������η����7�A  &$@  �w����~1��(�����W��������i���ώ�n�Yl6�_A!�á���saX��*�3�^���+���&g-�;M��|0��ka��@����2tWp�nw��%Og[,X���fp�>�q)˛7���e-b���BD�����[�k��0�jUc�%02/���],3��k�����-/mW�~k���Q�f�}V��-1�:%w{[�ܒ����{��RR+#��ǈeF�E��g����1��rkM����Ѫ���l��୤�Q��n��Ǳꗥ�:O֦�f(ۂľ��������o����Y�]��ݰV��T�|��΋����y�P�S[c�TЄ�l�:S�����x��{舘�Q�Xe����I�~N�7���l��:㌋�5S[s`O�O�PR�_��i�sk?u
�|L�ǳ���8��X�e����C>fJ6]��&�[K%k5�����O>�A����{�sc�b����l�mX�Yk��qz���Hۣ5=T�V'y��6���ޕ���s+�Œo[��8Zk�k�*L<(nɕ|�*�����>?��T+���8)���u�m�΂�%�|�_)1�����6{�ß�G���A	����}U���Q۬�}�{�㏿o��>}�I������|�PI-Y����}>���d<��'o��iW��� iU[���~�ۓy �i� �`���ֶnS@���Z�t��/ĵmO	��hA.%,�O��ӕ6g
���{�5zJ`΃�]��~�8�1��Vۣ{��#2x�,�^�h���r�Y�}�
p*Y�D�����<,Ȝb\�+���B����*Ѽ��~�}o�q:��<���{��ɯ�.vv��5f��k�SA_�M%?l��| ��|m%]F��j�k��Ǔ]�V����}Zm��z�X@��6>�ڢ��w�wv_<��.V��%`K>��:��%���e�*�t�j��:�5���_/mi4�,zk[��V���mM���� ��ߗ�RJ*���E���e��|=��~��ci�8��@��vd�t��l<N��i���q�cvz��j�,��uQrv.����/�l	w�k��m��Z҂�]\��%�k����{�Ȝ�ZX�/j�y�[�KP�5g���S>G�y��y>x�����JsY��_�t_�z(��}��Q����zɆ�l�`��㬵��6X���v{{M-��4V�5B�ܔ�Ӷi'l���kX�-=ako�^�0Z��갳�J
b+Q�_��۶][a��>���i�����+�lM�&������$�r�6����KY]��3j{�����ۊM���P|�K]X�&�U���CY ���\�:Q�g�V���OY;&�G]�C��~��~�_OlM�N��j⦱����~mrC� c����>��q�z�H,�@z�]������rmz�S+c-A1y���\��t��kc����x,��.bn��r��7��F[;�����;ںk��(������1_���/z%�����l���k~i�μM������.�����tY'xL�Kx=��J�M���3��c���|��w����k>���k1����q�ϗ�~j���~�ہ$ �ς `Ӵ�Gj����*?�G�o���9��{�Uf�m����fG��;KjجG���2Ki�K��:�����j��Pz/���C��Ҵ�AF���?�4��Z���2�9�s	��äv�V/���ꊥ;:[݃s�fF��C�35�2�V6MS�#�e�r��m����o|?���/��z�e&�Ս���U���^�����$4q�F�w��5��n����,��|�½��:hчx�v�٭���ݗY�
�u�fFf�����c�y��y�|�Q�_FO,���R�S�hZ�x�u��2;=��ԪAj��n=w��������B���z�ǩ��,�N�r� �O��ė�P���f�*�Q����B��*I�K���D�ك�
>+�1-�m�l�iX�A*UB>�tY���'9��q%�����x�͎f�~v���'�m�d�'�^�!P��V˫aX��P_�dǠVZM���5��ѹ{c���r�q����?��&�|kaY���-�lFjc��fk�����C۠�-ܾ�3_�D���[G�͛O����Mxzz>���tx���lɠ���z��qN�4m��dɘ�ۇ�6O?�]��ߕ�W~OQӪ��E�W�h�|U!�X�4X�S��@�ֹ�qT����~��E���9�i�U�U=�x�d�W���꿦�VCY{�i.-tj%����٘���Ft	��~�-��z3��̖�ʝ�Do�^y��ci��=G�����s�?ۯ]l=_�fo+I��*�������틙�VM��m�z"ξΑ�JjX��Ҭ3�U�u/By�H�x�e�ǒP���}&��n���q������d�Ӻ_k��_���}@��d�U����e���Zɓ|���k��+Y��[[$\�}�k(5֊O-��?Vok�t664�'K�����/�lm��dGWZ���y���j��=�Y�u1g;F�\�NA�R�-m�< <�S��k{�V�uR��nʏ����nh]T:����Awk�9:���$��z �vt�W��������~��;�6C� ����
ڥ��+����.���d��%�����t�/)]n� ~��-�l{�kRO-���=!��*��am�(|�^��^�k�*�z�[.��0����}���[iZ^SiK9�uNT�T�C{.��赼��e|<xk��]�:�1\׍��K�����F�V���^�Ke��c̒��\��SI��}��58��X��ܗ���^�-K���Q�Z0�%�]k�/���9����G-iio��=m���SF_�ê�u��B��\ˍ_�e;���з�[�\��Z��j-{�D�WOe���x*Un~���`%::�'���%��qWb�_��w�u�����=վ��ѵ9ؚ2ݝn��޿�_z���_��{>��ꏩw���#I ��	 �f�����o��b9�˷�����I������+m߿?��εE��{�m�ed4%�V?[�}�}�k�؂ %��5ޫ������V���8ciuӔ ��YQ{����mg��J�K:k������A3����'ZkWU���>��Ͻ-}�k{DN�w[���_�l�Ǩ-�x�\5�-��L�����l�W�O��ﮭ.jPӒR�%�y[닮?��
�d�����h�"�o��.K|Z�NӬI�XΣ�S���٥j��%?Z;C�v%)��@�f0�V�_����
�:�[3�-������U��������1Y ێ����+�GT!P��Foy�L�x�-����������`��i��C��=
Ћ*Lj���%@��u��G���bm����h�$0�M��&d��PeB��W�,%@�݋-0��Z�I�J��mSI���vj�֏i���@^l�-���\��Ok��m=���?�<��ܕE��@��gU���+}Խ�������}ث%��*���.����n����׿���?}���������|��F��s��9<?=Y����݃��xz���5�&QSֳ���uNv��Zҩ�N,��[ox�p�m�C;t޾F��چ.��k�\v��>(M	�����:Ҹ������_��¯7I�P|�ʬb-�l�����N�G�������x{���,^�V���lҹ<)�Jk���')H��ٓ�~�K�NE��q�.D�k�6��v��v����Үg �Mע�^��USY'�ZE_��*�t'���ۼ��;+d6Ƶ�t�j���{e��]�a]#Bm}�^*�Ub�g�X�,�\ۄ��	bOlL�M`i!���'���kkEo���[Y�y���}=	-"?�����7Z�`��5��%��:���u�y~��X#j7i����Z��X:^s�XX�n��qk�TΑ���A�j[�|nK۬�T(\��V�UZ�K�/m���C�2K[Hc�5f~{}�˚Ve݊��n���F,	��(���%���$���vg�����N���2K�eMF��j,�ea���U���n,�ec�|}]&-����_o홺���/q����u�d�η�{�����X����kM4e=��em�V+$�H�{��]YB����ɓ�6�!��_R�]��c��\IԊ_��.��6�q�\�ju��;ձͪ^J�:�e1ZrZə��Ur<��V����5k���fI@^��1��]F���{��Y�U��V?��8u��q�J�&'��0��`���uc������{{]S��bk�56�}{������۟-�����z|5��KmO���H���]3%��b����|]�������U׾ZϽɯa�|�����/����h��<�*�;�۳,}���U�OK�?=���àY��a�j��M"	 ��" ج&�v}�W/������Q8�_����?���S�}v]
0��E�3�kr$�E_k��v����>���u�viY"����5sO��ۦ|�/��-ȟ��t*\��;�V_�ӧҪb)�5�0�m+�1����n(�ǧu�i�P��%	b��5s{i��#�@��~��bIy���A�>0_������'�q��قУ�8���D���f���������X�������3&�I�5[d���QoK�,/���X����*�q=F����|�q��1Yu������
"���5�R�j%K=f�&�4�������+�L�-
� ����7����x����p��VM9���ŪmQ�R5T�:�
�+�Q��!\���9\�Z똮�&�n�L���}��̶�ߗ��x�^��=����� Y_�I���ϧ�K���<�'F|�Ԓ붒Żި2)Xp�<=���8�ó�hm�;BƲ��1���Z��\M8/��i�y���.w�i�c���܇�>��yoK��o�Qil��~��C��?��-������>}
ϧg��~:�c��Rdm}�%��N��ӷvB�x%[�\��k�2��8�-�Ex}���Էʠ�*�|�x�"���i��l��&���5ө��X�
�R%�����)�2�;���(��|�kJ'�����ڦ��5p-�g��B�����Z˝�?�P�]N�5Ц���Y-���Z��&�,8����ݯ���T���d�JдeL�{J2j��x���zmsM0XB.�7�7/�%Yb�TE���eL[����S]�!*wW��ɒ���z���k�`� ��;o�����/Z�ZI���0���q��5L��ji�ay���*�R�g���,o���Y[V�*�d$�����$S�:S�<^t�4{\�4֢NCMn''�߯��:Nۥ���Fk����$�[�"�}���n�q���~�|_���ak�D��1�0���|�y�j�N���MUI�^��N����IY���7	�k��'<�����忕 �D+���p�E���ֱ�*U�(��Z[�HU<�gvem��*`|�p��[�>z�K�l�u��f�Y�y�i����J�!�3k��<��%��$Ȭ�`�IK�,e�h����dS\�6ubʬd՘��/�����mK��c:]�U�$�֪�˹�1��`�E�K���#��n�V��5�j��h���}��ٺnʚ`���5�l����]Ǚ��u}kҰ����<v}NeG,�z��:��&��!�7Վ/�$g��&�l]�'�}m�T.���5a}�V�,��_��?�*-���p����^�������|^��4�Ov���GKpM]I�M�|����-�����Mu�|��<���}���RF)���W�[�?�_�� ��e�͟�I�#��ȫ���;g3�� ���Y�L4�h2�i�L&��2�$�l�$W"����]W�
��^DT}��G��uבGddd��s����h+����mmk��l�O~P������m�|�<N��������RMboļ�K��
��C��2\�g%D],k����T|��x�_4x�s���U�&?��BˍD���\m?D��X�Ȋ�Z**��Jn�S����'^�p�)�k���TLr�xf�C9�2�AU®������j�z[ű�]��y���ڝU��܆�����{`?�$��k��TX
92{�M�������:�Ȏ��>
�c�߰���/ 	,�
��h��I����*�X:@=��H�P�-��3AB��?�c=CO	���5���N�vL����z6�[�G�����W��[XE=~�� ?왆鬄AV\���I�ns���d�i�4A� A��N[wj�58-N2��Wo�5R��7�������@k��(]ĦcL�0/�ɬ�n8��@��)�-D��8yw<�Z�=Si�f�Ҏ`,A�i� �x�fT���6t�Y���><������

��o={F0���G�Z����pp_����ꗟ(�u8�݋x�^�~�B�ǳ؏U���+'!�TQT�	 �KP�O�@*�?Sux	�Χ��	j?7/FHi v+
��K�9�t���N�tÜHڶ��*C��1�)1������s�02		��W[�Bj��2w ���!h8��� >��VevFBϪ����p���>�
e��Ԙ�Q0쿅sa� JuVq�_ %�@Rň>#�Z��U���wfw��҈_����h�d���ҟVaO�B��03CdJ qSIΒ������8:����I�;(e�J�0��,�,k(��VPLwY�H��3j�(Hj��Մ�&{.ZOM\&TS0����V�?�@2�r(�(5"�s*+�T ��u��l�^�L4:�*�r���([�{�o�v��/n�,K2g&��q}���L��@|������T�
���E]a�`�Y���1�c!$;��z�U�x�햏�VO�$�UTa8�C��򾓱��4��҆����a~�/��y��'Yg>���F91�
���62�qM�fUN�y���L�gq?f�(I��kN�O�K��µ��f̕YԚP�V��Lc�I��_��d�\�d����`oy��l,6��:�h�I`/��ۈ�ՙ�'$=/f%qe��%�M51Ϟ֋�s��{���2x?��Gd�	�1��n~%d"�s<��7��p��H6y~�����IZ{U4-F��2gLB���y��=UG8t��@�8e�(l��mpO�<qO���@Ҵ��v{۰=��'^�@�o`�W�(,
_���k��y���n���y\��Ϗ���}��������[��ֶ������Vdmk[����{�>��4�y{����oW���0����α2���;�ʷ*�0�B5�CUb%�-��B���'��T�O9t��@W�t��K����Im�<��ڏ��  i�K���fd��_+Abv�jA���`��.=�+������	Sc$0��Q����E|������ ��k� ����`�����9��:����w=Id:p�P]���]Ǿ�{��X- @��J����l�cǧ"H�*j�Y|�GUk�r��Y�'؅�+��L� u�Y%��@˴�z@��ާ]�0q�k� X���_�Y)�w%G�)�������T&H�5-� ���)H�X�;���D4?cĂ�~�LPEUb$��-�S��6C�h8ff)u�6)m�jͱ��c[h��t8f�&����~����W�� �i�	�}}�RɕÞ�'��l�����4�����@h��o� ��f�����p�>���Y�)4f�ܿ�8|�����%sF^0k�;��9�8�i"�l�fQ ܘ��� �FZPq1�[r_ �ّ�M�y�P�YIP�;�>T�R�; }��× �n���oƘW�If	�h���e�� v.�c��@���W��*l���'�fs2�����0�9����p� �/̣��epq����ʕ�R�C	E�r�����dU�e��3+���.s2ZS����Pr�@p���hFI�?ޟRGV^�j*�@pc:��ZQ1BƋ�m<Nb����Dd׬�{G���g3�ASw%�d0A5����%ƺ�$t�H���	JP�,�!|��>E,4]�<���Eh�s�4���j�4q���:�N�1.6���Nj��@�V��)���"dn����t�����y��H��4X��J%~��8��Zjdߥ�a"�y^%)��xF��"�rI�O��Y-��|�N�2����i$�ַ�L�,_*�0�4g����n<<wLiC��:Y���/��^C���)�;� Y7"TLD�<N��g��y��7b"��)-_0j*R^��\�P��/-� �'ف���9��s�����dL���K��$:x?$�����v�>���pN2Q�-�~j���%_��RL��U��E#i8�{=ڈ�b�&v�bi��/�(��=\�G_��A�����!�LV#�>?�d2�F�KA��}��0ɜ)��r���ۚ�d�a^Ø�=�,�����Vm��y��r��>��s�2�����P%�6 �����w��h歶��~Ӆ8��8�����H�� k[��ֶ�k[	���mmk[��]k���i<����G��ߏ���~��k��X9>&p��i;�1�O2&Qq���E������,ᜮ+%Qf����>x��f3 �1��S�@R%��"^̋dK��-� ���h���;�bI��B%dK���!fm�H��TtE�� *sk�SH5�o�,�9�o豏\� ��8�;�oG�� X��&۴��+L���m�m�x�:��X��� <�C�^���	`Q�'~�ժ5��9�RI	K-��������dl���y�ϡ� ͓���T�?��� Z�-�ɟ���,��P��k��^�TszVv���3�X0u` ��b����jk�Za0�C"PLYa��F�VVB:����7�3?������Ո�A��)9pBP�^����m,U�B�4��HՆO� �sc}�ՐV��5TJK�T�ۘP��M�a�`��x���Y��ڟ�������bQ9ȿ� �]|��k!5���)��8����y�
p��� V߸��g<�x���z�4��� ���x8�ׯ�����;���)r�?��9����z �,�^(@��5�$���lObT�s������6�� ъF胂��X�5Y�[���9H�Ūfv9A���{���<v��
�R�2a��ìs� ��Y�I�3��ɡ�  �*��BWMȹ; �F"ӓ�r�}4i�C���M��&V.����w2nq�O����u�oP��y>��0�5��s���9�1�}Ns�&` ��t����9p��b

�n�N-��0�B�Y,�p=��j'Y�Di�(%�z����d>%O�qn�P�՚��B��J��9��#�Pɵ�^Z��:�Hp����R�������
uaE�r�y-[���r�ɝ�)�o�.�s� �� Tߔ� ��k��!y7BT`? 0;/ny\��$  �����pLy�Q��P��Y:�%�XI����W���*#*
�#���$������=#rF*ב�A��`8�~�:n��0���cۺ�:���"DA��C���?H�I��Q�]l��^(!���u�����4�Fĩ$�~B �m����l;�,6�\{�r�K��c��ߧA�CF��q�ϝ�����\�E�_x�Ly<Ἢ���c*�tb���4r��}U�HVG� �	��I~8]��q��s�!�jƽZ�_�5�:���d�j��?T��A�9�=I�L����=��K�C1��|�P�)
�8�"ؼ��-�����}8�݋�����'��x�=z�c������������/�װ��~A�DAT/����v����m�3=����<���������7�nmk[��ֶ�����ֶ��������ǟ}��ov]��e�������\���XY|� �ZU�)�2��
R�!���%U%���Rg��@��n�]��Ϣ˲�dV��S�F�j��5l�0mG T���������nv7�C�b��u������b �Uϖ!����1.kO� !���}7��j!` �>��!^�a�7S"<L�aU�Xƈ���V46�T�Ǉ����d�gu#D�SP�J���F,�H|�A!�ͩ�E�G� ;��Q��
g�x�C�#�%�*<�Z៭(*���!ʥ�}n���sH���`��N�BǇ�L�N�^RH�T�י�Z�d[e�Q��}�6}έ�ߴ�Qe �K8 ��o\��uT7����%3cP��e���#�^�#ԛ�r�j�IA�V�odʠ�0��|�vc�*�@��a_@�}(]��a�.U!�F�9� �=`���+��+r�؞�o��x����	��E�)L�I,� �WanŤ��� �{��� �h�7�2�8!��b�m���w�{��}�9�ss` .����/�'��[���g?g���?�q����i(@��-�w�*����n�@�c�fƸ���I�IT�C��Ǫ#!�q��?������~�U�MMo���~ ��̳n��x8T��VL��ݪ�bUd����Z���`���M�b����*Hy�3�?�T� T�H�>�\���<6H�.xV#?s�8:��H��\����m�V�D[:|? ;y��jfz�,� ������ ����� � ;���}SI&�4�����I�4$��\w�VJu-�T9�9�Y2 �O��A����B�`�Kg�+��X��AZ�F^2�f�p���aܟ�������#�PZՒU��Ǔ;�:�8�����Q w��7�L8�B��031"��:����qc����K�N�b �d�8W�����僑,r�u��7Ǆ(j��e�r��,��K2��)*��8��v��Y̅>΋�2���**HĦD>�}�!^�G�$�^99nΣQU_L���H@�fUXm�B��dI�ډu�|E^Юk�Tì}��3��T��wL	�V����Kץ�qCRʽT�H�	I�T�4r/g�&X��(��It�*��q�K*U�L�X��8'��K�e?�z��d���.ܗt�Tİ����I�b�ѷ*lѱ����}�:��U���%Np��,J����F^�7��+��M��z��}�▖�H���sQh�������9���s���}����dc��l\7�����]߇�<���6��p����݆8��~����tk[��ֶ����� k[��ֶ�ߛ�����e<�7,���<�Q�����Ӷ�6�������D� U��V�I@�@�n��ϔ�!�8���f��N�#����-�P��:y�3�'�Ou
0uZ��GQ*O�������d���RA�Ǐ��ֵ �Ԗ�E�g�O�N��ٱ.�U�r�C'� INmH���צRk������'K#�gG�1K�o; Ė��R��ת
�h�D肯�JM������&.W�S�ڶ�!����F���K�U�A*X�mz%FX	)�(� Xb����w�g<��V")�d\�i��X�a�qx���ܓ�[Z��
��̘H#$�"*��~8N;T���T@\���~&�d�H�v[	�?{ 
X	�!�J� r�A2��T%�Ѩ�Ȉ��I 1 ؞aF�t��V�����ϸ|#%̊
$��X�� 9B��fGP�,���Q��*��-�%�Y�������M�hꞺ^�JeK�G���,��V��w�x��>�K�3�e��� of,r U���q~跍�$���	��v�� �p� Ԡ���όg�f�r����<ۛU$��B�;lp��ҐQH�9�Tڅ�| �²��Ӷ�܀}i���8�8�؇�����%���ÃX���|��+����W_��ǟ�/f!�dH�Y-}��#x�K���@�J�M�Ψs��c8wN��|���މE@A � ̰?+�P�,���'�DM��UA&d&�u��!��^��x��VN���xñAL��������G{��S���n\�(;�9��Z����@t���Ǖ�S��ϩ΂��v0q.�N���9����>����UL@�(����n�q5ֹq���> ���K�=ƹ�f<�����}�N��� ��߭fJXh:	l�f1[&yM�b���dX�r�k	&{.�D�&�t����H�W���J�壘
.|O��d�Z�N2�e��H .��h��)by���<ݮS ڱXa��Jd	i��g*qd�ȉU�I2K�C��em ���
�1��x(_�m���2��.]ho��]C�2 ����H��{$DX\l[�66���(����%���kfs�����[�wމ������"y�{��✀�$	ݡ�~q������>��:Ι����K���k;˜�g�$A ����<5(Qa��P�`�bM���,��=��>^k0�*�1���x~6�!�3�+��ms0~Av$۸��~��xu]����T����M��q�LBt���؃a�z�u��d�	!2u;���Ǭ�����zR�}�z[��щz�	���p�,>�|�
�9�<N��vlRo��o�M�N1(��U]P%
I*����'R��L���*���V�Ÿ��8�޻�������������/����O?��=������}��W�Vi�>ާ�݆�Y��Y$�3u;������w�����o���mkt�J��mmk[��~c[	���mmk[��EC�G�7��}�>	.�Q��7�C荫����H�6��l3��
�  �A���hAA>#?rF����]`0�a�K���߇��	R7b�d%R]^�~� v�T?9�C+A�TլPgu���AU��"dN�p  '�љ`��90`V�����G���O�e�b��/@�����!)A,l`S�@��.��g��SO�þ�d����x���� ��7+�������b3.�T�\Ț��@&�)ed�wS�BLU Va�ZAUI�`�s�`�j�% ���S�lxL�P*:,�bV@��%?!}��e�V�V�y�G���0u�Q-��@���S����f�D���1�= +p���7���t;K�,�ײAll����T�2��Ϧ:��w!m7�wws疆��i_pΠ�0��gJv[v�m�Z��ݖj�AI�������c��G}�L��,M�4�B2y��x�zo����ϋ����(^�$�Dȕ��?u�ݦ�1�'�a�| �G����������/�W/_���$V[ ׆��#�+�h�/�A�r$k,c�NU����`g6��*�7k�;�׶�
���l�%3g�/�1���j�4�����!q�T@�Cs@?�)����|�gOӞs^���2�\wB~�`ٓ��b�8	I䤢_B�d��Pê�:�<	a��nlx��mY��%8��2�b�/��@(sP��������5B�U���:�#����BV����&>����.ҍ U�u Ǜ���*�����B�7h|f���1� ~��5�9,���d
1�;
��n#s�]'�+/�q�4L����p�>��(�ĎL��kwq�H`8�o�~ױ%�˛'O�N#�Z��`�׵�A����p+��ؼ�{O��1cߖ|�a��(�S�-ҿ2-o�J�ׅ�{����F�G����x�CG��eٹ�f��}�]���8�WڸG���|չM�a��M��s�<"8~��x��[�w�q1������BP:����?��/�/�{y��|�C��Q3�F�GZz�Nb�@��|�ʊ�~6�JҋZ��i��岤9����������q�o�Q�uV�Z�u���"'*&��2��6[���)ʗ����S웒=��)I2�;�rw<T���#W��&|�b_i�u՟rVtf�m�e�1��a%��AULPhQi�W�����*m`pJ �	��!����7ލצ{~d��E[�D8�~��s�wM�H���u�ұ���������Ǉ��?��?���mmk[��~M[	���mmk[��|�����o�+��e�߉O�?�����~�'��lS4���� lp��V��F��ZI|���Nת2$gr�\�Z���W���T���Â�a}�@��@d��\Z��ij� �[��{����7�<�	��k�N�������P��
�
���i��]�u�Z1������"@��Dp�����e�1%�2Y�P�X���>�v�6!�x�o���j�؁$�e�d���J� ��=Vڶb/A{_�!��!U��( �Y��'�4��l�HĄ�<��q0��Ϛ&�&-[b�8��a	u���{��b�|���ZU �b9S	��Ăt�H�� � �8ި����� {��И�DZ�҅�#
����s ˛
K.�c�T��C�tD���d�E�pY4�U�s\H���	*7��$��'b�Sӻ $�A	R���o|�C֙Ձ,
�td]�j#$��궃$�2�B�	*���VgfܮD�'9:)�*�����]Q���T�h4ƅǘS�E�>���x<5ns��� T��]���iI�1o	bo6]<�5<��ѹ�x�0Xf=n<I�:*��z��}��KV�ά0��!�����ix�X���&k�:7Nr.a[Y��v$q'���hpN!��h�J��ł��� �K݊� !,�pJ#����R��$ L��XB��&�n�*��U l��#�0��̡x> �G�¼H���^�2bGU��0�76i�\��OT�`<���q�o毀�bυ9�Zd�ԋ���jq�y��zn7���� �3� I�e�v\B�W+Q�A� �I�}ӫ��(���t�ER\��i��������k��JNo�HCV�9���$��6���6$�h#5����]���T�h�ZQX��zwb������Zm�?(��'�46��d��趸��Nsf��x�����D-�s�W ����"l��0N^��3�:rn�`w�.�V������>Q��񻐕�t�A@���r��wX@��ٳg��
��Y�(jh#4 �Lu��G����q{{t��g!vqݹ���,�Ah��7�?�E��É���$z��y���ի�8G�*�_���3�+o$WAN�����%�5}�
�� �M�q���`����T����w���rd[-����}�|[caB��e�e��k��H���bJ��v��S7�y%_2ɫq�G��E������$�����]�H�BAk�dP*z�wf'�(f�s�Rd*T&���<���2
�����&^>��C���
:(>�8����"��9�EeK�ڸM�n�i�Z*R�1^_�q�^�3��O�������ӿuk[��ֶ��}M[	���mmk[��tc��<}�-���H�����{�oǇ�����Va���.&�������I�)�`Z�U� ���K�TV���o���$�� ԅ��R�$���|{0�*�>���+�a!� b ���Wr��8�v����EX�-�t%CV��U0mb��x�;SoT�Rt��ՃSb�C>��U����g�Օ.���V �<1�U��>�����<lrb1"��x"0܅�;A���{V�9�6i&�i�#���y��7x��~ݓV#Nb�YF����T{p�
�����ګ2gQp��{fb�� T��H��� ���Q�d���X�J&K��
�~�b�Z���(.$��6��xf�a��U�O��Êw�Y#�n$��o� ����1���>Yv�QFd�b��VDK�4B���Z�h}"��ا��K�'�4��� @���^�(�`��N�3D�3�#������ CqL`�ST�I��b�T{�JAIC�ߧ� I�mk{w�ۺM�� ���q��ӹ���ً/܋W F^������Y"���� !��Q���vf
M#A{�!�����8-��m���jɢ�l�Bι����������'s���[$�V8�#-��벎ZIY>;�&#i��"�I@ݬ*��ր ���-	���Q {<�����ZLrd�8{����
�y�胅 �THԙ��PƵ�I8����Pm�����pp]��x}]l�q$�p��?���]]q�oo��� �
��_�5	�Y��)2�x~iw��6m�b?<�l����W<v��fXB�j;��x�J{����Ei�g��x�ww�(��2޲����/5��
IR��#
XՁ �fa�1���m��l�����d~1.s�\��\�]���InVU�듑� @8�,�Ru�]�07o�wi���Z�)��B�.��{��-�5���gs��/����Xq�i���
�x�y��#�#�;%�����~I�l�H�)4��?������_���ۿ��RrU��[�f�#�Cл���g _@���NCM5���'��l��K��r�e3���[����}׿�z��D�ʏr�]+1�u��# #�l6���ݡy/��D���~c���%$�+Hg��G���&�Jy��"؞��ΐ�s<�(p��|�ע�L�N�q.�tNE��/~A2t�Z�����9�qss�G�0���%�D��}���x��|W��=��`�o~�a�?����[��ֶ������ֶ����w��������O]�������}�L����t������՚���z�iV�[��h���To��9J4T��)��ϔ��d�)i��mb�U�r�|9�g�,���ҿ��w�ճN�M�V͢�^ �Z�hQ���A�9I�p�qY<���0���% G��<����&��.ۢo��<�I=�9�Ԟ�T�;F.��\� �G'A� P� M�*/V**�"��b[T�a�[��U����V�� Q�C�؆Ϯ.N�w ���K�)���Һ�b}
�.^-b�V 87�Y��H�~�jw����O����h�% (���*�Yl#�J�Ɨ�Nm�d��#Y��*�~ �3K�2��T+f�d�Җg*%+1#hM��0�"[P)ȉN^4|�� ���1���b���(������۶_F������������L�K��b�V���8)�rԌ
X� �.�3��#О���'QuU2**ڇ,B��z?.sH6S.׷
̞�V{�*�R�U�0O�s�����/ ����1G��:�<ݣ[w{�s���*hFz�S)w��M>���^�� ���|<��� �>�$ �o,U�z��;�m7�`�%�V�d1� {�|m/H�d�%|8����O�W��Z�i�2 "pn�j,l�,L��=#ʰL ��M��R��Ѐ`�g�� .�l��I��u
.�fOιE�K���Dr���i�0v~����yxH�9M\���F�O��n���~��1�]�~˲���6r���plT���fjƍ��{}��4�|a�E�W�J�K���{ۧ�mC�O׃�ld��%���]�P��k�8+1u���9��j���X��ꯪ�yI�}D�ǎ�C���8���R���HQV������V3���υ4�d�/�y���e����j+�K�:/T?ɥx���,�	����c�?7�
��
���=~|������s��[ �OvqO�xxp/^�ե��BTXX���$�ڬ������7gs\�$%π߇��Y�ݴ�L�\�ڕ��~�$(Ɍ���ܫ�k���,��ϖ״��li�Y��	I�軕�����<�Ɔ�؀�J�(7E�?���ҹ.��8�An�R�����|��C���6qP�f#�&Qe6���SY�L0(L���m�\���/\�ٺ'O�ۻI�\ϫ�
�#65B���q/��n�F�t��x^��UՌ����>Z~���[��ֶ����h+����mmk��l�'?��4O4}���4|�{��j�?|8���m��Oo[����� c@X8�][��R�ث]���x���l���Xj�*@�e���-k$H:�!�a%��Po.۬��!. 	��H��t�i��Q��@�� L��X�H%ߜ�{� Th��_ݻۛ���S#`|=0cw�s��Ņ
$�V�b���LV�쓽�/�%բS81Cd�r�#��'	��ֵ��^��5�AJ��K>�w%C�Ü�y�|fF ��:R�y�B)0ć��e_�z�����^�����İ��~��(�8�6�!�l�R��X.�{Y�\تI �?�� 2�|^�V�V���d��X�k����<7�]�\�2���Ӷ� �%���)�Y�w����n`�-��Q�Ňt�2; .!����>4��c ,օ*h�FX����?F���}��U(H?��Z���J���1v���l| ��w���<���1p;����O����h�c��Q��̋����O�J���?H�j���9{U���^& �ﰍ�QU���ůa��K�O�j�Yu�qkc����E���B9#��1Yv�̳q@�_ ��$��d�O��Y�a]��[=ng�#�Pi��8O��>X7�|���$��D ��E��R�&���ZQ��G�B�#���lZɲ)sj��C�#�]���9��M�씰| �%H*���;�W��r9���	�¢�3��j����i>�3|��M,"A&fe�l�rq������rc�U�3������R���� ���%��c�B !(�7�N "@�1G֓~Q_3���2!**QJ��!�? Y�J������l�,ꬠ]�c�Tb��U	�*s�4�q�sR���)�L��Z�hQ"We�{
W�49��D��'�e���I�)f���yzYH��*������I�@�c��&젏�9�m}�w���c��_��g�����ο�%UN	C��x���y�\m�;��L0|��䆼�����jaΊ�2P=Qsi}e��3[�S��R�W^���vn��J���t���r�~�RD����(��l�T�Q�P��>Eϯ�In�����qz��-��ܷ"�a��t��{δ�����mӹdj��q��{8'V��,��<C)�a�tK��㩝��>�Sl;
c^�~��?z��\*���d�TBtל7�12���$u?��!���-nI��?�������J��mmk[��R[	���mmk[��d�����Uߙ������<��ڟ���y�M��|�`����8/ᵠ��3���<(�����j]� ��O,�j�4��*m_��I�i���5��FQu��^I>�*��e/�!Xj��<*�'�@u��hVK5o�/i�:��	r
zZ5�6�t��2�����}N�|+�ѵ�ԫcOݞ�
�"���S��<Ϧ��-UjZeh�� �qH���-��c �F�更�
���K�W�	�_������%��T#Lj�����;	�����!]�(��s���O,��� bǅ�F�J�	 �
K��mJ@3]
E UR� �7�R�mT��Z��*R���2K�@w����5�&
��̬�h���  P���F>�<�����e�x�ٖ�*�/�e?�u�7Yo��@qZ��2[�Rmb ��sIh�v�*�V�2���W ��"bv2�{�$�
3Z8��R�@K ���� ��- �V�cۻY*oq��C8��O�7ڱV���^�����C�F_CY0	I��\�$�R���$T������o�J�T)�l�π<�r�8�bBƏT�S]�q�0�����b ��,�)���?�K������ �ֵ����gM��b����xQp 0�G�F�έ(2�jT+���:�f����M/vDÉ�7�����s��eR�[�؃xL+�z�ιl�G��I��i&S�X����GM��L�^��&Ύ�� ��sM�Ѥ��y̙G`��	�Bn$�������&�����ᜣzd_�Y���0�S���?5ƾ[X6��*�2 �򪾈e�`��K"��*�IΦ�*U[I��
�'��L��ad�p����1��w����G�s�/�w��
�2�C�A	�MR�pn=U�X�t��"�.���-�}]�<՟b��t�QQ �M�g�c��E��*�P����w$=��;�Ao�7�&F�Ko��v�S1�w�N�ϼ��FZH��\f��쮯A���f]�A`�%�J|}�L�:m�-ǔ(�����~#1q��(ɉ��Z�:t9��7�ZJ������T�C��*�)�Y�ڥ����%H��d@Q	R�-,!��$W=g����Q�T�d�e��Ⲛ��߃X��bRϸw��#�X�q��e@��,&ƶ�1� pj�:H1�?�R`H5&��=�˗B��9D��m���<�z��k^%��q��k�B�þ[�� �wh��Y��ֶ���m%@ֶ���mm�s�����?·������'�a�#7,ϫ����W�ū�����2	Y�� �S��M��Z	<�Au��{�����rV�
 b!�"�w����P�Dg�D�#P�r#����	��S�X�DR�NmBH��y��UCE7��gg�r���B g+��h�f��,pX�/
��IVB����� �$��P��&�ك,W�� ,lM��JI!�]�����-�H�8���9fu� �;����>&{�������U|�ڥbQ�|���= V3�3|!�Y� d� Є�E�[7w�����Pa �Y/0JHP۠I+p���a��V-�<0��Rm�0�@�s��(VK��9[��9 �K�nJ#"`5�� Ph`k"��Kd��I�4I�!ă#p8�礐���Ɏ�*l�T�>0���4F8�DE	rP+�P��� T����(�~��ŏ_�?�����((UV�k+�=X����p|3�����5� :@���{���I���Z �`Y�c8�t5�2�o��~`;�C;-�� �<$���q�fe%�Xw
���
 <wr��|�%��6�HOgQJ8z�HNھK}�8U����|<�����w�#yܚ� ��ގ/����^U�;�&V�'�j�`c��ګAYɭ"�a�<���w|�D�iL�����c�y2fFUn��p��N�H ;͈�9�RP�����s#Y�QA�ŗF�c��bN�iVe2?�U�	)�.;�.�/���A�e����"�h��p����#��T"������<	ʻ��F���N�S<�'ν��P����2D�snIDd9GL]���(����c�1#`v�z����(�74�P����8R?�O��,���QX1���'����N��wr�2��}A��D�e�8��/T:8���y�A �E�]HYH��|%�3K`=I>T��ꊽ�vU�+Q���i��<z�nw7�?����o�_���Q�b~�Ir]��^���H��uY>�]�T��r�GiM%�v�.�kH˷�y����l���] י�
�R�A)��\��Dɞ�Gb;�8����6_���59��d9L�h<��Z�&��P�@�A���1�	�A�m������ꤲ-[E�]T�8o�牪���I�;#׋ϣ��Ž%�������{!K��@�]� l�W_�p�^?���}�=z���A��{V�"���S��q�p�(:���֣�p:A���*�������������mmk��o+����mmk��j����O����������n8=k������p�7����(���pH`�6P�
�@��J�<�dU�!������hj!P�j�eQ��"9A�LP��zH]2zV���J�X��$fP��l�ǂ�������p�Ș���|v��`f��m���э�L ��=��M�q��W���Ä���7�ӷ�������������nn�IS�����a��E !�8aG,�G��R=hDH�5>�nPi���B��-��} R�:E=�e�6AB7����bh����O���k��v�&K�pB���2��Z5m�@e��ϱ������[�x����KVzPHp�I�]��z~z6,	���J�'Z5m�D4�%�(@d�`���&�2)B���2'�N�{�1�m�V*��A q�Ͳ
f (�hM����ei��=�g8wT��H	�T��sq��̦�8�'����mEŶ�:� �5��,�����*�=�'�� (�}�D��O��	�1@�ۛ�˵����4erȈ������y5}�g Ɯ�~�6�en��܈���s���rw���jK=��SQ�&�����PUInC�(��$�}�������O�T��!��.,A��7�?���6��Ϧö�D� �&�A��1�� =��|C%	M��P��NRy�u	@�G��#�T��}@S�4��@,,c�K�$C���@��
���!q�k�7 ʦN$T�8��s����i�s���o�7���|�<�	Aܰ�bVF�-�vq8�p麭��h�j�V�k��<�y>1�c��2ڵ����ϳ(1(��B��٩�	�=���8a<�r�`��W���9��P�r��SP����*�#����Ih�Qf�`a_H *x����/��AV�Tz�2���9���ʿ b���P	�x|!���|5̌e��8�ױ�[ZU#qA��WI;��3�<��{�%3�EM�4�i��p��	T�$%H]̋�\�:��2��u���u��H�y�'���vr�+���&#�7�����aYw�ךmHV� �A|��sE��칾y��c ��xM�,���4�+1������`_uT��=�"0��;űO5�/_q�XL"cL��ICSn�f3��$"Z���Pdlt���ϔ v�����d��@#��r�H}�Y{�y����e�E��riKm̔JD������4&Vd1?H�>�
��� �BR���|���<�B��<v��������zYM�pü�q,r���f�����g
>-�#�aQ��
�J,]�[T�M�s7[�k0�q�hz�1����-r<��j��޴�a�7j=���22�q|�9dT�W/^�ϋ\m��/��Þ6[ K�Y*Q���w���^)^{�n���)ˆ��~����ֶ���m%@ֶ���mm�;�����;�2~��'���{U�>�/?_��0���`�1���j� �� � ���tҪ7��b���W_5����~�=�G�$cf{��.��y�"��3$/$�-�y>�:G5f]dGt���܎���%m��������2 >�et�É`|c�N�a����cj}�9�C~�p/�	��e�"�+�"�|��=��B��n���? ��x�w���%$��%ˬd1a�KQ�y�;>��E�e�:��k�%�!�B� ���lO��O��]��uQ�]��X��U-S�з	l1�Q>����@�B��Ҫ�	�^��֕+ʫ����f$M:��nۦ�(�-l���� c�� 1���r�o^lpL��\0����ep��H� �7r���* ����1@3e��d������_��,�Zȑۻ���)�I����*�&��o�����7�g���Ős�:9s�@"�ފZx�2B@*}�t�Y�����'�����1G�80�m\�xt�D�@9ш�%���8G�����,6����0�$����9�Y�4R�2�'  9n��������8_m�g�6`�����E�^� �l<�o�ҹ���@z���Y�oc
`�vIVͤ��T�����`U���~��Ĝ�<��L�Ի��B��ܩ��7���$�h��!��-m��7���E��uI���O�9��0&�l5�d��y��̴�jC���W���~��P�� ��z�w;F�:�`ųH�@v��~Kȥz��#�+(�[SIBeۦU V�88�X'��p8&��RSi(x�r{h����\nwq�K���bk�|�"��ӈ�f钪@3��ܰ�r��>M�ʫ8�w�F	�8�!+��:�y��QEՇ)�*�7�0{%�k�W)�,�j���.)t0G�jT�ԖR���<e�ˋ�ͫ/���sw�*��;Ƕ�m�rG�bKYZU�<����C&��z]_�e���*O���'qV�\ν�}]�{c�.[&Q~�g�2L����$Nʌ������!��2�H�xD+�ebI�9�?q �@eik5�8F�0�ͩc�I����r)��e����/�P��{X��bu����)?S�ͬY4KP5c`q����A݄��s=P�ڦ,���(���Os,�/_����\����S�w���$��ǰp .�A�����'�������v������W?�������_��[��ֶ���A�� Y��ֶ���N�����I|�������ն��_�w���.c��m�� |�[f� �Yu-9
���`m�)�:�-H&Q(GaDF
��kx(����sz�'����:��@�[�_)�^XD4B��ui:�PH�m'U��&U�8	j��<V��k؛X	81Dv��9�������'OE��J]�n��u���H�
��_�Ux��Ӛ�H�@�,nϡǺ����k�S�fa{U'�m���Q쬕$I���߶4�R
Ġ:��6F���i#�*�$�&dT��0��>g����kK(�s�۴����(בǘ����t�2 .ÖD3[.��U�C�c�7e�#�,F��	U�f�����s L�s���I��$�]9P�@M#%����-m�l̕a�f[v��=6�@9+`8Rma�_�Z�q�s��G�]o���9�7ValD�L�(�J�ZV�{�1N�&+�������^+I#�d�2Ye�&�D�V9����/ ��<�c�j�r0/t��%�$�d�3�i@aTu���� `�)mZ�%9L�I@@ �$q��!æ�	��Jߕ�j�Y���¿��+��9���ߵj˷ ��_���M�<����kAM2xQ�l��W�TJ��B�8�A��w����M�M�$�[@_\H6Gv�8�`�7����byv�9��e���6�o��6�K;�rJK9���Os��qe�Ţy֠l�x�����'���B�
@���d!Þ����K�*�K��y��Y�:���k��>�Z�K���/d�j()��9����l6n6_X�b��ƶӪ��Z�oc�L����$C����H�� Z�/�l/��0�pܙ�E���Oq�A1�ݓ�2�ı�1L�"{X�_|���Z����i�m.�yF�J�U��܁YO����5�"S�To����Ž���%x� .�
/�X�O�8v�{�6X8�e�m��$ ��^���wy���������0����zu�X��P��%,�[F���1Qs�A.o��s�RZ�L�GoUy_�����6��ĥ嫔W￲ҥ�n�ءB��	/	��X�n��F�yu�9���QTO�Y�k(4��v���0��*;n�|�x:Ү�{�>{�n�����>��3��p@�2�yJ�Y]���3�V�a~g��]�|��w߿�������ֶ��������ֶ��������?�G�G�Ov���G�O�����i|d������r�YAz+ :[E�>4���K�U�q�a��|����8)0+`Ǣq������;RMj��\N�.�QB�7�n��X��,��@���٣�k>��!��������=��NH�&[��FH���ƪ��p�H�5*0-��B�r&��;��gB�+)�B���`�ys�w�A���
���(� �"���J%��]p&���
����:pV���*I���A K����E�0�N�1V�C�jK� ���T7�"�|���-�˥���݅�0K#Vl9<��b������j��g
�ʇm��bYǦ�� }IT�5�F���ڗ�	k֟���=S��k'�����������֯P��zL��l*I��a�#Ŭ���#rl�옔�o�P9�;V�]��-��� �;�y��3�#���u���Q���ƛ��LK��Z�$R&K2�p����~�
���W��X�j�Hߵj������/���F��)����[˱��e�b���բ�i&H])�^*�Nj}�4^b1��2��j6/ę���̄g>�6ɓ	,�;l,[�HYYnc�$dK���JNڹt�dK�� �9;��[_�w#S,�����*�l�h¥����	�}ksN�]���ck�O�˂�4"�H���$nq��T;��r���l�������$��u#h�,(������1۹���r�8�W��ܨ6�� qiT��Eq���a�{�9D��r��R��&�n�?��Ƀ��8�S�[�����0��T&�b�>h��*t.	
�5��&���K먜���L�U���m��%�\_�5��!d� �Z)"��/�yr97��љ*6�  ԧm!!/��8���^�Nd��q-l$'
��]DN;�Ɣ��+��r��8�-kdOZ��,ErE����`1������1ryΈ�1���29L�}��,�'q\�r�К��20�b�yb]�$'l!��P���jA"����\���s�p�=�{B�<Ι�?�j��~7����,�'�,n��q]����K7W/��Wdmk[�����J��mmk[��~k����-ׄw�ŧ������6m��������y~8����oU|�ښ
	���T�
������X�縆��L�c�� �f!EL7B��V/�E��1��,Y����4(	��k'A�^�>X�l�jĳ�|P�M�#�rCm�(m���V~�5<��Cz���VS���s���34_}�E|�~��r%'�Mm�FXqᶡ����n)�	�,�K��]��D�vL*Ֆ鯫���e#A�mê5�/P��|��fA���R�8K�)^\t�,?����X|߯m�J�
J󛠲{��$'p����J� p�C8sY��u@�5y  ~��u��.-�$2�ݪ�N��uj��TN��p���ZVJ#7��%�F��-HJ���*�h�:�ed��9�;-��-����of����@U@4RƔ,F�`��訪��a�(�TU����"��V�̣�H��<��K��l�p|7���c٦
f����j�:�!Ѥ�`('m�6�l_ݿ�c%VD�GF���ďD��B���K�s����'	
�5�	��#�ƙdm�`G����n:�|�E�V֧\'��ޝO��P�V\Q�1n�:0�$9�JXp����Tyf5 pD?a��ÉY'h���؈�S�5$��N�{Ih�R]!�#x8��0k�RIf�'��M��/�;�p-�������9g;7��s�R�+犥�	�U]a�ɤ��1�^��Pd@0���s�86��Y�㸉��B�TJ����bX�`��3F�b|���ZX(0_������ �K@>?�p��ypI�~KU&��1�C��~�siL���F�(�6O���κJ�9�Ǣ�lI U�/�4�ڹj��	�F��*sp&km�?�q�'%�D�c,C�+`WV�O����7u����}m�#A�Ugd�u��l��\�%b�D��������Z���{M"fk�:�Ox/��~���(�׽����x\�	�ɓ�s��|LlB���8�z?ϟ�s�����G�ղѬ�Z�h����$>3�j���l��iU��i}��(ߝ�P�v�Ī���i��x�-���=v"?@����:��
��}x/#�y�����}�8�h+ɱW�v�V�o��$�&�z��m}�ꥻ������~�����������M��6n�m<cߎ�$�R�_~��;����~�ֶ���mm�m%@ֶ���mm���/��?�x��~��Y��{�a���8��[�wO��4>S=��*>�Iஅ�@C�
�N��@�.Ԭ:8HV�k���S��m��%#B���Q�S>U��#!$UG"E���b�StQ��^A-�������+VXB�(!�dU��$��va�!B�C��S���p諭�%ѓ�O��/�?��g�?�r�>;1w�"~�Ϊ
HD�K�"i�K+,S�ь4H��hrT��.���d{e�֫���/�s��N�y�ը3Pf �U��U������_�L��QA*X3 �$5l{����5SY�-��OH���ܜ7b$��D�U��)�WH*����F0"�\�Uj���Us[���!�OJr�5��3��*�K�� ~#GаT��6eF��}Q�) �����>)����ƅBh�}#�l�I�P�[���u����%W7��������R �2���m,	2�Lb�ۍ� p���r���Ҹ�u�ud�����?'m�2����2	�xy̍�YI<;sW2����(FUX���}U�+��L�	��X-UQfׂ޴qoj��8���_�j���� ���)V��~S�9_q���T�R-Ȑ(�S1}Ykߵ��[G	.�2U�:fr�x�y�q�y3�u'Vg>�s�!+�.�{J���R2��l{dlK?�Ǡ���Wv��[*Ռl;�|��|d�N���罇�Ĉ���B`4���>�ْё i���
����uR��}��P҂D�6������N��z
�$�l��{��X�������>��o����Y�*_.���T��T�?��%Q�U)�����2fp���l]o� �$9@V��D�0�Y���o�k}|�]�x����pr�x�u��V���Nl�J�1X=���=�[�X�~��׾aH0 Kc�RW�`Kr����$�K��*i�ۆ��HW���<��͖D���Ǭ�@PbH7x��d��r����EsAp��������z�ⵣ5"���P�?��뾹ݹ���α������9ε���ߏnA�G+�� 7�E(`?�x��l�R�Ƴ��x&~��+W�X�J��mmk[�h[	���mmk[�o]��@v���������j>���oڻ��t�J�a4˕Z+�Z�L�jy�����*�)Huh9C�!�U���>>����~&*R�����V>3 D��� r��%�X�>�U�py^@9�:F�{>�1e0�c���a�	���⨭x�
G[u:��u����oݰ�����1�&�@?�Zy:ek+4���2�n���I�l@୺��^ �ɛ��%R�n��
���fyu��d�t1��.3�c�2�c�O�6 ��x����wJEC��R�������~� ��3�"����Z�O)7�^����ƈm�YW��DT���0Y�����@)	4AFKa��2o����ۤ���10�����=G%?�2�1 �$�{�"�~�٢H�S%��^/	�k[�tz�l�T�m�n`jy�m,����9 ��2�����.�k�OL����u[gt����s�!�d["��*I;���S�����9�-GM�։��{~���f+"��d��P`�d3 [�bGV�InG�%��K���߭��u�ص�@n;���S:�|�}SlK�-����*F��qm�m�;�����6���]q�h�$�Tɶ���綳��? 9[��
�d��-l[�q�t�M݂Sc���.��k�z��z<D�X'��\Ye�Q��Ma'w~c.�dF�J�G9�$]1���MX&˸���	t#�D�"�`V^b%xI��i|��'�q�s9���ÐP��{� ���5��q��}�*�8g����*�����@�s�����s��(b~	��+zR����[�|��0)[~����	^��>[׶��u��K�;{*P.e.�����f���㻋��U\��P��A���]��Au���.�i�D"��vu��m�=����)V��t��H��x�%�{N�����y3)&GQ̉CrIJ���2�s�i9 �-�蓅�^��_�)���w؏����D?�n�G�M��p?[�3�=?e�oI�T��;�?�麀{����7���G�� ������v��	�Vlۦ�t������T_�z�������?��vk[��ֶ�?�� k[��ֶ�ߪ�������ߊ�bߏ��?���ߏ�~��ղkC�=ć @�� ���U�;y�C�)�J*'Z�6~v�B<ъ{���b���"( ��uࢥr�#j��Y�Z;J,2�ϼ����i�9 �z�łK��䇬cQ�R���Ku�|�'�%W0B�
����e�;:Vc�GZ*�;w�۹W/�ݯ~�+�΃u@|�|��)�i��4 ��q��5�P�N�lTv���F�0'���ER�g0�H��K_�7%!��d�W�w��;(q��1����9 5�@kA�+�p�.�ɪ�/C�]z�}��VX�`�$7X#0� S	���aVUe5�R��g��9��,2@�Td�*��J ��7�&��᭪	x� �
��&U�����VV��{jmVY��|σ˕��e.HYeod�3�B�����ܗkK #G Db}���ƳeV&�J����dW	`[��>:%�����X�F� ����M�RZ�H�쿨0r�\�e��w�	����������vBu�����Z�I��D�J���y��#V(�)U����ش��������Zv�)	8���5�R�d� �;�aJ%,��*�R�Q��)�3�U�d�t�������ח1P9QC�W7�Ty���9L��p�sM~�c�Z�7e�ؾfR�)�p�P�ThA��l�y܊9_�]���$Lp��(h�l�%6kY�r=wۜp�/%1U���V�4�s5��QF�q~
9��#hF&H�tL�|Z4�H����W�ĔqP��k��Rv\d�fUܔ���"�4�oӼ��uAwb�����=SI�1ۅ �K�\��o�^�R�qi���ɍԐ�����l!���Pt���k�_*z�]���]#��$$uD�� �Ht�Rj���n���%�BZ�9���x�%��-������ ���=IL�)����x��-�Y�Ң�N�P��S&?p��{H�ix!�m<2w�/r
����uAZ۵Z�9@:̰��=0�c��P ����Q��5a�ey�q2�盫.�Iܣ�6��D�k 
�*���8w?�{�?y&Ǖ��Bev�V���0]�q?���n��U��eY�_���mmk[�d[	���mmk[�oM���q=�'���G�?�\���UC����]| ��{b�ֵ�.e �Gy����
��K@4�@����0V<�U
~�!,�APs����	�z���1��и���T����5<�1��ߕ��F4��x��a�:m���>YG��#,�V.��C%��t��T9��4�ɓǴ^8N���+�9���x��*丏˨%3b�?pC�15?�u�o� ��0� l���+���'�h�$�  l�[��������_)15C���%�C��Y<��u�:F,�����ء��-	�G3Ox<��x����b�<�o���F����] �ږU�a@	վ��!e�*�<�w���d\W��@���:�A�|h@��f�E��B�c����>�l��T�?�>,�Ϊ����|����eZ���P�w�?p-�Zl�KŃUu m����qZ��z���������q ����@��X6�~l�e��}i�Vf`��.s�DDi[d`�5`m6M��dk���4�_��4��]U m,�m]&��3���|b+�9f�*�� �,��z��	�Ԕ�~�ʭ�ݟN�u�� �-@?�O�B_�x[��9�C�!����4�a�9�J���j������.�J��Kzm�|���m�GZ΁ľ`.iP� t`�Mq�m�5���}ɾ�ݙ _V��2�|�:��p���.�{��1�b�[n������2�u;�m,�
��q�싑=�����G���m
B��9Ӓ�Q_��Ȓ���|��$��%�b��-��zU@�i9�
W�>�xa���x,��o��ZQ���yi6|�$����:�<W�?_�6/Z�ۿ��7��a:�'Z)�ħ(�� �:�f�l�+�A$���`�k�S�m6[W���a��%������>ڸ�o�v׻��k��[o�f����H���F�x͝��H�c�p��'�E��ŵ�S�cvbOU
�k�[�޴��u�6�C�a�_B��Ò�N[R�E�*�լ��j��ɘW'�ק��|{����F���7$k7$�B�f<y���}$=�<����pA>��-�9A����-���3�T?�:��وr	E��y/���8U����U�	�$�	�IU��A��-�> b�(h0k�eI�G-�{ ���0☀� Iq�xM8�΢$��(h�r?��Z�g���|��W�?�y�"^�����Ǿ�jN�$vX���؎sf�LO�&~#��7�=�w}���?���uk[��ֶ�?�� k[��ֶ�ߊ��o���R}Z��G����˲|+>�<���	�<���V�m�sW#}���8OI�1( c�X�H���f�9Δ���幑�{�٢�9�!�
�_��-���qFI%+BfE1R��BP���̐����Jno� �\!WXe�\���`�*�֪а(p�j�����}��� ���3Vf�Ҕ "� %��`&���D%�D���
byxH>�TH&�+Bϝ}�'�dB��n��o|p�|����y���.i�Q �K�<_}C�0��d��OQ������� �bV8���
s�J��Ҋ%Ub�do����g��JkV���U�s9g�T_�ƿ�l� !��n�T?Pk�<���%�a˱�3��*�Ͳ�H����֏�6� x0v;���^	�w������Z	b�fI2!�N�Y_�f���7#F�oly%�a�k	�}ݱ30׶� ZSEX����K�?�$S9nq��2��˒�J�M9�9�G������Y����bZtœ�H��b;J��GX����ȷ�)���hւ��=%Ŏ }eފ-�Z�c���x�5uZ�+U'�/s;�v>ڶ��S�r|�U�����Jʇ�1����U&׊�QC�K{�rn���xr{�L:^+,��3�*s9?��.��(-�\�_Y�S�!c�4��8]�>�/�e猑M��)��L!�u�W9�^ؙ����3��>W���3�M#J���)���L7���2ql�F�y)$z�E?�t�V�TY���I.�LB�l�D�Ҥ�t�B�J����4l��~�������U��'DȐ��rM�v�ۖ�_^��uozUL�\��i^��>)��Ql�cv߈�ܢc�J�C�P�L��}h�(�!yaD�_�u-J�c��B@m��\�����v�S6�HV7�Z ��I֎0q|-���&�G���z���.[Ұ-HN�S%Ȃ~��W�J�9-�}�q��r�w#����b���S�I�-\�H<�<;�l^p͎��#����iX����{�&I��H����̬��g� w�1 d� �p
���!e) ���swW�~�T�S��Q5�~�^�vk���8���r7է��7��O~���m�gܥ��e/{�˷���^�����忋26�w�u���1������՗K�|�7�;��.������A��).*3��<�m���jVSM��2�cg�H"��ڔ�$AP�%ѩM�њ��,��bKc�$G�F�����2���%�ϔ�C@;��Q�@�
>����U��k;���������눨��u���k�B?=Y���:� H�dA�=6�xb8!�Zm��n�pe|��#����&(FVW�x�I�}V>Nh�r��t�� ��j{��)�����G�H�C�-I�[K슱�wCc$���YOx��W5@�C��c����#%(�qX���_���z=󻗋�W����Tؿ%
h��uFR_�5W�ET.�s���uL�Y�F�o#��@w_�>>=��V�!�^`g(uܘ� ^{$��Ή����F��4t.���g}6*m4t�H\�l�2���N����q"����'Ѵ5	8��h�u�f�G۹S�I�\%"�W���o�>���ඪ�"!��jl�]H�Zt1"�A.$*�<�^sW���k|��k����By>����[1Bc���p������e�Ƶ@��	 �J��ɑ�6h�?S���ZS@��ȭ��ڋ~�uÂ0��jOe�9��g^+2��VN��[����uK�a��TM�5W����ً�;)��ʚ�%���?���怵I�@m�;i)�=��2��m]�#)�k�91��>w���<���٬6^ўk��ff����-�~vͫ���S��jٳiL�v��Q�7���Ū�o��1@^�� �H�8�Ֆ��d!]�k5Ǌ�N����L5~�h�����6;^�Iʋ�d������%�Gxˏ��!�~W�)?Nj.�K���|�"%��ʱ��"�
A���������k��»w�Y�| ���9(|���]�Ӗ������	�j�rQ�����߬�Z�^Z�,��3��#��$��i�7����e|��lZm�{?M�ĺ��kӔ�J��ќ|$m���>���ւ���h�O|��1]&�#<���)�Iy<�*v`q��Img*��$��ח���M��7��oR�ާ��e/{�˷���^������/��������˼O��O��|���ݵ_�-�;$���M�) �V0�����%�۶��c����W"t�GӨ��yns�^(4(˫Γ�T�1]	*�t`rޕ�	ĕ���� �*�e�� Ȳ�����S}��3����-y�Y!�l��{$ �P��~���d��Fg��]��p޻���<a�ovL�9uܐbS�r1p�"��m��H�Qb���kCv��v*߯��˲�W�,�VI�:ל��>?"r��u`Ϳ�+o��H�3��G1�c���}#0 R���C������5�ut�5m��E�4U��OE�ǜL70e�}k�$E�@��GK�鈤�ꀢ�x1�߈J��PxKX�d�"t=1�p�xq 5O����eU�
Xo�.�<�-�(�~�U�ĶP�*z?Z{ERD�q�g��x}:nl�s��H�l��q�V9=��1��i-*�5�m���� )��=l�馯�B� ���`B� ZZ��!]�q�~��#�Gm�k�D��R�A ��P���5��Y�v4�5ϣRD�e��B��ј��*�0�DZiL��~��~֫�Q����e�f!!*�QJ͛[�]m-���S[���[1�=αҏM͗ac��˵���h\�O%5㼌 6�o��f����*�]}(uQ]����JE�"�jB��dqT����덊���d�m[UB�J�~�6��
���CQ���N�A�k�չ�}��k��.Ʉ�K��sj�8��������(B��d�WFmx��Nʍ���ZE'l�;ݔ9|_��k`�ߖ���!�ܷJ��V%kl� 潀b	���?��	O#����ս�8=���ӱ�,W�Ϙ�ړ<{a�����2���~C��с�TF��|�|s}W��몱h���s�Jj7���c��%�srⓚ"Y��,Z5�"�^ƌ��ć�_c�:O�]����Ϸ�+�E���xN��\'�\g�w ���x�G�̠"��ݫW�����.�Y1��9���c7��i�^�,Mz��ݫ���������q��^����|k�N��e/{��^������0-�����f��4��K���:��4�λX1LH��7��g� 0�)�$�46��Z�p�0>K �H6z�-P��@ތv��4��d����Fl	���,�D�-�Peg�*��;�	�%�e����ͩn`Q�g�Ҧj�U����<&�|M+�t�6:��:/��=L=���Bb���.�A���e��=��}h�waH����O�R�ypn自����5�ڸ��,��X<�hk��k o*�Q� ���T��-���
A~ʃ#�XU���vn!`�DN/[�$D{K- �@�|�!��bA�2RM0m`���#�]��]�=�p����(���F�G���j�s�-� ���6�����]�U� 5EF��8S��U�#E�d\��ͅJ�ӵń����_���//� -�4*,�4�ǱL[:��� � �� ��\4��R��]��Ɏ��P6ł�ɿ�hn���-C�!�ԗj���Q��jɐ��]MD�@c�r���TKM@�Qu��E�����j!�<L�,�򘅵�jk�@�@ ���,���P�%}h�θ�s���kJ��9t�S"p�g&⽖�Q�ı�v�A[�;�9S.��G�� q��G�_7�O
#��k}!���v"�iQ�h��z_�҄{HP�4���v0v~E�m�~m�}��4��i[���e��������V	8����x��:���{��=�2�6��0�-/�\�Ğ� ?h����[kq]��8�㼿���=�S$��:�9q.�% c����s%������⳥j��.F����Ǣ�@�M����j ٰ`�<�_�H�_��%p�5�#f��/���3�b*Wܘg*-;'?bK�m�5!zr��#E�ڦ��BD�^����㽱�$]Q�h\~��*�A9�����S�G�x�"1u�P����&&��mҖ���=*d<w===�����4�ׯ^��y�0�K!������-noJe��ꏮ�?d��׻Vć�������Q�֍<'�ވ�Fb'M�>�윖��·`-�Ȋ8ViE�H9��5pl�P�'��֯��	bϢ\�Z���љ
$R�  ��/��y���&��	kD~���e=p�[�"�O�/���˷ZLNܴ����"�����v���e/{���� ��^����|c������8?�~��?�{�/��7'�}��G�7%��,	���2�ctYC �,��van���l����6�i)���ɐ-�����M�B� ��-0��"�Q���lIzi��YG�B9`D�bD�1����|���E�@M��� "���W|?׻��R����-�Y/�0
S]��߃5�j	9a5�Ǵ�swX����Hn ��Y�tū��
}��y�5ح�C���w��C�M[hr>_7�����
��l�7tF?Z��5���-������#�|�
ղdk]�E��I5�:8^��n���?y��0Ar:l��M#���5"Y�5��o r��e'"�#*9HG@��R�Ȗ��q.�g���&��T���,�߭j�������QMU�?�?]���1z[ǐ��\@�m�)��\ G��<���*LI�q.�2� �-(Z��U�m�z��d-�j�yUJ̋�%���쇚͹�r�K��d"x|kg��ek�"�9�!X�I�AG����������3���y
��-I�Q��yܨ 8W{�J~�l��Ϩ��m���g$�W{��~`9��b���ϭ�L��j�x>�1�k����>,���my�����h[��y�n�F$KU�w#1�9�4#�*QX��i3��Ҹ�x���b%���\�Un�1 �����<4��D]��1�^��(����oT����Fa�T��-y�u�,�����[��
D�8��J�kN�o�LM��8��l��k7�ǃ�>/�����Czxugsl�Z�l'd9v� �P�H��q���>.��3R��"1�b������͑>�6)��G�� ����^�&�?� 9�#�:����5}��W$O'K:�^$9@��=�y
��%nwr$Ɛ��$����-�j9B�ɟq�l�I���ύ?�8�L�!��a�)��HQ\|�����3��ZI�����#֙�,��u[��	�F�۵H�  ��Ǩ��L>�1ObG?��]Qe]mή���fyl�`Oϩ}��΂w�'k���֣�xgN�|��M�����|�L˫����e/{�V�� ��^����|#��w�e3O��?^��O���Gy��������,�w�}޶����Idp��S �S�2��+bx8��q�Z?�����@���;D�!��3�k��`���
6��E:
�\�n�52��twOb� ��VU�~����lP�� ţ���ޕ�XxI#��E�ǖ����#��h�ᮑ�O ��]��e�ə��	rMN6�拎�Y��36� xF�M键���cA���hOs�Z
QbWykEQ�"|���������.Z���>���E$H�,t^�F�l@P�b�� /���}-�ddǝ���yX��$y;�F���b��9 �X-{�㩴����ƚ%��A�E6<�V�]�A&O���#�-��׹|�&Gv:�
���ѻ"E��K �e�"�fF V@� 0�3Q��0�I�SU���QH���	��\L�1��D,-���J�w<HI&��a;{t-���w���I�%7T�Qc"�5Xco-�3��z+F��H����|Sˬ�����ұsC]q������Pč$b �	eHnwD`�6n�6A�ƕ
�Ϟ�6�7��H��;z�i�WK��gS��*��5�m16�k�j��8��N�U��Z7rL�C�a�s?��93��c�����cGc]�d��D�/�=˿b�;�1��؈8\Tl��G��?��R)ณ R~�X��$W���nm�ӕĻ�V�%�}�6Qs�jǧ�D�~��P�Dk:�/��HNf�;��ީ��v�P�$u$�A�|Rx-�Y�dQ��w��,�xJ�&.�=g'~�h��=�]�<���nm�|=��+)G��v���u���5�}U�@i����w���uZ�3)E�h{�,�����"H�?ל\s�����P��c�)>@>���K��~U���������+ Pj]���&��0���up�N�d3��6�_}���}��Mn�w�3�H���/���.w�4>���bE;2��m}s�B�[��N�9�&
�s]�J�u��M�֒���Z�V;S�س.3f �z�+�u�G�
A����\b/ϸ��h���)����yx�⵴�,ְ҇�q��I��s^��q�v�h�j��R�gQEl>w���ǡ�&?oQC��'�X�9ݡ{5�����?o�7��O�������I{��^���oE�	���e/{��7R���ym0?O�*o|�7l��[���u}��w��%�^�h���3@^��[�V�YTDY�Da�p�< ��6K �*��<����r8k]�͒6�%	�]��c�ά
}7��%B0ý�}����:l�1ۑH� ,2�Ƣa�M)j�!
�Q>�J�T��*+`�������{?/]�՘��v�-�)P`��F��$�]6�=[u�r\�򣵤�����Y���)O*%�� ������`�@�΀�)،���/��Sd�u8M��ٿ�(f�R�P>W}�dA�<��U�<-��O�"@"`h㫪2,Q��H���.��%ɶd
����'�z�YlY2�
�	_����@J� �T'�ε\���Q�P	Q�Mj��hk��-��qp��	�ԑ���ǁ%T�$i�y�.�BL��1���)1�^�X"�Y��`
��<��3��9� ��J�(A<>��QUu�{<V{�T]�sMk� �5�Vy�k�b]�ES�ʹ�OR���:��"�"Qb��(�	W���sLR�ρ���QU  ��m���@ƫ���G�s��Fy��q����}\C��[�$`�̓�TD���n�b�1P�<m�A;�
�VJţ��'5N\��$1 ~��i4��t�*�Y�u�B���YP�DR|M@t%m#[�
{})}R@R_�o�"+��C���(��eh�(o�rj���Du%��+�dU=5���+��*��"���H�g��R�N�e��&�Su/{c6�:OG��wM�v�f%ג�{��UN��[�6F>vC���nT� 9l��Fy\�������>Y�9�43�u�q�ٝ��$֦:`|�8������<��В���9X�H�V�1�x�[l����^�/>�,}��������^����|خ6E�P�q�*m5+*�t@�c,�������e����U�]o�n,��r�qNb]�ua��g�,�6�G�S�CN��,�P��-��$��\ںF*�H
�.���<X0[Y���3�$-m�F6���󹵵g�sn{���i˱����%�>@����4^�y\�o���K�<��MB�Al/{��^��[_vd/{��^��/�˿����_�����M��e����|�<o�������#���ڼq�������������cn��.�i�;q�x�{��#���&o�W�-$BG>�����VFJ��n�?6b3��fnL��6}ؼ�����ag�6�uk)A��w��(��џ,ؗ.�=b�[$�f����7�p 8 �[�	�ǼQ=�������E�����%�͛�n. ��w�f"x�[��X�5�:-%��]>U �Ч��7�S� S��w ��� �s=�/Q�sUq�6@C-�}�7���8&�X�%G���<�\�-�"v��VQ�t������7��A�M�J� aYZ�U�Ld���1�qI�#��(Dp�.�w:&�-rR�y�kiX-�Y q�t �k��0 �T�=^&����q�D�j �����X��F�) =�71����6&F�#�=��y"�ñ�o ��T#�L@f1[#��
0<5�-S���7"�ݔ���O�Mc }��,�i�h��1��Y��^��9up����$�ԷTt�KM�#�A�ݳ�]z�ӯ~�Z��_.V��@���x��������#_A$�j,X�!&�bN
W��<��ɇ��y>�2�Ϧ09�{�~�����-���6/!�F� ��c-�DJɓ���_\����t�z��־}������⩨�8�D��Tf��2>����V{� a�~!��[b�h���W�?�(� X�}�;(=�ݖ	9d&���}NN��+"'��\��D.����@p:�j�4 ���c]��^:��I�{���ud�I�Ź0/��4\_��s�0�}~�.�B�t� 8�e �xvD��nW���ñw�ĸ�K!e�S�r,$�1��N��D��sP�X�=?��q��;��=�~9���x���]!��ېr[{��Qݘ� ����X�V`\{��2U@���)�T!a"�H�h�	
ko5Qx��q�_6V"'e7UI��I���:g
��ND������l�T�D(+�&b�EJ6N��`wJn{V��,י%TOL }�|�8�Gpr# �ϟ�zG�������?O}��������k�@p�yʫؐ�F����糬-Cn�q#�^��8�B��A� 1��+�ﺱ����!�,���G5J���r���y|)���j���
�/��֮=�b
ׯ�>��$<ޙ�bA�x��|1:�����Gy� ��]��x�YM5U�3��u��pu�W�>LK%'�Z�<��a�y��J=�K^�/W��Z��
O��w�7�۠B\�;�g)��C��y��YyO�+֐3�D�1����ckuJ����]z�ß$p�>�����\ac�փ~0%�\C���6��֦�o>��ꌵg�\s�=�'L��^�1 ��54���.���q�ol�C����a}8\�*��^�����֗� ��^������K3Ok7�ɻ��6����ʻ�.w��nC�ȸ�Rv�c��&��ƱY�-S��m�Ǳ<��tHJ�M�����1j��
ج�e����)���	z�7n\�o�t ���s�Q�kk�*]tb�8'����HƤ��&K��K���ojR	2w�ހI�����Ű7���[�.�K�� ���;�S��"X�<�i�F�Q�&H�XBbD�H�j{�o��p��Ĭ�f#���$ &�{�SX�Ù�C���]�ę|ʃ\��mO��kȈ|$�z8�Z.��ݯ�+3�r�sjj�e�Kn���C��2�
S�~��I�k�\�� ��o�6�
����w�摀
`	�|��u.Q���E�5�|�c�����%�'��{�܏���<�D�HjΈ�-�� K���hO�'t>��C_@�[e�ƪT8@E�+�BL.?:0��u�h�%Pt]�r,��9�LL�c��HpH�>�����uAcXW=#it���p0*qT�B���p�a�Y,��X���%�v))�J�<sj} �h�8+�<�u���ߦ�8�ʉ"3Z��؉m�ׯ�י~�v~SMa�8�vR���uƈwS��su�����܈-�����j��Eu�Ǝ)��vrՖ�ZT�ڗ��ak�T�&��������n����k��%o-����f�	�X�9�eE�I*!3Z����j��Y!�=�>���W���Ѳ��Ef��S����5%$f|�D˶�5wLڨs��m^��܉c��m�.��Tc��u�%��AC9~��C.�f^Kx�����A��,�߻�S!�_�5?~������kԺ�0���"�;m�'n���T�E���ʐz�7�����Xsk������e$���"�K;�� ���Z�ދ�BFd&�Lmx��|gkz�����_�{�czz|J?�яH�� Y�Nw$�*Y'�L~���*�W���8��c�'֚�_ʳ$�֮�#��T��e�
�Z*�ݨZ�yZE�<�B<�4)$S��r�����֏���;TM���a]�u��h�6~���2�K�;���_A
R����;La�4���P��Zd�g��A$MHO��X��:�m��w���М��0�����e/{�˷���^������7^�v��&��F�M����c׵ݒB��d�W�<�������i��ʣ���|X��	�on��Ĝ�o�b{@��T(�(񝹡!��������u�eWz�E��V�� �q!!�k#gZ�0���Nt�����A�XK���[��Yl~��L �,���,�,-J��Mb������c@�0e��.�8"�I��ᴈ#*V�WOH��%�Q^f��m�:CvHi�9s�����+�5f^,:X�rM��`�Ir3n�^�+�xYk[D=��G\��u��mM����#���
�'1�6v�TQ,~�8�1Owqs]��W���P��녾����S��cm4�r�N��#�7Su\z#��U[�h-	�7 �E�D+$�;�Խ�
���ڌ`o��Ax̹&��V3ñ��� L.�[�|�J�2��ܴ(�-�#` ��h���c�Ե� �U�D��G�J""hy��cp�%����ϫW�w�NE%�Vd��c��D��9�x+rmv +�i�ﮐT�2E�ߥ �]ƨ�G%�Y�1��4·月v^��}�2s�#���M�k�k̊Pj0�W�D���*F��Cw(�H/�WQЇ�㦔�6��~��M��dQ	1rE��cX�'�q�UZT�M�	`�4����%7�0]ݲ)-���j��ҵ�����r��e[�@~ּQ]���tE{a��:W��ꊢC�Ϫ�b��O�8�:U�)�-���� �'}_ר�k^$���%���`*�m�WYb����<�Oum�ws��'����~��_�{�]zx���y<އ1֛-��)����&x!��������Ԑ�L1eG�\]�	*�1�z[��]*3�գ|�_�2�9ؚ���,�����ʧ�~�������o��o�/�����!�~xM�.k��I����qd=�+�7��4+�2'Z{Ƅ���aPB�U���Ξ)��L������c�@`��4��+H�BgS|���*R.v�n��c^���3bޑ2{r�q2gຶ�`�yյ~�Nk�4�3�,�@*��:?/�����ym�@N'�;GS���5\A��\G�Ed�Y�\ώ){��ӓu/{��^��[Yvd/{��^��/��6���p�kک���#/l��m��YU�s_�>�9�͛Y�D u�wz�� �#���)G7xm�pS��mh7��:Z�[!C�9�I�+.�^�$�r���{L��Z=*CTfW�)�$mץ
a[�&mh�/Zz#��Bf�9� 1Y0��6�7�/�,�`��(�ucmH�� 3�5ӗzA��Y�H@����Jj~c���IH�r�<X�\&�u�Afn�?U>��l�*�^�(O|۴J:�<
w�(E#�
h��P�ˀ����;��C �A`2���9҆-�N��7X����i'%����y���G9_,�4��,B�j��o��兟`�3ͥnl��ٺD�Y�D�C}ߓ��i+�/PR}.�QDS�\�AU�&���@�����_ĉ��C�pS�O����l����������.Z���"H"�G �%��."��p�HƮ�$�zP���B n�� ����+��������иP�q���haU�λ��>��]�@��c�H����X N��^�3�v#9�M������*W4v4�6s=��R�sO껬n��Qm�>_�Z�qR�8f��C�I��&��J�8�Ԏ8�+���g���m��E91D�5V��a�7āΩ1�6�5��B��vS��R9Er���<(��e�]��{$.����0�1����'��(UaR��~��o���7��V�?�0��J����P�)q<�
	��X۱�JW����4	z������]z��F�'�?�"���+Z!����rR�̞gcN5����Ɉ���
����C��^��1������l�GH��Cq�h2{ʮ�~P@n�Vui�,X�
�):ݿ�z�%��ʽ)�_^�J��|��v�gڻ6 ̼�����Â@����p-}O�'�x#І���eqeV�|B溗���^�}`�ZA?9Z<2P�zh���MI�˕�޴�q_0e/�>z_��&���á�e	�]L��r���������5�y�`uNx��&Ӊϣv}Zop��/��	5,.���17�1(.WĆ��l�̽�e/{�˷���^������7^V צ��q>�W�6V�>�H'�2 ���6�<�7؀0%��������H}�gg	Hɂ7���ƔN�q��pK)*+��L� H��<��i�m��R�x�e��K�����ZE_3��Dh�Ƿ0�mvlv[�Ʊl�y�Β�2�1�y�+�(���β�R�XU$��&3����Rl�M��	I8Z�?�y锪�m�%{o�\t-5�_��@� |��C�~%M�[J$d�Z>�5��B�m�"���i��75@�ȶ���擓�C�%�{2o��ȭ@�e}'׬��a�M,".�z��}1�%D�2a�
��r�t��1z"�\ |�f�爴�>��|�\�[�95Y�o%�0-P�Z~�LD`Uƻw�,��KI2U�6�ʀ�k7�����G�I$%����b�G�#�m���6�7>�D���ɯG7F�k����� �d��H�qM�|�D���"١k�qu�j�6+���<Y�?����en���XO��3��o��`ok�;�7���o�HC��Fզ�+J�H����cY
�����\�*v�8�����NmLuM� �F1�*�6�M$y�mW�'ޛ4�u���J�5�I�(�����*�{�z��I��������U>˿kN��,5�m��D�k�͑t37M!��-�$K��̎k��@t�l�x���R��}*ye�̊c4+���ȟH��������nI|S��_)5�nV�d;Nt=q���g\ه��'���^�ˣdd�]�C-�6A�E�������\��=x$QZ��|��>�"�~�&aO��h��1��(��H���|�6�s�ݽb����V������3Շ��Gg��R<lؿ��<OZ��R��Z�
|.�E�B���9�\��g?�)��@�}���0��	�K9��x����ƻ��_�[��5'��{��R���s@\'i��@<�?�/r�ZB�����Z�U)	��� H�xR�'��i��-
µ>+"xC���?OFK�5m����jy��4q�>w��R���Gg�5�A`��g����W���ʠ�|_a;1 `���������\���^������+��������7�y��� ����h��=��)Pi4� LF�w�����j��A[�MNp�͆x��T��p��B��@�MJ.zb���-�
��ǖ�7����֣P#˚��E�9K�T�M�9b��M��c��6'	�؆{v6R���F����E"5�4��]{���*�E�Cޔ.�����j��2Q}b���n'ԣ��Wt�������c]�������I+��y)�� m�-�A=�n]=�1A��l��J	��i�`>3OBn��q?!{�˅��y�C�Cc�
80��?2s}|���ئH���HP}��Z>�{ccQ�:Ɔl�Dh%��R����8(�C�
�j7�����PFۢ�;�ZF�������d�@c�� (�z���T�4��"Zs�'~���wڜO��y�#�c����� eTE�Mb�9Ƣ��5D�� $+W��]��D`�(Zk����c��-j�ůEצ�mE&Ee�Ɛl�t�"4"i��}�l*�(�H%���n,x_ĥ�"�I�ы׆��d����}	�VSU#	���#�-L]�ej6D�l�bDT��'R-�Mtn�S�gl�[��S��㬁�E��%���ۃ���(S�ͦ�e�ڡ�K��uv�e|�yo�gZ'�G1�=�CT�~AQ}�n5wKl��^u�F������f-��(�;�[�w�>�qӎ�é�i:_G#A�":��������p�������b/>����g,��A�Ž�%E���\oɅ銥Ֆ8��w���`yA�����:�ޏ
Ck�l!?�r�TE��iN�c�>� !�!�zxE{+�D}����{��s�c��'n����;|�chd���4=,����rݩP�	�O:f����]���Q� �1�[X�5e-!�,c�Vu�@.��i{;]�$�dj$!�BD�2T�u5�d��#hd��6��f����Xz��Ίϫ�}w 	5@e�u�k\���u�����p �@�0	�Ք� ���|L~�e/{��^~��N��e/{��^~��)oD�Q:m3zyy!�ʛ۟9 �7ܤ��Yx���66����7���Q�7��ɠ뵘",I~��n6a�Y�#o���AJ~.%������d��cUU�Ge��5m���7�7־Av���)-u��Ǻ\��v~ԅĎ�� ��c�����;v���m)��� Y<'C�NH���y��DH�U$�d���3 �#f?��� �4(r�X`��^_*�Q@�����٠_[:�A��&����q��0괞,�~������T*,EI�v+���U1T|0z���#�Pؘ��|�A���0��|�܏W�"%XߛG�0\�~׹�,$�G]�yL�u��vI,��{m�Gd!�6�� �fp�eaRl���6��:p#{/����d�˸�{(Q�E��|��e]�Z��x<*D��FH�gb4v�-O%�n�� ТDд�Tp7*bbu��1��@�M��a1r���I ��-�d�4�H�vm�˕�/��ҵcY~���C�S@��1�y��5X�y{�h�0<�٭U��˭`k%p1��"OԖ ���@�C�נ�(�Tk������g2=�G1_������f�ض�5�Jj* ��ǖ�Q
��w�Ȃ��	~I9��Ƨ�-�>���2��mg��4�'*X���g��$E��.by,̍_7#�'�S�2���G���x�V7I�7��n���+��A�ĥr�DҊ�]�ͼ���ek%f�m�}׉$4u�A� �u$T��U%�☕��xv�	�tPuh�j��Z4.$O�}dO�J���������e�g�Q��8�R�k�?.��
��y��;P3�V����S}qH�]�z�ʦ��,��@~�NW����]���E)�{�H���nӇ<eP��N�<����f���p�j$t���A&���W����;Q
+,�l�i?9r���j�`���UL��O��ϲ�<t=I0���մ
���Y��ς|N��}�봚j�A3��A�������۩�:e*�H�t�f����TF@N�x��z퉳�q�*���d��m-��u���jc���d���Y}z�oS^M�:�x�XMg���o^��[=ls{��M~V�w�yq��^������[Svd/{��^��mn� �W��R�'(];'@ �w{nJL���1ms�q���M�%&�R�&P5�7�*Kr�����%6����/��׵�&�0J���Z�b��R$�F�q�L�f�7��ŹW{��o�}q���XP)R�͢�&O����������� �`ѲXQ�`1@��)�LMk�.y
p��F f��^��Lۦ��R#޻�k�%1��Z�F�2	�\ ��#B7��#�C�,U_��l�lKd�ق��5M�k�:�ZMhCR �h�T-nd)���n�V�,��d��ߑ0�����F����%1m1��@��I�Xq��F���><��M���K��n���sb�����@eBj]M���"ɔ���>"����婀�%��G�
����9 ����\������z~.cTvS��DL��v�J�&U<M�ob �8~T�D#����6Xo޼a�ȏ���c�\&Q��~�m�9��0@���	����7�E0li��R�'*v�6�{�H<�U��Q/�!��R��|�<���F�)Qu��]�m^�@N�\ jG �l��"���+�0���8��Ol�h}�s���o����Ȧ���ׇc��Վ��-����9@���N푨�}��g`�V�K�O��{W��J�i[	L]sL:�6�׍u���jWF����c�$��Qmu�GkQ�kԸ������(��E�Cת�H��vL�꫾)s2_�7Z����REu�w�@�W���eH��c�s�#��c�3���sL!�@ڵN��vm$��z�x��k���������W��]�}{;�"R6V�Ǌ������{�
�����"�]ߕ[6�&}��1�`8�$H��n���5���4�U�5Ucv{��j��-���!	{�8XԼ�*π���U$́��5R=[�<>�����{3�#�^R����	�e3V�K�i7�+���0�<Bf�����}�}h�s~�.R&�cQ����a> yG�=(:0��Ƽ�-�)������7��T>�O���km�L�4A^:��Ր�ȷ����e/{���� ��^����|c�LD�}�73��%�z�:}x|Jk޿<�6F��1MWVW-� ��Y�:DJ_r�t����M����7�ؐ��)�Oy�o�D{���xy4���¦�X����K��k7	�S�$�2'�^^,5<��y�L����?h7�<��2_�����7ɸfD-�����z&���"�=��؍��cs{+�լ	������2��S��P�B� i�bW�ҡo�uUySn����c��;{�&�`�p��bvyG�O%����@��:_7*�Z��K����`�6ϊf&�;���5��IG[�I�Ba芥�2����n(��t4��Nε�`3�\�P��[4���
�
�����|�d�8XBʟ<�s���xz��h)�6n5a
�������>�q6-�3P}�8\@�@�c�&����#�y�}�ln ���|�߰n���m`�P�#�F	�A�\^�Dh˗��^'��  ��IDATw�U�_u����Y���a_��"�(�.�ɽ�^��d�#z��2p�q�kXu��$b���6�_����(؊��J�. T�	&�=_,J�q��|]��?X[�f:�[���� ��̕s��0 �q*I�eǃ���"/��&-_}��kRI�L�xp���ߥ��m�z�����q�sƨr�K��"D )"ߢ���r���kQ;`��ߟ���9%0�@.�������r#��1�"��R�(����`%�,*�>�]鯘||n<ֆ��7΃9��zcN�d̪��[G���'��������$����@)`œ$�F�D���nW-�x?ZD�]]�R�A����#�4�j7��;�ƹ��ji5l��-*`"I"R�WXS�nx��Rw�T�cl(��;}V�J������b!x15dT���s!)Ep����bx�}�|.���ګY������k��a%֤��s�J�QC�TR��啩�hı���W���R�#��`9�&xy����Kw�Z����{�����O����%�8��K'%>7�Ē�� ����l��l�l\�vp)Xa!(��$��ʱAv�P­������\���>�A�����s	��i�<�"��5u��g?�Az��b�j�r˘ee,\��g޹乃ѕ��E$��m�Mv�����\��kw�1�2	�����:��e<SՊ�� {N���Z���;��̆c�޾��nӆ<~��rz�i���Ҁ���u���g�v{�Z�Z������u��3�x������ty~��@��p���Q<$��ܟW\{��^���oM�	���e/{��o� �7@htK�Cs4��e� �� ���#9غLf�Ck*D�+�yg	bk𚀼��H�6�6W�'JNf#0l��RIn���Bg��{�O�Z�PyΗ��:���"��_3�&��v�K�[l���,���l�
�;9�#�XA5�ٙH����$Z���_���h�����&;-]�[���%/���I��E�p! e��U�d��֯;�C,��\���z�0�KH��?��̛��O���k�]���w�i��y��#�c��B��ؠ��XM�: ~a2Yڇ��@k��� U9�<q-}�-Ë%1�����u�<=�� 90�S�_$���0�=���Lc��C:���N��C���s��z|o@�x=�i0�K* F�G�2R#4�^���(����W���,cQ.�1
Z+�;F�~
< 0uGA��ӵ����(���sz~"�G$GT�h��TF	_k�r�LQ�8�)>F��v�U"������J�1�KQh\Ky#����8�}ӍPm5_Ug��'I��R'�U_���zP4�}QX���y�
D�)�z�Upۈ�J��8j7�[O���O��n"Q	�~��t�����&`N����5�p�hk�M�K�E����ږ��{k��Tk,� ���q>�y��x�8�Me�As�mj.�-{��c4{���ɨ��j�ml���c����5�2�����٫bR�E+�x-Ŏ���ڥ�W���zm�P~��a����װY>����L�g��iU�f&	�����uFt�8�d6��3���u^����''U��I)"�%SON��,��>�~���D�/����2�6�dm(�2�:Q�z_g���,�e�d���T���l�ʘj���/0� ]�{P���9)�[)K�6L!� ����ɕ@��~�d��B��y�`��E�E�m'uu$���Bbp���9<�!Y��`�DT��!���y�c�D�T��!�%)b^V�����y�Ç���30x
�x~(�E������]����e/߶� {��^���o� BԉQl�5�C��`I����{�f� �&��6�Rd0�~2 ���E��7vT̫ѵʬa.F�����-�T�Ǥ� %2G_�$��#mU��䓤p.$�|s�m�X ��X�H]��ȫ��}���ф�G�|�[*h�b-0�ظӡ\��p��J�48�+2S� �\��	8��2�f���v��I^�?�6XKW��⅟ *Dt�[K,)@j��ͷ�=�ߐĢE��f�癊�e��1ݧ��)�A�LDk�5Ћ�.�������0x�5ۍ #�&�GЉ�ew��6�K���_/3I�V��p��	�Q���s�ꗿL��7@���������<��-��΢`�󟥗܇�_Q#`r�`u>�Y�'tu0�谅D��5r�h��
�c�SA��x6U��t}�V��A�p*� ��ER�&HV��=�20R�j5�.���R���z_�i�)�Qҗ�Q��w �X yDxM޻M>Ad�1�N��q���r蒯O �%R��	��y6;�!��u�o���6%�#��E^W$�_�J���W�
�W"z�8�W���J_�0�X@!���VYV�ݧ�z#!U�(ޮ���Y��,�`	��k��%�ˈD���h\(7���$ZF�~�9�jc�Oy��5HuAu�x�$�Q�s^�ns�HP4mU�E�O�0�s!�m^/��D��5n��LTj�:��f:�H�H~���ҍZ"�`�=��J��+�k���c�bO"(���ǊcL�E���?�k��î���L���W�3~mT�D����\�,����Lc4��g�e Ӑף��D��}����R�r������nQe��d|x�r?���������&��n��R{����H���|��}h���d`����^���}!Q�v�yc ;���p�`S�A��ߺ�Xk�`����<o��t�f���}��X��K8g�7����8�q�#�*�&T�c��1ŮOךu,�1fiUmո����e���8��o%�>y���t��9��C(T�����N�ħf�[R*���Jn� ����P�LKzyzN�����'�� �6���{��^��-.;����e/{��6�ؼ�!).6aC_�$���o�EO� = �޻~2ȋ�@�s�\�Ѹ����vz�EZ��cV�҃�E�"Wm&+��z��wd9�4�����l�=�[��蠘�uw�|���m����X�M�i���@d4ܲ8Xo@��xΐ9$Mm��ƀ��"��D��ZҸP�����?(� �e��A�k��8�-R������ã�S�"/��g��7���`<R�?Y���'�Gzz�˛~�D���w `�j�1F x��
����K���ݻ�h�q�{��D
�E+3��䠼eL~��ў
`h��^,�J�͕"rX<��Cv��	�s������O/��> ���6��/黿�/���!�z��-�����>6<?l�68.�M9�� 	ȇ�D�@@��5�G�c�6:y��XX��4�SH8�i�,y�l�d�Ku��P�
���ES7��c�6������\פs���&b[u�b#@/�F�}V�����c��$�߰zb>��m��Q�e�%J�3���#Y���#���(��%w�����Q���r���Z:�$�j߭��D����T�.�c-�k
�%�R������C�j�h<(���I}�5�(\�BVH�9��t�+"#�!�M0��9^7��r��z"�ǨH�s-��d���	 �n���n�Tz/~&�Qi��Blc��)���$孉� ~��|"oU?�E1H�IN.K�ǂ*��o�����(��G��2��r��(���V<�&nZ�"k�ߋ)~`�e���;7"��ﺒi�[wvln��9�yP�5(=t��{.WeGU|h���Y)�VOϗX?pG=8y�>t�����Ib(o/���~�zBnsSQiP3��vDñ�wu��1�-���rձ�{�\U�m����ϗu��e�fwV�RY���ڧ�̨g���I��]z�ϟ�ȭ�ϣƮ��j@F�Y��XԻ�q"�����h��G�i]K��鎁3�OyFښ�.�5�[}�zm�FA�:�����,$�GS�<?_��e��'K�!i�����e/��e'@�����e/����^�w�1oT�70& ��}�p bqɢ|]m�&��HA1�G�;	t��a)m�����ϳ����͛����&=q���%FLv�r�l�D��U��9�|�N^$Sk�n����YS�qV� ���IK������Oac�z};֏��d@�<�o�/F重<�~0/�X���Y~ ll-�f碏�����i�`�5]�O]Ϸ�]�]m��NѠ��_i�����}�t�O8n�Y>����aH�}�.��M��c��W������~�E����-�yL�?<����+�/�_��/�L_~�m������������L�}�惘�@'��JR0y��'���+U"]�d��'<��ߖ�yWz��f
 �=���y��?�8�엿HMߥϾ���������^}�;�~D>	K���
�E��j�P�y��󲂽����� �e�`��K%P`'BK}�/�-�ȳ�Q��1��}�������"ZU��$�ugf �-�\έ��3�vEp�8�
��Xp	�`��RN ��!��-��6e��^$b�q�I���| �d�#�i/�mm��ݩ2�6��e���)��jhQ	���4[�-��j�j�6�h����<I[rIJ�_J�z��u�>r ?U`Q}w��^���l�1�_���/�L���G%������G;���D����v_+ﳲҲk�d��{�|wwܴ�L���/ʔ	hS(Ж� h��`!`�C�׉?QI�&�Z�ӛ���f0������k݌{�KgRahE���r��sh\a�Ȏʗ[;��,�MC�q_'A
�8;�x-���c�Z?�eqN����׉V��8[�&��>��%f������}c�� ?d논#�V�i���"y ��rrXDB*���o���l��0E믓i�������6墕t8v�Yo8�>�l3\�󓑾�m�6Y�g�5��  $�ƺ�|R���L8��k#�1��X�T7�s��rX@��<��:ۿy�F{����e
cd���ʤ�21S3(]�Du�Hos�;F��,���[>���	J�$����Z**�����=�t�?O��/�����������Փ�O��d���0����X�N��Ɵ���[�&���5$�������2����=s	���^����|��N��e/{��^���M6�m�M\�(��<_��V�Q֍jxX�`gM��
j�Al�ŕ+<���FD>��x��uM�T[�Lx�d��cH���ϛ�@���Ȕf+�'钪���L�rl$~j�rKPKf�\��}� )���{]C��F�`���.��1<Nr�8�e�1D��!q��O�d�4xb`�@)RfO��:whm�J�25�v�.l4jQ�g��M�G$��ȣ��M�h9��HJ�ik�������������H_�{����.��_�U���]�������{����� �W�ߧ�������'�o�}N[��}���c����E�2���_�5s�&�Mؑ4���������M�~K������%��*�������\�ǯӏ~���?���פ��7�?�Uz��]�������k)Y�q�yF΂dØG2�ˋ���D�J$�?J��� )�F���ʋ�m�n�R&ؼ���k1?��qd���'x�\���?�5G@�cn� 7Ar}���Ht�f�W��h�Ij��A_}/*Xg�}Q"�Y�T#.#Ies�Λ[ە�z����3j{�Ui��W�#�q�69"��]s�p�5W�!*w�*g���:i��P�}���J#:�6�\�� �ƚڿzL�/ON�^���9Wn��D"������5Z�Ѣ�s�PU�	��o����n���D���b�4�q�$��*e���f\F�n-����U��cY|�A����Y5�h��~R���y�P��
�H6N�<n��O)?����s����t��? ��\֘�do$�d�T��JJݮuۻ����g��n՘����V�F^7s"�b��ٞ�	����)dc�c�����ޘg��ץ��D�>�×4�b�ו[$E����������{�O���ϝ�3S�L�c:�h�j�|N��FPL����B��.pSs3��j���q��>���k��@��I��P����Ϫ�����^���)��vAm�g����R)ʟ��u&���gB��U��R���]븏
�2汎�� f��IU����gn����J�E6$E�'��UY�%�CbΏ����pL���ԭvo �s�Y��k�-}{;������e/��e'@�����e/�X�N�t�Ql�lS��G���2fDX�K��L���(\l`�'8��U�=��DYb����������M)6N��#��}�M�fhl��z;�$�!1$�.=��H��C���D"Ŭ�Z��=�=%�l������m�R�`�=�ugPS ��# �ҫ�6���Xɞh���*8�zT��z��d@�����"i�������/}/��(�D�	b�����X"�a�1ٯ�����+H~�����/��/���o�<�пM����m���q���H���������Qaq]���r!q�����/������㔾������qn�đ�~i{Z��H������	p4�Z��4������L�jJ��� Z��8�?�������J?��?���GF�N�	���?H_|��{h�WpξSB�Ţ��c*��*� �aNX�̜���t{}��Kw�A���95�fk%�B��^X�#�m���C�P��*(��V��� �
P��`>-��M$��e�8"�i}N�Gj��M]�-���h� �^'a� ��ȷ¯�_�&r�zm,W;n5 ��7��g�-! 8*
Ц�k�k��A�M��Z��D!��"L����*����'��G]���7UV�몊0�������.�4�mN���{��	[i#���[���V9y�?
�3��p��W_�о]S���Co�>� C۳/���6�U�M"���Ff�^��@���Ѐ���Y*��c� ���A뮵\#��<F���z l:�xTo�)�c�J���[J��cx�%*�� �\��J%��h�@�q	�[�-�֚D>�a���i��QD`D��{\o�K��@��c}�"�'����J��O�e^�����Lu k<F�3O�B� ��^��槥K?�mxv'�m�s�x��Us9�ڬ��rs߮$H(hK=Ȏ� �2OZ��K�'�|Sl���;��f�g5�.��<����no�,E�*۫	�l܋�-���Pj�?m�I�]�1�W*A��ֹ��Z�j���6p<_-�����$cז �Ԛ��g��]��
�7<�aL�°�=�v<��f۲]X��l���2t���ҋX'}l��,���r�N��*�H Y�ծlk��d�ԣO����:�I2�縯O�3�(�q��X9����e/{��/;����e/{�F����I��uWoM}' "�E`���D�ۨ] ��#���֐u�#�	�@R;ȒĀ���Z����k�;����9Xq̂�@Tc^�%�x� JQ��|��T��3a��<��q�"Qq>W"hqH�<�_�j�&��A�Nfd ک]��%���Gz	���a.v+����ůvG�d��\+��:ɔ;L�9O�7�ɲ�o�I�'�� ���y���ѣ ʅ�e,�)�Rs}�bIJ��Y��*k�k���-C���DCwH�^�����?������?D˥�����oޥ9W����N�~L�����d���w�E��rN�7����s!����;� ���2�:����,� 6!Bx!it��6�kE�ϋGq�̛3s�]��$? �������?��?����kΥc�V�ҏ����������;��]�������N�7'�SKY��[@�1y�Z��h~ *�5@�(�;Z����b�CS#���S���oY�Ȫ��@���*G6T1:Zu �%��-��Q���%<FW� �]�Oc�v���@=�Ũ���,1�>��O�圷���^е���F}O���>2��^j�	��P#�`F"%*8`h�_���X�k�X"�їxė^��I-�?o�g}���1��m{WΩ�q�?�E�G�����2��X�j[���A��?��9_K��ԕ2���7�S�}, �w��qPt��6H���e��h��&�Rnǜ�w
�Z���H�ɭ���݁DV�Ńj���aX#"	ҸB�HW=M�q(WZw"�JZ�D�� Q�o�7
�T�뭽�8ѣ1(�E�T��Χ9�'0X�I�k��� ���䓅�=�E�#H���5��S"OPy��9��)/�2�י�g)5k��G��	��gn	�B��4*8gS�bY?[N((�SCc��+DWO2u8蜾�2�c��$m�̗�y��b9�Ю-�c��u6U�Gsc�gL�}�3��kgT�|}�q� ;���3�Xy�x��8�X\��˳��=�I�2��$�����dG�9Q����-�e�CB��-��ڪ����>۴����(�ڒ�D�sq����6�1P�Ɣm�5i��(�8�;g��֬��Z��e/{��^�]e'@�����e/�X�f?��76*��><�Oo_�I'Z0XD.��4����.:�̼�W�y�}r�~f�7yW���)~ڽc�W��@}��G�?���6	�+��yU��t$���"),��\l��,���|�INH�=�::(��#��� 7�&�v]N��	V5PL9A%���-ʎ��Vy@��}d�2�Zv���Q����_H!��������@A�̳y�����-)�y�c
�
��'�3��� a3�Sz\^���j9�4��?�E�f�Ѷb�-��啑���Ɨ�x7'~�`���VZ�n 8֬��q��� ��������������qҦ��_��o?3����b�۔�V{J�W��՛4�����?K��/&���%�ɟ�	�@�É�V��0����SՊ`-��/�ĠNy~��V���W_����tz8���]ϩ]�,�9χ�\�#I�?�z�0�y�����O~������~�w�����Xq�Η3���`ő_ǹ�"0�|~���,�G,[����{�*������7o��_}����d�Qq���.U�ЦϿ��\�3��(� 4��V�7k�e�%$[���#Д�� ��ӱB|x�P����/G�n=�M̯!�g���hu�]M��{*���ɳ	D��\� ��zE��o�Wb���_m�z�ݎ�i@���B���+t�.$ PdDĲ)O��|*'���;0w ��5���U!T������J�5;�!|;FF��l��3�Z��IXW�H����DP��mm�_=��[�}�4!��~n�8t��fL4*�l݆���^�'d ����n(y��f��R��ļ$�FV`���Q�׏򘛖b}$��u�*�T
YИ�фM2׼����X|�NNN��qJO/O6f?TBݩg~�����4�i����hۓ��i�-b>7�K�-�w\f#Ćܷ�����1�g�_O�L��&�Thܞs��d������#B�X!Z֖��:WIdt���b���}����>pL�^����	��<s��\ �&��a��J"VU�6�xV������`���ø��'�۬�zΓ�+������ �x�k>r�im��|��{��k��^ҾN��#����@��|��]z��u���~�,� ����Z�V�2:'I��i��߸gK������5�xP:���>�L��U��t���`�O��ڱNA݀<o#�~WE���J�>ACr^�5U�E�e�?R�-\�J����G<�~>����<>=��ʞ���I��L�2�Gm�e������e�o��b��S�|O����1_��}�}^�/\�7׌g��h��/g*��>��q�E� 7��"���5>���
�7O�k�2Z�_������/�+X��~1B����k��[�^=�5�@�k�ϼO�\w;w.�b[� ��}���s-��)�e/{��^�=e'@�����e/�������7m�0D"sD�5�鑳�c����`�Z^����3e��۶Q��)�j��7���a�	��+��g�pr2ѐ#�N���(K$]���K��YN�#0���['bf ���)_�����Z#]�&�9B:�X6庘�r5���
��{N�BD�f�q$р��E �<&��5��j�R#���EI�{�$�,r	ES:��5�MEU������^d�D��\iA^\�5�(�y���_/�>s��̖#�&H�d볆 ��q�\K�\�4]&���Q�)Ni�o�]�'�����������Ny������!-��N#mf]Y���9����!�<`bv ��f � ��<��вv2		G��������_���|�����IoK��i�,� �8  ���|~W:�y#xk.��0�Dϻ����I�������rI�Sc �WR	��!8�jĵ�E9��Y���&�V.�h�����ע\ � �	�TTYO���t'�}�'��}�M��Y7�*B@���E�M���-���)�\��^���1��F��Tq�۸�`uuΥ��(��)v����//O� �1�T�QT4�+�VK��M��	��=Z�*�g���X���0->���z���
���'��ukS5j���f��Rg�(kW�`�i�)*?F���q�r�6a�*[u��W��/ Bj���j��gG�Pɢ�ڧ(T֥(�⚖��.���.Fʤ&��I�د�׺��Q��U$w�ys�8���5 �g�G�Q6{QqT��W���9X���+Zq���~k��[Ib�^�W��3RP� ��\�bӁ�v(m���4nH����uk�ɩ��ۘ�k��x7���T~u%_�&7H�o9rMQ�Y^O7�~��W��˱YqĎX"p#���#�G����\�YV�����_|��u�2��m���8_���њ���: %��0M��$��uLvY�wQ�a���ɏ��Ǿ-��4��Մ�F�/�L���:������ߔ��ͻ�����C�-V��Ü� r��-�'pp= E��c$�y.��5W�򔜼�P�*�XA_���z�i��9����5�C����WgjI�Qx���4�ka�����Dn�<|�@��\�O��YyI{��^���oQ�	���e/{��7RFW t�6���7:����	�S���A���N��bY�j�6t���f�S"J��'��_�A�&8VVxU�� ���É�	��{yyN��K�.�uF&�>.S9���:���'��Ebx�k�I�0I\+��%H_�1� �r�$O��ׇͶ�1����f �E@�<3#�l����|�й$��z[�qK�������LQ���>7��N޷�B 5yQ�t`*ILW^����;_��\>c�fq�K~�D��� �u�,ՒEi�}��>��Ɍ�*��Q��T�'cO���9�ݽJ�����~�������i���9� O���P���̅��L��y!���Ax�ɾ��}�1lQ�-���������4��g?e�4��s,�mź �eĭ���vc�L#�x:��G@�lU"���x�ð��W ��:о�+�~�qK�+O6Aa����hy��VΘ��}3���Rch�8fn��H{u����� ���iC.D�V����R>]�� Z[�H��j�����`��t��$�quB��H♠��q-	��Fl(�ʤ�y�X��!X,��9�0*��E��l����wT�ȊK����DЯY=��6zc�"���jC��=�=Tl�[�.���K�tk�ǿ�
���ѹ�+��rV�kC_jLX]��_����q�~��J�#�TPIH�{����1�M>�� -�+��8gT��~�Ē�V�Uϱ-���8�s�D���V��7�nq��5+�{������������z�v��UV<�H	O3I<�Uɑ�˴l�U�^q\jLЯ����X�WIR���i�5���}�
��D+�k9+�ɴ��!��6uG����
��`{ՙ������6>Y\BI��\�X���	����@=��5�����	��L�ֹ�j��<ORg
*#�L���<sB9�T�Ƽ�����TW+����7m�G�D����Ȭ�ّ�'�V�����3�ݕ��� U�0zeu�.�.�;*#� A US5{�ٞO�u���XY��Դ�����\�N��|�	�C�C5���x� |H��w��@[ ��k���5�mO�3.�lr�r��&[�p��촧�V�x�e��cb���5s�m�}5�1P@^4[�������d�8�� �� m�m_ ���j����N���>�O��:�Q�r�����A��(G9�Q��2\�4�� m��&��o�6�H��|��&�v�l L N��$"�O�i��+���v��p6O�d�6YRpE�E_o�/��t���#��貞�Eo(�jIpa�pY/�*[3 �%����B"[�N1��B�؄��Co�C��"�)��?���6�O�sB�T-�(�� ��~�G�ꚙ��7��;�(�X�(8'6�JHo���ZT��]�'�������5�0`�hwo?Zwі"�^0��6 �:�`Ѓ��6ld���X��7؈w��򟥜� ����??�ؿ��3���?���q�i�r_�۽j���g˛���$�O�>}��t�~���߯l)$U�ړ��/�Kh�P��	;%]=�AsJ����1�� �a;7@���#��+�xǎ`�����($H �P_��y����3K��{��-J��+�b���-IX�ȃ? �M�a����#�Ia͏D�m�o��K~�r��%@��}[�fSK ����`�>����J;	��y�&
�u��&W�G{�+X�0�kU��vG�}�C�#ǧ+�?*=P�����d�{=p?��H� ωX�@�A%��\��S����X�G����.��8'������e�W��$��"�~��B��7����#��R�)%��F$ph�����5�^���)�#�[�W<O$Ţ�C����2.��:��/��4�����d��q�{�C?"4~U�e�ς��������}Fm��$u��aT=��x�S�Z�
)�J^�V�7�i*�ޢP�Ơ�Y�p^&�;�|0t�BPq�j*��y��8.�|Tס���q�\:��wǱ[%]�󉓉%
��۶<��,�@�¶J�K�ھ�ZV���-�(	���;�����:`���ԥ3B�>���=�����y]��F�\�����|=���ꮮ�������jG�&RF��|h�lS�s����+}�#J�H=_��z4�{�A���3e4H&k�=oAj���q�u0������l
��3���b�	��0���J�D�Y�u��m��fKJ�֒�c��!�ڵ]Y3`]�6���[�j���ա,�����kN��q���zK�Gi����G�v60�jl����'-l��^<�;�Nw[�v9j�r���(��� @�r���(P����<�,��iE���7Ą=:���
����he��K��(!���%Ɏ����p��t�h`~n�	�im������b����HB����Ž���mz}y)чU}���37����;aaFb�����$��=MKM�n�(;��?=�m	�έY�b�=|�X���a�����`�t�6��42*2{t�΁�:6�9k. ��OJD_v+ot;�l���6�B@I�Iش;�e�� VR�'@���:�O���/S��n�!&5o��v+0,_�w�<y+}�;�A_�"�3�	������m��4ݷ���y�9��$�����>OL�����v� �ay2����:H��h҆ٚ+� ���	��^�f/�����~����ƻ��J�@/��D�.�bE���8ߩV ��Tp����l���M���S +�G�;��QyUH�N�; M�T�܊�B6o�[ �WP�@���vɼՇ��edc���PIՆH�7EGl���d��ۭZ�"�M�d��Ie�6bɶ�����$�ৢ��[�TU�(��"ӱN� q���k��H:D�E�cN�V��Ol#k�s�C����\������sI�	�h�$�=�:����"	��X�#i��K?LU�R�M�o砳��HM��ᜫ�"����Fb�ZQ%?WP%���"K���4�#��]��݇����OJ�5�FX�9I+��)�y!^��x�뤖�khZ��s2���Uk�b[��5�K͙Q�7����$ŏ�G]㣪**�ѽx$ND�D�ؐ9a��rJ��1�����<C�ؤ痋��与a����� ^
���:��GC�m�L	�q�q�b��T���K"xν�c���R��~pmA�"�d1���$��6��>ۡ�\:S֠XQn�Z7�*��v����˨��)]�/�A.�h2��s��x �>_#0 �pܟ��-h�7,��<3�sb-�Į�}�(H�|�s�y�s����G܊��`��C �g��2�5�R�{)���+�7��bY6��A>�Z��Z�?����C Ɖkd#+�������d�C�|r�X�M�_:���
uepF�S�uK�{`����މ3S���t<�?/�9��H��$syN�mԕv��]�?`�%�e@��=r��o�cU��}�r���(�r G9�Q�r�?�L ��j�5�R���P�#��@D##�Z�襏�yD4�zWxX�,HF�iͩ"p�ލ��k�}��jD�}yyIO��0Abз�7S�4JJn�<�D�G�6�zH;��� K�m԰�8�{hD���
�)�����8b�
���ef4�N\��#�n���5�,�+�r� ���¨A,���1���1r�g��6#�'�}k� %K��N�d��׹�����|y�=Y.�T��Q��^�>����0 oV�`���ˉ$@ߙ*�ꃾ���q�m3p�l�f����g��>C��x����~e_E2R��a���Tд���\�~�8��|y1����{�nu	@��< {+�o$4F�.����_-2R��!�}wɞ�;���s��}��K���W�
���C���]
�slT��Gй�[ޚ>M[?��� �!B�J�e	װ����a��7�0�E�y���"�ʷ��/)�>[I��W����K`Ƕ��H��U{(�$��'P�1^�RԲ�#�B��,�����AmC��T#��Y.�f)�Q����e�0x�>���Tw�����(E������H��ʳT��+�QiI���R�Z���w�ZE��Qy�C�����<��%"<W�D̡몺�fK���^G�MǑ")ZEſEP�T��D���"��2��w�G$�T���u���?쪟~$/�^TC��)��:w����Ύ����|�$jT�%�ҺE6xe��Z���)Sk��l����{K��0\`Ctcݮ����}峼��!0����t��\oJY��q`	"+,�T��l��J��=Am�����Nn��Zs�>ep�Ж9k4\ǧ�3����������"'��T$;�Zu
�������{߳�/=�HQi$#p-�"[�d*������LUW�wmW�q���ȩ(G�C$��⸝����j�/�%G����*�p��[w�����/����v���2�8О���.��{�z������F����[�[��0U��Ĝ�w' kL���a�`sN�r��cp�&e����{�g�'��=� kl�x�-�T�{��(G9�Q��')r���(G�C�4eF�N�mCw��?*���L�nH�o�y�_���BѦnY�?�T����~��Z#)��짰A��t�����6z�^�a{Y��~��)���܈c��d��潀e�5�L�A���e���YZu�O���62����S9����<4@��̻Q=�a�a�,Z���Y~~>q�ˤ���`[�������\r�4��2��e�����e;.���B�y�+?�j�5���r��%6�Y<��8%�I|�A�
��$�� �Zݢ'�
����t��m�\ ͆<�GuP;<�� ,�idD("Z��"HJnR-��>� Ҷc� �m�P?��k��^�4���w#Z�:-����q�ۃ�0�uq�����ݝr���X�>v��ha�|�*�㴼�gn�h�<�n%#������0r��;X�_	'�Z�Yau5VPR��@XޗYO�p����mP��ܨ#�-�[�O²)��+1m���ň�ıVA`K�s�c��(GvQ6j�E��V+��n���v

�� Ej��k@+�/�V�n-"�:�������$�R6�D���w� ���y.�:�l�`��ə����m ��c��\96�>��%:��PR0����Q���2V�5������?�]�pB���y�W�8h�����;�����v�d�I�-�"�{e��NłR�X�]����xU�MsRN�����9㲶s�cq*���#ZL�}���j�������k���iM����P�CT����R�kE0�vdkT�Ȣ*��<?���`'������>�y�tN����;��'���>�pM_�~M_^δK��xK�'��2%�+8�ڶ�9�gvZ|L�@^x��|�.B���3�9t�)H�v��}J�~N����9^�r F����M�3���D�
˞8|����:۫1En�ڒ�.�� 1�~�÷�iN�]=��G�5h�u.��T'�l<@�r�-�3xj�2���e��X+ê*�R�rݧ;-��<A��lI�z'V������Ͽlsȅm�#-ٶ���m|�+C�R�;�s�pj�����^KC�[>>o��h��YZ.|�����|)����*��҉��q�|^��ӅA>��e�ߡ8Św�~��j�*:��o�(G9�Q���)r���(G���+�U ,n��"h1KӆUG ��@�����6��C�Vg�RE�6I6v^�`�{8�h3�x�V&�eM�$� ��k��~�.߿ݮeS�:�)"Ge�@�ц�ϡ,���� k�Q�q~���٢����\�ׯ?q�������� A��!]��ۦ��[k_S�(�p�����]����6�'&ϔ_u,���x��q��¦�[k�r��ׯiڎyp�:�o6ds������b`� +g7������� <
$��%b,O��HCr[l�70���L�jI���_Fƿ|���m=��A?C۬�/���}�����n�*������w�VrPΠn۽>5E|���⑑+�=�[SsX�aXc��>dH����&4�.f�iy�u���g Jd/P-��G �i�=a��rnH�������-*Y�E8G%��wk!�uz���,�6G�Y��H��}El�N1�\������KT��@��h�<�\}��B &l-�Z�~іJ}�7��1�I>���#@����q�6��yTc�H���"��c�-y�=)Q�}Q��g����C�	|W8U:��'b�mQsq�z['����!����E�G�C�IuzTCh,�>�<���o���g ��^G�,��:� �wt"t����񪶅�Om�!��QMU#jw�?ٖi,���؟��uߥ�y�Q��V�sE�#�;���]���tԽ�������n�`|�bA��s�Ķ*ch�R��0L��CJ6�;)�f>w]E����w�,<�@��� ��s`>�o�������?�ǿ���G�+-7���HZX9��t]���J%��k�oU�X@B����<��Oo�y���4��񖞰�������_ :�G�rS\���(���c���y�iw�}pNAP�Z׍8��$���K���O�i��Ef�MP�������W�%���(��"�Q�Y����eLgSM��O$��b�~�u#��j��Z��~��k`�߷�%ڎ�R>���(f�U�8MN�_�;��,�|�����l�l�.��r��.�_�@����+�Nk[���t�=��+�{�
h?-�;��NɔI�������c�(G9�Q��'(r���(G�C���x�f4)b�j4��ب!Z����#���	-36Y���	&��`�����{,��ܢF2���m�� azؠ�xRXԞ�����q�=����6���]�G�Z����J+%�2o���7B�?������w������%�."q���&F�o�븝����88�Χ�7Sf��:E}q��b���q�u���I{�K��_�|ۑ|�hlV/�mj���T�E���d������M�h4��n�F=�G�6�d�U	"5�����qY~���F�w��ۿ� c������[�|�|K_�;�r_�a�+Sc��8��
p������N��H������=��������~�9=�huÉD?�vA� �U�DM?���Ұ�$�~�fQ�}Nn�w��G�¹[	�
�!�:�T��\�G����1 �%q��A���!b�Dv"�����e���+LzB�A"����������A{�h��$�Q��h;%"�9CP�g�;�+�Xcc�aU.X�b��������s:�r�����1z]N��)]�	�"fb�U;�
��b,��"�dW%��H��bj�a˭�P*��Rm�#��V��% W?g�c��T��5/2s%ƺ@ШS�G��_��g�7VG��O��!K�| ������� "(�9�Y��ݑ8�E,�|)�/���JI�H5������K!�I*�7"���7�f��H��5}�6��J�R�HQ~�8>�w�=��ӊ���2b�7"�Օ�wc����u�?QWX%a������e�}�qT,��|H�\��������q�"[5ޏ����/�T���[�' Z��n!t }�ϝ��(�JZ�j\!�<����S��:����<�K�/� ��h��K�{Zr�B�u<�N�z���^��}�f<�4���s��A����\7�����uZ���j�$#���|8����,XGܩ�"A���R-.m=`J�1�(�_dc�1��c����1�eâ��o�d�����c��uS?<��~�����qK걶1r,QUI�տg����/�l6��J$H8ϸ�Wk!�;O8NRկQd ����,*���Aj WK��~@����}l�DҋB� ��׌#�4$VX$ז�?i�v��r,B�"���r��d������่��g2T* �p>���E�4�_{6#����2��6Ys��Q�0F�����_�����3
�J^�3�y�׼�I�;ш�l��| G9�Q��'+r���(G��wG`i�#|N�(�g"hFޭ�LO�l���Vh�F
�����[�NR���yh
	Ҷ�<��cfY���1��"����@������5��rhI�ō�D@@�rF�����"wF�M$s�������`���ۧ-�����6�J(�k���	\�h�lv �Eb*ڮ���j]-O��I��[�v?f�
�=G�8)"����6���]��Pt�ʲ�$�=���	��~2�_��h)oHL���R�v��o�~nF���&Q��=Bz���}�cd�2��m��?��/��IH�T����1eO�ۋ�vX�� ������b��}ü 2������tH��:���7��]ͣ�4����uH�>#��9X��X��̌ �9s�$�x=�bc�l�`47`y*��H�v����(E���h#����Pf�^"���{�O����=�9D���۱ ~ZB�S9��X�����"`�zI�����c\�֖Umb���:W4{;,���cnKuU����'���^_�S�jͮ�����Q��/bD��kO/��0�$�ꧼ&�cD�죢�G��T��jߨ4��ٱ�n)(b�D{U�DF�T$HlW��:�N����=�_�3�4m�� |��r�NT��5>	�Oc�c;Gk�����4r�ɓ7Eu�ы8,�V�)���ڶzMר��F$�����0&��u��H�}��E}8����골�yy��-��X_�m?6o��U�aUw��������)���C���EmW�s��vCU�@�m\`=�B0�5L��믿�v[k\8�Z^5]��@[��h��tM��4].�\�?ʲԗ�������IJ-vk�g��m�3Y<?�l�Y��$7�)(����'��I�3�83��ן�ʺ�WU�j��y`\OY����fw*�A�?�''��0�����$�.�w"���}5F�d�� q]
r$�����D�Y�C���r��f�����w�)E&��T�v� q-�Wu��c�Gm�����y��������g��n���wqogZ�����%��>����b�$t�Rk-���Ts������Џr����V�(G9�Q��O/�����;�ۗ�g��
"ĝ�Q��'6@e�<	��.� 	�	�K�h�b!�	'���v �.����� �qS.�u��(���L�N��� D�0�p۸r����\{n�R2��e�@`jF_�S�˦*�����3_�n�oͷ���N ���ʶB�)�F������l�E`��T�A�$�������Y=ԨlD �;ܬ�At���I����c��ٿ�mW(
g(
�Q@�T��{2#�"'{��L����+�p�����w���-=?����ѕ'�~�=��H�ڑh�����#�^� r�0�x��N^�7g:b"����=�G���'~��������r+�~;~o�l��r�0��@�@��"�9�6����^1o�i܆�!H��h� ��1�܆�� s��կ����qL��ٶ��S�}�{�c>@�Cd�'�YA�!$��_-RW�,r����@+��_ ��3|/T؈$�*�)żBE!���"�1 ���~�8��	��$� �:F꽌��Q��2�[�q��ɏ�lLL���5_����E�K�2������\"׭���6��$洝c�>3��}+[�AȞ,* ����X}�s7����G�����9�+��q̨��o�o�E2�k����"����/(�2��H���+�z�pl<�"�I�H D� `-I�\�+<Kmw��$ɮ�0Ҫ)�l
��k 44�b�U���i� �6gE}�����x��y$�D�H]�v�����JT)ŢkZ����杲+~P���DT�$_h;twB��/��q�wu�C��Rڠ��v'���'���������?��/?����'Wx�`=r����}�܇!��2�������ȏ}��G�K�p%����m��H5��h�j��I�!nG�~�}�w���覒n xo�J�Z?5�+����9#y�DxX"w�V�}0��V��詺 ���<���b��"��b�b�u�VvN>@u�|�XI.��8��Tq�1I� �f�.֋$I|��f�kźf��
��Y��F7�A�ǐ���$iZ����vƽ��EZ��1ԝ��n�2�n�3�����ld������"wت"w\���F��ύ۴��6��#o�j�C����(G9�Q�T� @�r���(��a� ]h��OlZi�(����!ygl��` �B�(A=T��fo:�&ieGЖ�����"nf彜K�;6��\Z�E���X��|�q�����7����ya������9�<�M�8���������������޾�H��_6��H�%�l��f����`o���6���p���RW��ƶS�J� 5�\lg��d^��|c�mZ��w@���"����X�Z!BN�B��%�zm	���O~�����o��/����He�x	��r˔ǭu;�u7�����{����GΓ�d`$'�[_�H�M0vۘ�S�,Ej_𮢌�'HE���P�@�[�pX�_�4�制E-����i\h�e�q��V��YW�<_``������<� C�� ��>
	� H��W�q�?����5�c.�Y%��E-s���CT>A�e�Y9�F���}*���b�;:�H�J�c,�}v���cS����\0�"@\�R��K��9����z�"*d*��r���	���m���(: ΁{+0P6]����4��'���>�Y����EEm-U���������K�N� *s�9� ������5�>�`�����J4�gAN�����x����N*l�i��;�<_jw�@�U)@"�!�BE�W�f��VՎlҤ�Q�c����g�|R>�@��X���V$�ԏ�%מ�y�r��!��\��hn2��gy=�{����������=���q�%k��hv�F�Rb?�u�m���[��=�*�y��KA�;<��E�Z�PP{g���zmk���sP�XN*)nW.�~��,JM�,$� x_����.����ͩHꤐ�K���5b��׶��z��,挘�����S��rOW'�����ў��N��,)Ǔ)q5�c�������x#+V�>zS�B����P\�3g�Ie>��v��`ׅ���\����iM��>�3��zXƂ�YS9.UNP(o��<�΃�g�]n���4������$R� .Z_��P�|��k��AfD�Y���k.ktؔ��6_�ychY�^��چ�K�_:W�,�H���#�(G9�Q��\�(G9�Q���#��,t���m���`1#�Z����������"�D^ؿu��_^����&���"��.���H�
0���8�}�^�Yld����rc}rK�ax6���F��*��};����eL/�/�Ǝ>D��E�sS����F۬��(_�<o�����a�n2��Έ�F��c��Z`�-RT{2Hm\Kk�5���B2���Er�D�+�g���i;������veG���DG����>6���A��χ�v��9� Hs�.�9��7����q��=�i]Ni240�r��E�*�-���k��1�����ך5$�� ��LXh��Ѭm��d��10}|������A�j���ʣ�CĶ�Xł(�����K��+	p��������C4��J� ��fe����w�sQN��B`�
F�D�L��"�;PW@wS׽�Sͽ1`R�|a߆��*�^���nFT��s�T`V���#H���hǣ~���e$���|1�z�v�G�?�����祐3��^���y��k{��cT�5�.o����v%��&.�3��1�����E��Sm~D�0��g�[L^��ed ��)��+��pBA��il'�Џ��uJ��EĎ@m�(�����8�>�:�17�Ȯ�?��H,DRu��
��N�%ڮ}�Q��ֲf��Y m��<A~!܃��PP!��)?I����O�y�y(*gtmq�5I��jͦ�y��ʑ��9D����Qt�Ն;�W����͖�P�.�;���c�{��{)��!ZCU�MMn�"��wb���U�-��8���j�!��a%6{.���>����T2w$�x��4n?�Ę�Ҳ۽����?���,�8�.'ZG�h��^H�����5<w鲭��peB�=:*!xn���9��]G��i��ھք)/��,P>�|F�����g��(}юJ��`��s��ڽ`��*<Ӑ�9<�),u�	���l�1����k�V���lkI�Qԋj#�J�ʒ��cޮk�ۯ~�
\hI�d?_��쥿��$�zS�����p�v.�$�w�vs�T<��b��,c;j��.@jl�#�g[��>Aq�����1�W���
����( �(G9�Q��/U�(G9�Q���<��������%:y�JTcQ{Ц*�H�GEJ|��x��'%2����ܚW�'�TΏ��f&���#��^Ϋ�;��3�E�s�� �l^��ㄼ HV��h�u�Y0�8���4����M������Q�f`��c,|>;h1���{HݓY����mӾ�(IŲAv>����Ah���AE�5���g)�k&�7��	k�T��m�7cNđ8_�(�SG����N�DیT���<*u	��e��ar��ܻ^��׿�5����֦�)�K��15뉑�bwN�I�V���l`[a������ H��:Xެ�x2�����Fdn54��n (S�� �P�mr�5#�F�����������y ;MS"	��&`��9A����;(Nީ��<G��!� ^$��ÁbZ[�H��8Ș�Ca�' /�%�Q��-Ibn������Dx�#�� KC�ҀY�[��p�A.�V�>�����Q$$EF<�]=�+��PkD;����ϻ�����
���|p{)�N/�����Orb�*���~J�sE���ox�6-r$֧�: 8ݩ�b��$����Oۺ"�x�#�"pZv\�կ��![Q�ɠH����#u(}>&/��E;*��mT:����	��$�u���������-�G��^��7Mލo��H�E�0y����G䑮��#�]T)�����f����b�5?��B4�����>H���?o��7ݛHrF5�&���	o�K%��v�6�,������2�⸟o�;�}#'"'^��]v��r�?H��ǵ��.�AI����X�j���ڐ"�c8��X%!l)A��/�G0��M*�a��¼ıjs��4�Y�� ��q�J�#�;��M-�%�uw��R~�>�d������R���#��H.�#�៷�[g��r�A�5`mО�[�

	ʑ�=�z���B�"��ec%�T�>G�m=EV�5�Z�}�u�O�2Ճ� �8���#�{Ɯ�ر5�<�\Ǚ�S�GEBw����y�ډj\���}w�R��Q�r����V�(G9�Q���̔���m��4 �\� �E=��J��S�6W�]�x��2"ODI�&ހ P�qO����k- �[rL��k���_�\��P%L-�4@�~��k�lP��D�#��#��.��Y_��ɓ`����sS�/�����wn�mP���z��F>s3lQ~[[A5��m'���O�G��0i@���[Kn)Ord�&�3�_���Y9
/!���
�<�%�^�a/yTc����?�p�J����!rNt�G�T�
P�3}�n�� C�6`N�!#P��Z�3�wv��1k���=�����fۜ��_��0R�@�Tr��1?����f�ts��b�#�L�v����mP4N�����T	'��ɕ W����h�D��m���� ���}~�����Y;�M="^�#�%F�*	z��^�����ߛ+U�JI�D,��{�1# \��M��������oL�>Mk�<6�}^�~�"0V-W��b�����,m"�X���ʚ+��@s!<��G�&��p�j���:��QE��/V;V@R$�b	}��z-� ��A�}$n����X�H�j�U1���]#�����Гۗ$�����Yd���O�Ve�?��J:������Z�������PY�yF���8��u<�M"Ӣ�� y_əG��M��1ǎ�{*�����j�u��װ~$8�]Ԏ�m�2.*a�O:h���gm_�� �I�]�����_c]c;>��x�B��U�����1���ls�X�?Z�E�ZU��p���hv]�wͺ��ٙ]Q�.�����O�� v����׵3�A���]ܚ��{7X��I����|�m����
�өc���/���|Xnv���oT����]��iǖ�g$s\t��-[S���ף�k9�ŬZ�%_�vn%e�Q���l4%������b9<����B�Z�2(h����sq�3�X�L�Hܮ��:�p���=���=��C��:��)W8g����䋍�����Њ*o���`l��9����o���@�F	���eOl�|}u���Z�a]
"I2!H-���V���;�����e{~�����,T� @b[tmrk���x=�Q�r���k�� 9�Q�r����|��o�Ex�����ۡcT���ɱQYa��0���,(j�nM�����,)��-�Ã����F�u��6V̓���ߨ>A$�YU(W���3�"D"7# �'7�j�-A���/'�{ ��dn�^_^��e`>���wF�Y��lZ���aQy�mCyJ�2R{;��	���۷o�g�"[>D��<?Y�!�*��I}!;l��3��BH}d�!Қ�����vM�i��	���5M�\T��,��!�jd��/E�J�Q��}������Ak�����f��i�{��� ?���,=������ӹ'�5�5۠�d��.�)ػ5�	$2�:���U���U�����rж�¨Q�_�l��:+�\�:>7�2�_�AP�Ĝ"��0�ctG~tV��`����R �j#g� ����� 8����i������Y�~hCt��g?��h��v)�aIT+@��@A���'�.@v�~>F��5X_A!`tO2���bi�������&�\"��J�'���s1�E�c;N����|�$1Q��Y?"@	&�Y�@� �a�~0��~�v�j˹a$�E�j��9W�U~�x����6D:,�����~�Lf��E���w�UN�D��0���m��`;���)b�>�"��=��c)t���5O�������	�i+c��D��?�АR੬�̂�����I]�kq<���dW%K�M�5x��ZH�Z�^1oJ$4#Pw�'*�D�n3)��vl�yZ0�J�y~h��<1(8�P'<�6�_?j�8V�Z$UW�t�qc��$��K�0#�?Y�xl�mM_�$$+��%n)��.��������:��y������IX�T��(����SyFC�K�߄(Hb�)=���cr�s�\����L 	�ٞ��S黰 �Q@�+X{�_@�)�A�{��t\�pe�O��d�Zd�3%�������'"���t��3�l׹�9�y_R�U�ܶ=W���K����� �3��pE�.^Ú�`��]WH�����(Ϗ֨X]��SocuS>:���ϜP�����j�g��ԛ���ž:�4��;�^��k���'����)H@�"��K�/̯���~8H���(G���� 9�Q�r����e�6P��ɍ ����X��l��������������\�V��H����a�ja]`%�@U�$�G�v L>�m�-�o®�@m����l��48����9��6I���lΘ��شb��m�N{Do���7�̪6�G�7�� 9�A���9����k��^س[n��m"O�w���q��� (^	n ᷩ)��H_���Z������}��ƮQ�gE��A�a>e*\4}��	~�N �"���P5#ż�N��'�&�4,�m���]U��4�H�j�A2������Xx��TP޼l�g�&*���P/�/�ry��kz%�;�y����������K�F�[��i��o�ڷ���*��b��Vؚm��S�}�#]�o���7��r���u����ɦ���r������-8��z���5l���#�5l��^sjOO�>���Fw������ǽ�h�޼�o|kJ"US��T! 7�� �#K ��Kȕ�@���y�O��H������a���K͉�| ������<����Dϰk��8OЖl�gH���K��{�u�����Ӌ�m��R�<�T87\�ek���9j��*t:*�F�޶{���X�<]LBu�d�1w��W[�3��%�FO��Y�엗WS� ��Y����t��]u�v��xE�	���'ԕ���˚�����gW�|rNUrn\^�� sK_���uK�$�im���Y��o<@�@�v|�� O8 v��`����{Q4<mmոj��[��z�>��mf�_�W�`?>�q�����5¿�=��8'�|�������ۉ��P�?��d�'�*���73����6�kP�<���B$>3ͣEw����n�c�m�GC�F}J���zy~%(�\F�e���x_}���Sh�L?`���N������7���y �;	�`%��)�-���U@x^Q����1�\$hO^;:���3T[3� �}&�v{�eͅ�kg�3��/'W�Y`�H�vIFc��U�%�\��վZ}�j��ԕ�}�%�Z#�.�'���f�>/��	�ՉZ���x�{c��tn�wn��� �1o�Jn]�bmk_��g�ʭ���\k����>ok��m�rl����6vN��������%����,W_�<<]8~޷~�g�1v�����	B����$�|�Ld`!%qǮ���,�rD�Rɇk�V�&�<��s�2��F�,sQ"��'��H(eM��n�5k���<� 0�s��AhA�Ƕ���O��1��
�P ���E!��j���sl0S�<%����(�/��r' ��Qκ�˙kM��}��Kn%j���>� '�`�+�y��E6���>���<u�5��;�9{�:�k�ٔTc�X�������q^���l\m�B�a��D�V'ޮ�ȍɟ���B��ۘ+�kC�s�B�m���+�~��W�*]g�D�I�XWL��3�}���J��(G9ʟ��Q�r���)���-��������- �ֽ�����\�圼�����U�̮�ȍ[>aS8[r��Z�jn�����6�xo�X�{=�����jHޘ�QRF�U� -L��br#���l��f��(t �f��������_�t�m��8����7��j��E2�u�>W_~~��gc@�(�~L�I���D��&���e�4�u�k��ߊCQ`�l��$>��Y�������Ȋ<Eh��  �F�lN�\�d�������m]���:�,L3 cD���\��n��-��Q�MOuA�, �1�i��<og`,O@����>Ѕuo,��`="����K��E���rh�{�զ;|�G�#Rl0f&�VR�ʥL��|��W�ȲsR�Z�o�����<@Du���ˠe���x{;cǱ$�K�W�&��8U%�vVK"ۢu�~���(���Q�#	Y+��hm��� G��ȦȆ|���S��W)D4(�ꩿq��6��B����b�X RAJ`���ޏ9��|R�D�E��	��vY�(���\/��*
�X=���1�W��,��퐢��(�[���Y ���|�
��Q���b(�:�]��>�*�"(�
E�+�e�_ν�D�n��)�\�`�}9�@�z��s���:X�ye,�W�R��g��Nfy� c��H��uἔ��>�<RL���,kBK.n�	��j=Ws������*�h��{(Eb�t�54{�1$`��H�T�k�v�MA�R�����M����b�["�m4�DՋ�Qy8d�����ؒ�գ�(5U#�뱘�i0*�1=����f[c��Ҷ�qw���g��6g!�u�}��8�p���<��ܫ�IuTɒh'������9&��j-B�v�Pr��|B����!}�r9�p�|�6�)���q&���k$l�zo�s¸�%��m]�qM�x��$)����x�۳l`�8�˖��2�kb)���v����>?�ͥ��P熪	���>--X�Zڠ�j�z�9����5q�UBd�D�� <��K�̹lϻ%X�!i;r��rj����<�bf���>jcjg�u�_%/�_��{S0�}��b��i���(��g�>������մ����r���(��� @�r���(H�cN��r^������q���)6�-#	�J~�?�h�rsō@�z�ai�V2��6I9���wl�-Q: ���Z�A��R�K����X �rI�6fn��X��v��S�ٙ��2����5
ރ� ��ag��&��a����a�� *CD~�,t� ,K�Ip����g��%	���lK\K��Ҥ� L�7&r�����m�O�+��?�0�1`��-��`_�*��4J�Փ���}�?�峝�`�B�04+w����i�[��o￦_����Jy�!AFD?��� 9�<9q��!��m��Obur�`I[��$�D���X��'g�ܧ�j��4�"`է	 �uIoo����s�OP�l�p=?����̶�H��ÞS� oZ@�qAp�"�<�����902܀ؕ�=��f1@�5^��Q��)��E�Ӓ���(��m���g�߿s̛����ڷ-���ɲ����8fU�Y���¸x��\RD�)��>)�]��	<�;��Ϟ���ȣ�Z*�&����2����5��a���~y������~_����8�}ކZWl�D�H��d1��KT�绰��P�㨈XA�Yvy� ��-��õ���!����i3�H��:t�t�����v�Փ�ޢ���5 �\O���[�Ob���t��y��Z�����0�@��=i�Y������k�2�j��{�t��"���lm���<�v{�kPܨ���jg��� r7Lnv��N��� <�0��ڣ?�xfr�eOz�>��ج!g��?����(�cj�8f�=_�k�|����;�+��1'J�Vg�8;��:A�x��X�?���FĽ���;7�@��T�=k���7�u����kS|tny��L����>w�)Ad��B�mlp�8ߨ��}��cc��$��>w��Q�iJ��F��3Ȅ����QD��z�$k��d�q��LQ���d@��7���
{�'� ��(_�QT���"��vukXo+�勭iIP��ԉV��z��(��}�S��2N���.�'_[%*H� ����g������G:� G�ͥX3Q�WK�JF���Kݱ�oE�.\Kq�6���~>o���A"P�h��*(F�������QW(Q����YqM$^�7�0hKء���X��|(y?֏r���(�r G9�Q�r�~A~X�8�۟`�� ��΁@��@ّ�#62 �F���1��c�{�sӅc�4;Hʻ�M\T���h��T���f�&���ـ���ɬ�!��(��O%����f�ju�VڔbË���'�oo�駟~J/���������F����7�/O��t>y�-f{�Ɏ�?[k�Y~���}>6�J@Lh1�em����=�a�B�A|�o�2:y�Op_	��R��|�RL�Zsír��m��G��d@����c�\_Sw~1^�.�۬ue�Z@Nl��m�O�Ϣs��B�%�lՎ� y&�ײ��i��~���rIۑ�}�f5���#}������~k9�g��٘�`q�Sg�?{�v��M^��Hv�?���<5Y�1��+0��S��os!P=/ ]�$�3UPU������8@��ߗ�"*#�9z�	��>�(~O@�����_���2W@e�:�<��Q�c�1�ZY�<=M��T�\ �59P�Zn��zS��Gu���Q�e.uC��
�Ns��	m���bq7��C�_�L�
E�~*�����w"�,5��kR�DU��ȝ���<�F�<�s�N����]}�1��RW�5�c�F�D�f��D�h���ʛ�����H��ޖ:�$љ��/�T
	XE�R��5�OX�&W��ϕ$����w�#�'��xODY��r�qW$}�"UUT�Am����������u�)�%�C�WnD�����@�S�T�Pm�,�{�`Q�4~�^17���ȉ��~l����`sp�w�\��KDv��kJ"�Z�-���a'*:�gk[\q�yB���ܑl�zͮ��0����syk�X������ }�T�7A>��5�̙�?�b=�bi"�������%]��J0t�
����	�k�zhl����H��G�0�%�ݬ\3�,b&
Krޕk�s�[!u���2mSg��|�ց${ ���v�żXM���:�'K�s8�C�D�۞�
�AВ�7
�M�J%�i��L@�ye�_-z�T�s-��Л��`f�a�N�s�u}QU�Z�n>��ܓ���]A@ �p0������ҳo��(G9�Q���*r���(G��
�, �V-N��B ����(A��Eύp�u̲!�=�G(�Gb���h������cY-:4�T͛b�E�|{�����I�f�e��o��F�چy���`��b b���� �Rl�jB	2l����/�����=�/��?q���ͳ�bU0������ۣ 9��3��4� kkI�﷒s�k�>�[�Y�k����U�;ﭯ��p?'5��@u,5Zv�0r��ɀ��a� Η����o�Y,�J��b�u霖�(��A,���- �ȏ����;ee����Q$�ɁM�ke�>��84h�&R�����.O��TsJ�����w�Q4ns�c�x�l��Co�,��&Ex����J���٥�G��$� 2E\���b��ܡ�YY$�pQ���Z*F싼XXfܙO��z�Jv���$ �
�bJ�����1��@�����B�a l��V����Y�YR��U�
E�AT���<p6�%��O�y�_���Tm�<�����(	z��לm|��c����h��G�K�8��� j����
���'�0���_v�&`W�h"�u=�?��=�I�s1uA��	ݣ�k��y1�v$@T����p"R����� �쭮�g�9�z,���-u�����Q";��@���Bz���m��_��Ӊ�Lp�rXվ����>ޟv���@e,zT{Ttq�'SZ&��+�"�<)a0/����]��T���v-�{&��"nu��s�Cׯ11\�e����
�q� ��K�ivcNc=*M�H�Gk*���GT��2k�$����Hj��oϽ�ѐ��5XT�`�Z��aC�������*�hs����d�	I�`뚖�����p��#]\Q���}�>cjѪ�g�40��䙑:Ak��g#��A�4<D��w�����ɴOx.�T�"_Z�����Re���@�t�{�^�0��d=GO\MU�0��b�]E��m/-D�X�͔L�s�YJ&��J"���!<_`�%B���R4Z6x�Y��}��9gSy��� �V���`��&�)Ա� �voa��<���TZv��"��_J���T�28Hu�֏�3��]�im�D��yb�`Fެ��(G9ʟ��Q�r���^~AB�˘��>-�B�K�H��? 0��)��`��o�"�GuG!*��Va�{ߍ?'�拓P�fUd��r/�mc�!y1Og�����bI�;k����D�D��`�ԶVl ���h�ed����"��)C��4�����yVT�'
�-|9���9�9(�u�,�5�2:�A �Y�����큋ߔ6UBK	׺����4z���s��u�r2��m��H�/TZ�������FEC�h���R"k���T���e�=˵B ��ؒ�nL�8-�3�c����b�o��Ą���������ׯ��: �f ��K��TT9H� ���GC�7��6���W����;��>ڳ����[�������F��1�1/p<Z�<��(
[J�k("Yd��y-�D��Z'����l^�� X62�>W��@R�զ"�F���%"F#�	|)*��o Ԓ�%��U���uϢ�"F�G� �����U[�5�+}O�_��T)�EQ}c0�"�	�H��<Q:��N�4 �-���Y���R��ں��[W��'J@m��XWAی����h���$]�3��}~2p��R~�#��l�u}�����|���k�$oQod��af-XԴ�PӘ�����7����>g���G5����nϑ���<Q��� ���9N���7*�J_ʵ���Nk��q��D\�6������=����u~��k'����_0���C���8����(��$2N�g9׸0��Z1bn�wt$�s�' �*�@�#��@�P�bsԦj�մ|�*H���w`)�d&g��*y�p����dI���ժ����จ��d�};/���
vl��J���4�Ҏd����zC��Lu�\��t��"��8X�����3�)�/YpA�q�}���dT6l��rs��u�IǖkU��VsU�r]������cH �J{&O���M��O$[�z�c� �r.�r�j��_�-W��0�a�[˜/#�4f�:Ψ�<۹�p���(G�s�� 9�Q�r����˶:͈����y��i����L%� w����
�]�>'�J���BJ	�=������H!R�����������}WM�������vg��0���%�^</���BN@� ?:S�,n;�z�N���M��֧��#����ǿ��(Z,�&6�����������z{^�&���kvd���g��8ؿ&ۜˎ���zG��r32a6 -;ӂ�j�#y�x�Ry�T�*A��}���q�����\#xQ���_�O?}�~���ۭ���ք��@��j��5�{]&�E���+pA`~`�8;(&�)y�:�`����Zxg��D`�g���RCf=i1B)[�vy��R#`��13q��0k���}���=���+US��N�K��۰�e1���@�_�W`����1N����n66�b��V4!�e�@L��R�Tb6(vN؀�~��ޛ�Ni�d��k��_
�ϫ6T�"�����B�(z�@�["͞c�v,m V�S%fto�y�Ǻ?����D�)چ����??�(�a��{�����VY����$	��׹"Ю�,מ��c�~*u�k������o���˺K��X^��7��j��m�*����"�#j�N1�z�S
P�>Vs���Q{���^{��C����4W���!�#J��{���Έ����ύcX^v'�� 2!�$���Hy�X>o���Q�'��٥2������FL��_�I��4ky��z���{��{���5���0'�"O"?q��cC6Xj�X�7&��^k����C�<;�j��sP��x.�)u��i1%���]�-����$�
A���*J3�D�t�����>�I�O�^����r�^TF�`���{Bs������H,��0��|�3@:�@PH^��������8��1|~Ǻ�	�٤u%W۱M;E�j�uC��,[n4��QW�?g�B��*��W˫�&"����VVz>��K�r�cz#�楬iM�c*L�Q惚���j�W����k=
�����~���A���0uk�'�Ӣ[p�E����K�0#��b[f���CLh?n��f*9?ʺ#5���ƻT�-�k�.�rev��l!��=����k����(G9ʟ��Q�r���+��%M���V��.-��mdq�a�/����\��v;[r�G|nG~��7Eb%�@K�	�q�$�F$XG�{Z��D�Zk:��"~��oaC�$��ڹ�hJ$eYhHP�f�E�����6����$5�7>6��Ѭ��ǂ-��~I��ƨ�y�4�d�EV�9��A��	�1�Z�)�=m�0/i%uN�,��{�]�f��"j�s�.cI,����Q��#��l��Vw���I��9ut�F��8H�}v��kl,��t9T��K3��'\��6 �r$2� 1�|�L��@��ɧ��@�L����j�4m��Ԙ�ɢ,�� ��x�3�����TBHn����+�pչF�?���ZUy����n��iR��- �M�� +�@�X��J��h��#)/�0�(�o��^y�k���'j�Y����I�,vM*"�w$���F�W1�?��=E��h�1�'��nP�p{*����m�b�m�H� Q��J��[��*�u�$���#�x�r�%��=��b���B[��(iv��j�^��x=�׬k�xc?���HLI9��-U��񠺃 ���ʪ&�A���ƬA��]�q)��&�%�;�#]�T���^�!���B�AwW�bjc尡u�t�[��/jw�#��y�d�8v�w�NJ�u�Q�$<S�r�#qַ+�	0)�p=���3|��V�(����q�b�+��ET;i�\ ���"DP?}6��8���h3����e|ϳ��ǜ#RB�и���sͤ�9�1�M��t[���\�d�೷�������?TK���t�u\��c:��ف�Nd�T3=��K�I�`V[����e�":W"1o�[a٘��\]-1�޵e��~������k0�g���y�#LD ���l 'F鯮��z�Y�&$i�>�H�;�=ׅoo�-����-^ɯC�˞S��:ok3�!@"�̋��͟���`�@���n[Xþ�����IuN�~g9U�Le�2�!�s��2g��sX_�6�3E�4���Ї����)ybt��l�����z!�V'��t�>���lv����5��6��Y�Q�r�����A��(G9�Q��e|��Ţ�I�h�W���F��{�/��(�F��6���hZTِ:�B1H��h%��ؘ��yg�-���䉲�
��Zv����)Sr,�Ǩ?	D��[?�t@��������E̵] �V#>d��(�%�e�h֮��[���w�W�'S�	���~` _p�~IO�F���tل��W���"n �|��h��n}����"����>���(7ŧK�B�f_��̚���B6�T��J;-S�8���l!^*��'���|9m?�f$�������'��-���S��IbX�j����|�����F`����Y�lMs�>���;K�g��]�b��:F�C��l6Yfo����~0���.��=?=(���OL(��>~ڽl�h��)Q��Q��t�%������YV>��0��V$� Z���#8���	�RR��i9jf.�"��<q��f��}nA<�X������<���}��=J��b��eݑі�m�$�\��[�Y��-�3�p�w(�"�ډvVLd�]"kk�{od2��SJ�''_GՆ�o$,��@R<B���w"���wT������穌	)e�/�+,����B>Y$Wיּ�	}p�vI����A�C����d��gg;�m�//}���п+�(�R�n7%�Zu��q>(��W�3#xv���s�m���*�B|v��n�_l�q���iʺ��z�y/�]-������� ��y- :/g7xO��r��> n`÷4��XH(�Q����p�Ht�A��T�e]����nlg^�4�q�q�tFD�zj�<�DI�T|�dy�2r�+�5ҘU��g1W�}�+�]�]�[�G�x�yn���q���1�8��$�{'�@dMn'd��*q� ��*��^�c�?=?{>�m}����o�ΆlU� ��`�Ә�|�>=�<&1���?��nW	�V��G����9�.��YH�.'��^�g#�ǌ��y�I�Ӿ;3��<�y��%�@�#"-z��ٞL�mj��v��������Zt8YRs(��m�HƟ�`��H���9Qir�eM���T��J�ٔ���z�,��qw���[���$���V�M�k��v!mA���xPR�����+�5�3k[�p삄8��a:���>;�K��m���	I���5��k��s$Z�aN@���:�}�M֣P�&'��^1Ɛ�������$�:�Mz�����f�yF��֛��1G9�Q�r�?W9f���(G9�^�a���Q[HԌMl��`E�Q|�*F��p�>���o���&M�����R�`��T�"�WD����}�Y���d�'�'+C��}$��;uy�Q��{ȺgU�gC�a��4��΢��|3ۀ^Zy-���r{���� �y(+���lg�jk�q
	�w�d�i"�t�~&y�[�R����
d�>,7���Z���.x]-zHrbd1e�gnj����JP��"	6����Mճ�,U����)I�|����>�\@Ia-�{R�9 l\���oj�]<�57�I
���v�Q����o�EϘN�Sr��?����g�ޮT>Y����V?�¨�"�nF+�e�sՒ,�d]<���#���=٠H��d^__Y/��ѾE�>k��CPI���;�g�5����H~]� N�_ n�= Puǹt]�4����C� ը�����\�QG�qU��T5��������6?��\��{,���bŢ����	 $%�bȀ��7$C,�g��������j�xO�O~d9-�T�b��V�����D�r�@�E�`�{�-Em!�Q���O�f�z��a8����-�b�V?�~f�D 4Kmr*c�}rl7�>�	@�7@]k�f�G�#�5�7��D���7�\��i"Vjty��'b*�>R YA�,��s�+k0fS*�ZDb������J{$Y��^Gy���>I�+]s%��r�Gŝ�]�/��pN߿�1n@9�h́R����b�q�v����k��c��+�8kI�>ur�Ҩ.�c�TBx��b!ځ�*�Ϭd9[X��y��P-Of��*8&Ɋ�^���m\'��7o���s��6P�f7X�>��)(�rQ����v/��;��Z���dc!xĬ�����q�n	����	�Ɨ��k�?�;��s�<��rA�ϼ�l��2���m/W��m��2��ݣ��`���� �3
|}�,�LY
����hZ�r!���ui�V�ŉ��1u
����� ���O����C͂�㳊�쮨M��`��ֱG9�Q�r��r G9�Q�r�?�`����q����F�#�l����7	1ِ�w�9e�&	;>��k�1�,��g���	���$$r�k��-��ކ�q�$⣣u���R�H�!+l�
��k�-b�j
��hѥ�$�G��R�!��=l�-i<6��.<=P�H�6�üO����u�*�Ӈ���d`vY�r��JCj����nJL���ң�
D{�̢)=�6��� K�(˓)A<)��I��y�1���=k���~�����|)`�E\.�r�ص!��" uO�x+7��ǉ�����m��ڦ���v �� X�������0���*"��f��z2	���l�;']�:�?�{>����P5�s��+8 xe$h��/��ґ�<g�0A���/�p�*����1ҭ�ɰ$д��v�n)�
��^\ͺ�,�:��f��y2xؖ�� �
�����9D
�t�~�{ %�8�{�a��1o>�]Q3PQ������w�UO�S8�(�Q?�l�a�{��6�m�jL퀱�1*�u�y��3j�Z�4�#|0���+���Z*���EǉJ�x�*� �
"��}�=W��?��{"�d#u��i$]�����ҏ�w�q��\T�4M��M�1��.+.�J��Ð�&��[�XW�N�)�J�f�@��Q���d}CWUi���Пٴ!j=YN"\�V�e�\O���������%��]�@ ���m��ۑ-�/z{>�R��$aNEU&�?��V!�gL��M$b��6����k���s&Z[I�$E����\�;�7���}OD��A���{�\?���� �9/n�/���hÉ}��\�?��'��:�If�y�#�o�+����J%֎ʠ�rY��]���Sl��Gp�Ӛ}��}�CS���Z�M��<} �/N �b��E�!x&k�bV��=s�4���?�v���L@M�7��D�K�KF>pA+�O��R�J��������c[�|�����ɴ,�Y�[}A�ޞ�i-�iZ���R�u�n��y���2T�ZD��ȋ��SYcX��ޓ�3/{l�a��d�h��Z'�]V����g��B��v�8i����d=�^��̕� ��4^��omz����:�*���g�>���yf_?,��r����\�(G9�Q��	I��n'�F�[4/"� �Z�rOX�@n� uwY=�ٯ��&&=w�`�D�i���m_eQ�� �IJ>.�
�jy���/6������Xv�Ŀ%_�X�N�Μܵ����cfI`�3�o��kʣ����c��5
1&��{�q;.���v!�|遅�L�è�J��g���,Z2�G��VE%S��h���S�m���>!1��KݥO��%M�qG������͇�������^���yo� g����d��_,�
(�9T<r�&��r6�5�(8�A����.b ��g�����I�`�=�@0;W�q�g����"� �@��q�׿�bG��`>J��T�ĨƐ�dr� %��2*��V+��u�h�"5~t]
����H� �x�Ő"���K�����\�X͗j�)퉇z=�V�����<����1R]m��Gj��_	���=�!�AD�K��^�s��w�/���m�D�	�4�u,������ȄG��Ӫi�;�;��H|�5�m��P�1�y�?;Q���>S� W����bk��e���3��6�cE������꫚�*�٘�#Yn��ݜ9_v��X�ȁ�7KmڒG��u%H�E����5�DWUU�T-�4�E�H}��ƶ쭢u��2񞊬��>���#I�kS�E��:u=� @2p^�&Q�7.#�m�|2��l�p��G%����s5�>u�'��c����[���sd�5� �G7����:~��zKs��٬�ln@�>����D��y���6'\��>�"�����@n�a�O���o_��X7!I�ǣgwG�'���2���{��a�c;��l-��n�<vx���jA(%��֟��9��z"��9a{�ߊu����h����q��g8���k�sw2���~�֊��@ k/���|o���"�/�-�6�[[b~�c�r��O���d9Rr�[�u�W��Ͻ����n�;�2st�'ؗ��������?�Q�r����� 9�Q�r���!�]�A��H���M�R�xO�T7�}�;�w���6VLN�������s�7Nd��:E����iFxޚ��� ڄb3��|��LBA���U��:�|��oR���}������\U���n&�����ޛ,�vdWb~�t���= d&���b�{Qf4�Ei@3M5�OhV�Q3���%�Hf2�FHV��4��dd��Lx�6q#�t^�����#�KZ�*q<���i�;�k��6�#�,�X��:�Vt2k�"��r���iR&ˬ ��JH@JL"��w����Q�r���5��hᆼq4g]B���y���0H$���~x�28�< L��!���0'�t!:�1/%f~^D6����s�
Y��E#,g�MYh���
�Z�L�MT����d6Sfj�/	ǃ�b�k"�Vߙ�!�"��S}bD/�#�8+ؗ�Z��2�V�0!�0������O�<,�?磀���#:����������\��Y~?I� ��b`�Il9 }wIue^��'Y�2�^H���̽�-*3LN'i�+�i'��y�}�"�QB�Q�}J��{�o�q//'��l�5�kǰ:����]
�x�0��:���7��W�t^t��R)H��5��.%��2�-fH�Z��\gw\G��c�seI�lԃ�H(����;I��
���`2f�?�`2�2�we�2p��y0�0IͅLH� �}�wX�P��BN_J Y��u�?� Y&J�;+9�e:�F�H��{�C"!�]ԙd'�l$��j%0ɾg}s�j)	2<�[D�#�|�~/��x6Σ��X���B�������bI�u��h�5��V	�m@���-J"ƞ�%ag�4ґ�z��/�|�����m�(�����c�X��6�K��Df��c��[��hߴ�\J0Y{�`���dq�WDo&��O�^:OVC��D�:N7
0�ϖyv�//��Y����O�D���y���!�:�/�.�V����a9i��鿅����O� Rd�o)�|��ssSo�~4_$WI�-�>������'�5Ϻ%͂�r�<��
�C�\)���I`		�x=��:����q��f���he���Q��.�Ap	IH�VY��$d!�JY�~�5�0�)PF>[�3�{��o���"^%G��܉�*���y��O��=�|���,6��9iT�;p�*��`dc��1�!!�D�+�j�^7�~k�<�~O����r��4�g~�2 kY�Z��],+����e-k�V�Q$\�)��`������p8�H�n'h#7��D6�*	@ҵz��z�G�Œ���5�^[�E(�lDůB��H+��*MT*Gas&��e��=�Y���/�V��(罼f�F����'�/U)�%��K(QF��w�I��3I�  wMS�I"	���-�Y�5�m�hF�����_�m�G5��%�`w�y�iV��m�yb�C��?u�i�oNjY����?\��п{�����L�u>-�{~~t�����N�P K�wK� �)C���<�g=�4�*�*pN9���� �=�D�M�I�-%0����#� z�<jT��np��	��w��l	��zӉ��$Ć l���9s�����>Y��Z��@�2��@�2ڿ�R��~�o00Ѿo}܎)�a���@�/3)/��4>!��_hJת��[��"�^U��P�~�ZM:	��(�?!�e��ܓE�[�[1��N�k_e������B���U)-S�I���l�w��r慵C)uM
ȸ�`�u��Ǵ{M����"��mg�`�X�3�#$�)�ڗd]y>�s%�_f�����=�%Y��T£�Oe�6���o0T�-����%���@s�`��|̋�$��>c}�u�5	�7���K�3.y���҇�'i��>ĶYD��<��P���&L�3���X���V�y����a�s�AZ0d���(�!g��l7�Mr�L#'���mN2Al�c����-��־���'�d���iީ��~��2���b#٥}�s�(3x��e��X��k�gk
� +�%!#z֙�.}?��[YR�¥�G���"DW���g�s_'�\\����;�8h�%��v��$�vC�<���)j֟'`/�r�rK�]q�1M��̫ThA�/�o1Tr>���yX$�H��N�f��a�+�]��鳧�xa�9����.�
���y�Xg�L&���\� ���1��q=L�T֗L�@X_���4�U��e��4p������'GY�����0u���5�DR��L����f0�Z������L��z�����C��@�6���#@
���du�77�J~�e-kY�w���Zֲ����[)ľpi�25��ĝl� V08�n��⥀����𳛾s-68�Ԙ��0��Q�a�b�U9Kd�Sܸ���/�o)K��2��Ltd`�I�&B��b�D�^�#.m�/^&���ͤ���86���(�����Ȧ�4p60*n:/�8ۈ��'�D�1�5��-�J�8���b��EdmX�'���z�lx�id�T(e7�ˤ��PF���aťF���Fx��� 2�����?��ؘ7�֥�������y�w���kw�3���%�X��&��&Xd�]\ֱG�#����@]���B1�2�ܫ!sO��R�	�ڌ�zW�3���R�d&�9e���$d^r�-@��� �v�,Y���3"ü2ʈd#,S������2�@� J\�L�G�^�W*g�3 P R���#�5"��7�	R�Լ��K����bJ�^ �h{����k���Xf���*�r h������c1%`j@�����7v)�n/�m���
�Q<S�*-���;���,����Q�e)�o�4�Ǣ���`����9��f�k)����[T= �:ĺ~z~$��v��i/�/J��-sȸ��z���(�:�?�y���Q�.������L�L�H���]f9y?��\���{zz����d��$���J�s����ֹ�xJ��������w��"c��K/�Z2T����珟틾g�b�Y��6:w�j�� ;�]�Vs�2Y���ցTQ�I�8s%	)�1�<}�]�DM�+���1���b�hVoV�UV��v�6ϖ�-=K��+�B&�Czۿ"%K�Xʢ$��.ǩ��V�'f��8�\f�F�3p!gvH��He9����ȲYY2����C�pq�]G�	�� �PJ\`�����������=����r��f�s������%\�I(�	!��e!�Xhl���;ˊ��I<E��y�$�k�l�̛Ր����*�H	8Ь�щD�����,5U�8>d�|q���1�>1��G��<8����0�f}����a�r����a}��O��g���\��ǅD��l9z�a��ܘ&��Ui��̫��=ɬ�Y�3�A�FdWwNH� v]�ˮe-kY�Z~��J��e-kY�Z���͗�Js�IlT� x���`���~�wwqS3����i�]pF&��7�qC�P.K@�Y�T����ĉ� �1�T���2�`�G���"�U�@0>�.:7�,G*@����e!$#�� &?PR6B�d�[z B�︱~��AQQ��+7 �Z�T�Ѩ=�ęU� ��/ 9��̹�4�N6��}1��Al�QI�ɲ9��+~�!|��@
�B`|�-�&�ZYY�,�����1��ab�1�^����H�U��e�I�����T/�X"xz�}q}l��)�S�s�%�~��B?�w�$Y<�̘���O���v<"�a(�I����ߡ��\��b�/ ����,A2O���o�Z �KON���4�c}N	�-���R r66,�]>�	�$�%d�����
V��q�`=~p8�&���H�|��8�Z(��10���J�X�� �3��p���ȿE�膺������JП�AƥɄI:� s�fS_eYT��uS�ĩ�w	�[[�y���w	�^g�� �u[^#K���c��]J�u��/���qoFp�>1�V���@"� .2��s;^h\���>,�oHr�$`	��m�n�h}����؍d���u� �����K�#Q����5�^�3��y44FĔ�Q�	��:�=�L�^!�u����gLYN]�d�o��ڛ���/ڔ�`z�0|	i>����S�d���ss�/�䗃����D< Db���y���q�s'Z}&�
2�U��׿K�Ԟ��cF�adFY��o��$�ݣ}�R]��PJzY2�&!E$��y�=/Ҏ�1�!$����1�u�W�0�)\�4K7r�2E�/gJ[�D�yP�rK��\>3��I?ts�-^��=�[��Z]�@��u*eFF
��iα�0Pk ���oB�����w��a�Z	I���:rQ��s[���X�z>3��ߴ"��@�ys�z�la	"�򘓬�}]ѷ�2N�ޗ���qM�!��d=L��a�s���� ��yJ�n�a$�u=���)~�.c�H��I�"�2���kǥUzo�N��Ifx���F=|�ᙄ�UQ��Ǘ�ZGIVJo!h&H���	1d6b��L��c'�s̜�x���tN�c\�|��;n-kY�Z���)+����e-k�֊d\ �q��x~9�u
>4L՟�B����n����i������Ě4��*�5�ㆳ��i)��	Bd.�w܀�
�Z$bUR2�ˁ࿚��X6����XŻ=�rl�F:f� ��fyV��i��Y�l���h�F5��Y�|�5���i�%����\���nUBǢ�A!��UC��m|������4��F�'h����&�PUx ���#������f�f�M��Nt�Ѵ�Cڐ3ݎ�J��(9CN��w�Xxj�K��Ly/G�:3V��!Y~ù:K���ZN#AH��g�5��!S��w.���S����J0�bP���{P]��z K�/�w�� H@�@�an�:<=�=�A�
��2ۧ�X�8L};��@" t=N��(b (���#^�{��#7�Tdt���W��4�����������(zdM+��n�~s�"�����Nߺj*dlt�q*�g�(8��f�"�pE{�ǌ��c�sC��o�A��E^kLQ� f�zIm�]�XX^�;��A!� �QI��q��i�b�z"���U��5�b�'���ґIr{{��I�L#kF�vm����q��s��J�4����/�J�c���Ec?�ܓ�=�C����಍7�y���  ��T���i���E���<�׎f9��Y&!g��:�A�\�2�hգ�E7g��V��0Y��`V�=t�H�6�}B�
s�sH��N�MBJ$�lM�z.#���RF -�x5M�� ���T�c�	>�q�4"euww#mρ��������l&�xdF����)��_�8��V!c�)���&�gx�ƺĳd� ��:3QTF���$��~��qIb�]��`<�������� �#sq֌3}|�C*���ee��	�1�g���" ������x���!�QH���Y�{�.�9�gH2i)�i�߁�'����'JCt���ĥ�="����B-A�e��#忴/!��0$�t�������"��b{�9���ߔS� �v��9w�]���r� ��YlD��3*�`ZV��ێ��q=4'B�����s.��RD���w��17��N �����$D�sJ%k�G{���S��x����� õa���s�N2ũ#�w��g�P_�Pd���1�A|װ:����xm���:�Ɛ�R�H�#!	-����D�t�t^��C�-;���I��y:q-rG�Wj��ް�l*�C��!T�E�B�p�d��[H^�~F��>���x�c�ߖR���8_����	y)�5��� �m�púw���w[��ẙ���DS��c��������q��g�	��+�D��������������{����z�,��L��r����3�o�7n-kY�Z���(+����e-k�����S�d1�����$&�v��P	����'�Q�+9�R��	�r)I��3f'$��ԯ�"IQ�0�R�ߊy�-����3ct!Fn^%
W#>��戻D$�Һ���T�,n�dW4��j�=]D96�B�4M6�<�Fա.2, !�h#bT�S$66�����|�:��ރf�$Ӻ���%!�MɅI�rHjBN�E}��|<2��
��ڧV@� O�����ͼ��D���s��%@x��s��-��!6td��<@
��tv���0K	Ѱ# ����H�M�C;/�@º@��T%�`�v�H�	-��10Z����fB|n:���	7b�&{��R�S�5����-��Q	�]�2]߸����lU߸���m*�FNk��z(4=w
p���%flnmUF�[��ɬXtsyl�#0�����{ �����(�d4���dW��M%(�1P:��t�&v�:�t�Z2L �ܭ�D��\��w�I���S�V�^%M������B1�@n�	�NՅ|�e� ]fx��%��~	�܇�M�����Jvӥ�x�Q��f�z/N��ʾ��U �h�7�gfXHF"�1�0��Q펀�׬,J���a׶��P�	���r0��>��ӜͫM���*��}?�R�u��o�"�_�$ƕ��eFK_dK�}��2eIc��o8�}a$!���ۻ�'w��e�����S�_ ���D�4����0ǕY&ii� o��If�1(����r?4i�҇�~D�T�,%gmk�Y�I�w:��t��S���{�y�������8-���Q���y~ y)�����V3Dj�ȇ&��]�ǽ��4K_�yMHZyF0*�B�2��Է�!�L۠NZfX8����]�_u�wI8;�h��ep�Ԑ��:�p]��!�Y歁R�S|��e�m&�t�<�|�<�8˾I#�9��\t�Z�nʬkH>�̪�9NS����C27ln��.�&�<����]m��&�R4��s�s�Kc����}�.砰�����i\HƯx����B�0��{�s���Q����,�/�]tM�:�'���3�ٲ.�A4��F�r���1���^c���1Ҵbrxz"�y�x������a�k���QJp�$�v�
�&]*��k-kY�Z��K]Vd-kY�Z��^z�P��(S�P��fg��,Щ������=��T�H`�Qv�
���rI��w�jҽ�I:����/�b��g��b�z��3�
����@r5�n|�-%s�qTSߙ���T�!�"��Fa��+3Z�yz�hC�_�Q�&P2V���cjr�F���Fd�#�^�B(1�>��	d�/"B�r��F�g�(�P�4��(�R�F�)e��5h�Ω�;����1ėb2Ny�|�q.��Rk�=�i�ؑ����ǦZ����$�����9�_(1"��Y�]�J�z���5�O����8���]U@��؟�Zd ,�W��4b�#��{F(#���8�AśA$1�
�B��\$?�2���t!�/ ��	8m;������;w:���R��/S��%��̵��'��@F�My�F��@���F��}dJ�Ԣ��oc�DT��βMv~�-$4��J|�X]]E{������P����5(ˡ6Hf��IX7�-ڮ ��$o�cI�@�ۺ �+� ��W��`�.Q��N	���-c2Kl]��%0�A�\�e)���w��ӿ�#}b�K�<��4(.�_�5���d~�}ʽ0C|��$]����S~�����x9�j��/ h�ߤ��33(�_x�F4��g��#�Rq�!+%���P*�� ���x����_�D)a�)3J��*	��;F�I�ʆ�{!�k��܌�/d��^N!����0�s�	&ȒT�d��.��-�a�i��g��'9��|v�l|d�.d���ik�	/�zfPn�"~�k���� )�8�0��z3qö[r�g�	����K��p�Q�����q�&�{!ܓׂ�VSZw�搌(�n��RN3=�H��3E�����5� k�9>��.�~�d���q�f�u�t1��$����i�)Ķ�<��= ۥU�,Α��cA"'*�m<.
�K���>�=��峬X�$¯��Y�Z��@!��J��L��<�V��&7�쀴� -�k�33UDʴe�4���}�ė��T�5�����:?!;��}ŏ�<x���kȁa�@�	���Oُ�7�A���ڀA��ߘs*Yâq��1���c6�҈�Z��p���ٝ�I�P���vCS�4N��@�x.�:z��F���:E �G�a�W�����
ҽ.`kY�Zֲ�_� kY�Zֲ�o��ӏ�8O7�]+@=��/��b3O��yǗg�	�hKݸ��{�XW�2��2,������{���Y�a��?��� �T��'����R�D�ٮi�`�����Yr��k%�{�\Da�"��sU��nxRUf<h�\?x;̄]�_3��r*s�-�:\��6�j�V�" �eV�;�ѬK�S6Aɭ�j#��XGTQ����c]{z��\"C�u������_h~�w/֗ �ن�<K6������<�DX����3S"� z!�q�iy�~?����+e�������D�;$^�[�~�E�(`�e������Ӂ<S������M�u����Y���H���B�R-]��������zu�h��Bev���%Xh�k�\FA�Y!(����cGܳfd�i�gߐ�5Rf��y��뺈2G�(��K�]$K6�b���h�����1�I"��e��ub��l�@z�8~��0%`�$/�������G(m�F�t_G0���N��D��s�np�����M��o�g� y�̗�
�����k^�3��׹��p��rj���g�D9�V�=y��,5�e���,�2�������Ӟe)�O�&3fY�T�'��OZV		}��f�Uq�6v�,S( Y]�	��2�.;�]�dk�[g)�b��dI����^Ȥ�ƺ:0���<��?G���e�XV���������$9p�����eɔ���>˿q.x)�$X9�m|��.�)g��.��O���랪D�`B$=�-�<c�ݔ�� �lo�o�5�{��k����u�ʵ6�Nk�B�"�$?���Ks,H5⡴`�7�c�~<A���,Zo�Ph��J�� c	��Y�w�H�,�����^Xѳ�X�H��e�-��� �^_~��`�|N��#��<�[���$�f���uI|r���z(���C�nй�BhF1?� �T��(��%ҮB��3c��g�����:O��@v\�l7��oa�z���6�����l���\��p�J3V:��o�{��n�>Y�d�A������0T?���Yג)�x)��l�x_��͝c}Tq��麪u���G�?�M��έe-kY�Z�3e%@ֲ���e-��[�~�y���T�7�s7�fx�Mm���!�B2PvA�z����:�#�ʛ�p9�a�
jH	� ~���8)!�bt�L�Q���9糂Ól�)�P%:A~�ˤw�D[��iک .3@2pl�Kp�d�y%6��fR(тϢ]�#2ْ3=��fʩ�T]֝m�+W&���ڂ'p��Ne� �"����f����������~މ9zQM
�
�א�)?|�>R�k�TG����Q����>q3��7V��$:"}��*Su&�u��6��P[�����"D�T�!Ԍ���x�M�	nA��E�����!� luM]��믿v��|/�M���u���q�f�l&/�%Ж��xO�������3��!���<ȹ�oQ�%h�@�*$y������I23 �eཥV�ר�R[����w��1))#7,"_�����(z10G{6��[���2��$�t��h����\�D\+	�6K��l&�8�<g¦�V�!��!���Z&.��D��������)3 윗��|X�{v�e�w�:�"c�]/���EL�kF1����9�������:���m�)l��<�dڙ�e��<�
����J�ﭿj��2	���R�B%�m�$����}��e%i��y��aGy�EX�Ԗe?1�ҲHG�e��2���q��h܎�5�(� �1}#m�v���oQ_W����>�/����H�Uu"VD��RNo��M��d��4R�}R�t�[_��혥|��e"��%������ѽ;�bu_� 6o��tI�&ˮ�>�Ae��>;�,�X��k���W��!�� �E�+���O�ynHD�oGf*b�A����,��Ԕe,7�H�N̢�Ԧ���G�}�g
���ߋ#!/RX"O9��X�Ǳ��*z�tl��pf61�8ߵ$���ĨH�ԉtM,2rݻ��V/��%yɒv���y�3�9;ϛ�wP��F *U����>X���x�_3٫�V'�r�}K��F��l����=�#Y� /�?)3y�,�՜���S�J�.���9�F֌3��Nh�s�i��ͽ�{������W[�'8�t������[���2���r��Y�x�W5��hb��*��Bu�_�W�����?��[�Zֲ���җ� Y�Zֲ������ >����.��H	�N��i���6��Lky	yc��D�K,�Wj������&�E��%���H�ޗ�#ADf�N��	��B����W�:Ȁ�b7��.��I�dGQ��I�x��ǉ�r��F��)�`�������,#�=����U���J}��ղ$X�f�Q�*�U9�� ��f�t���H" Q�A��v��$Qp���&�w(�����LjԦk���%��q;���B��mS!	p��|�U�����ah=�à4Ⱥ�K1N����;>>���q��R Bp�"���U�q����r S���� I�I�tY�{�m���{��o޺/?���|� 8"���w�x��m!{���v�6��=	%��@P�@����`ޫW���K�����I�X�y��B� �i����)M�A"���g@�IO��nMy�9�C�ʳF��ԗM����*;b:�Y6J���"Y�O
:���F�i1_��F����}��<��{s��^v��8�o�v��n�CȊa�e��@�����e�F	��o��஁���J��}?D�����6�܏��I4	�`�A*�s��iv�e��]������~�j��*�dn���B��A��W��u��u4~�FB����/I������׍���e�`�W��x��b1��c�����2;�28�{)A�2���m$Cy����y�s�L�]�k��QF�it:ɹ@�^^���9�$9:�>�k3�.fIhv�e|�ic�f>E�E��0*I�D�5b�~Mp��i�]�{{���ƻ���e&Y�X�,���K3�9σ�����`[��?�ܦ��[1��� }O�V�t촍��;�J�C�]����l<��ʮ>c��L�V�y)eD"׷�|�~�)8�d���M�̊Y��,%ed�(�}�^6�k�&���bulc�;�����́$��%֪XK�ܾ5YT�r0�4[vb��6wіi^p!y|�eIsH3�̙:-zq"?5�Ndb���` �y�{h6����~�,�X�3��Y˺I�$��5�Yw�ږ@���k%���7NB��̈́�'��9�о"��v���	�kµ�5e��Z��>Wg����F]�O�:w�)���O�c'��*~���f��	ӭ[�Zֲ��|'�J��e-kY�Z���{����Ɨ�9�G�"��q���H�N��%n�F��b�)$�� ɍ����ɖ���!���/.
�)!�\mJ�g<�]3�Rd�D�_���Sд�駁 zFe�M��M-ѱ��Y$�j54�Fډ��wB�,�}��۶�2��42����O/S�N_�N��#K�F/�X��Z�_�0ˡ��!���(�YKu�D������c<�����i���H��'�%�7��A"�Ɏ� ���t�x�v�%�|��Z3Kj!Bf� G۞{t7#�7�z�ƾe4z��v�l����j�mr�z���nŗb�*�d 8�9�j4�|A�7��m�7��)��s�k##:����Z`v���AV�c<�W_��}���>G�At��-'���n�f���W��)�.��A�2�'JM��:؀H�ّ�1P�x���P��i�L��R'��^�D��Mt��Ä��sa��L 3�oc;O���){xT�dC�؍���h���E��M��4�s���7䅁���N�����]F��?����DL۳���v��zI��I&"�J��B!s��S �R�Q��Lnfy!;�e��=����Z��R�%Xm�`
�=/�6YfgV�rm�]$#����e�2@�D ' މ���O��&�TqF(�ԍ��.&�����  �b~���{7B��LM^fa\g�\�y��s�R���3e;��e�o�Tf�ٽعD�r�f����%����2�R#���*�̔Af�I�.!ɩ�XFN�\x�̗�Jj�"MH�KY���,3qʬ����|_y�6��=k���:`���v�%�R�Řm.�L���o���c�c�[�q�2���ˣ-!�D�E#�ջj�� �x��Ie�\��܊�<����7D�o������>���3mY����V@�������n����?�/PWM������{z�q�"�st�R���,�D�^�ߩH�?E6�kN	�l�_� �������˳qN��X��[�$l3�V'�0C�M��n�);cۈwʲ�uQ|��NI��D�a����v���_q= �]�̚���&q�q1l㖙�.y�,�X+�l����"�[ S�zO�Z������ho���l�>�;X��x���\ȧ�����U�ۂ�N��{�ȝ�.X����ml�����'������7n-kY�Z��(+����e-k���N#Ӱ�:S�y�f��}�׍���y�5���`���L ��m���Z�F�ldPH�_h}��{����X�f L<!H,T j�&�L4��w{W�#.yV�N�$s2�{F�UU�6n��M+�%���rb:����+ T��c���1i0#�fݠ�%��F~�Y"��]�ԗ���N �m��/�.�>J/,Ne,ml�G�hq��c7AH` ��fjw�T@�M�<�f� h������J�D�B����n]��X/-��d`0������.�'���4��:����Q�4�5���	2A� $����Hdl����^��ȇ��ӣD�&�mJD ��x������۷oE��`A�N����[���N��B샀˒��	�Q��?'������*9��B
��@��

�o���\�t�����H�VG!�`�k+���I�'��S�v��KI�i��;�ѡE���m�a�_h���J�����u 4��&����E�g��_����9��6w���1��H��7 n.<>�A���E�K��J	��rJi̻,�D�5'Rh�G�"�[)�K�zuX��7A]	��g�f�i�3�0w �m���ǢS�9*�� OAFH����
�����[;^��_�GY��\�H�w�̜�ޭ��8	/�A��VP�k��EUD�["���U!q����:���w�Ҽۀ��M�R���e�s��"d�����6ޘq�s���'gI8�'�y�lPq�x��Yb�/ǡ��0�@2�(6������v(I�k��;��8,	�2����8༦�.�v1SlH0�����
5/gV��_;8���c|�l��Y�.����qS�yx<�c�5�
A���<;Ͱ��܏}�W%<�,�׉ױ��xƉ�kT-d��N�x����� N��?��D��5�o�M�,�"d�H���D���,�#�Y�c=��˴M��5��ȏ� F��T�SJ��,(k[%��ܟ5ӱ��j��Ō�XC\A�s���Y�=�l���;�|m�m��uw��>"9���-I�@�0�ü��uð�\ �k�e]�u!�Q�JD�a@�����Ձk���)+1p�mv$���R�H+��c����^�G�H���J���y	=�Fd�H�����	������Ė�ǹ����2��O�Ź�տ�W��?������K����e-k��.+����e-k�V�Ll
�Ycww<2#z�5'n��	���DM�%E5vqS4�5u�F�������q3�F!�X{���1s#F�.�!+���	*��b3�S`�DG��a���Нir��D�\dp��ۻx�g^
F{�����[��I<!ɍq���A%6�&�dQ��)��p=��y�3A)���~�=t�_G�A�"�@qO � 	d= ��m|�R���Z9���W�mH���͒���3|`fJ�ύ�d�xz�@��6n��!� J����6�����������Ne6f׃Y$NyQR��}W�@� 52@�H� ����!X �r�<� ^o����\����Wn{��|���U�F�}��>���S�9(��}��{`��F�� $h�J����_~�9A{�
�W�&�̸�����Zl���{||��{�HD/��}�Og e�В� ����l�x�� =�� �5:sO$\�h`d~�Op+(�f�� )�L�x����u��ܢ`�JR�x����v}��/�i(�w!Å>����k�'�b����|� x��c�c%@:Z���s�k��qb��>�8�l,|�ȑ?���>k$�׀���iP>�D~��%y�4�������^K��qX��[��v����F��)�au]�%����	U��O�,�v�`���_\/%��78���Ha/@�4���B���+D��6*˦$�ϲ��Fpc�ë}#�*"��H
���[#�Gm7k��̏2��2l��2���K�܈�d*%�ʬ!����,3�$�0n��#oLfɀ{�f`���P��e(���=pc�j�\Z��B�:�1�������;���K$#�>�)m��l����tZ%Yh#ܵ�)��ٸ3i�>������~~&kF���1��YE�hd��$x��.C#R��}��: {F��ϜM����&�~N}�3So/HU�����5R��1>�&ɬy��.HS�����#�u�`y��u��ox-&�%�t9>��V�U��*ͼ���&��1o��<dVVZ�� [��I�*��h�Ww�`��=�#���1 6�{��/�;�:xq�n�������$H�˥���W8'��tC����^$�jΛ5�%Frɜ-b��d�ԕ4�>s�D1�c�I�ǚ4�v��SM��|�Ye:��3.$�Fs��T���E�T�IZP����"{�'~e��P���Jɞ=�g���Ȥ��<|�fx�`��O�B���.������ ����kfE� ���l6���Z�J]7��xf]S��<H���O�~��tR?��������{�a���v�ɮ#�UO��q}�י�N����{>��}\h�{�;����x蘮e-kY�Z~��J��e-kY�Z�Qd'lV�$Q��W�_�$��t<Y�<	lָm� YHB��("�QHk #2@h�2�a�z��y~�$� �"sbQ"�We�ﵥ�ʎB pH����K �ѫ>� XMʰ Q�|T�e%���\ �x����I�мVM���s>g3K�AC�|��cXj�,[�S�+���E"N%2�|?L�_dj*��J|�
"t� �D�R��r-��j �MCI���i?M�������Oܗ?�Y����'zs, *dk�D�#n��M�4����}�0�?���F��W���Cmi�p4�}�Ğ5��k���u�wwn (r���^؞ �Qu�US��-��0���˒@mO�'�S���K�H���"�1Yǿ	V-��*vR�93��d�P.eNT)_�I����4(�%@���y� q��h�6��"��I�,%JY�23���0�rd]����f�l�F�v<�[�г��E����g� �5/���c�n�?�P�Ho��)����w�2\%m?�cuYF�/�]�+e$�5 �JDLIj��{	ؗ�[eVG�Q���<�k�*��<�}�"BP=wxy����,��˓a�N�o�f���������N�ޘ�6��<Vr��KmZ�עD�]��C�����)�_�M�wK��:�$6��e&�u;��d��>��Y��:C*I,�cev��⸋�u[c�r]3��u�/��Fp,���]����1�YY�6ϔ�fb9�X��w���J�����e@�}ƈ�2��~��.���˨q]����p.���î�U�=���|Ӓ������+J�>����=�����u�ۻ�s�p�A�V���0��Y�L�Zd�`z��LdY�:����Z$����둑к�������O�{���σ'��|p?��O�����;�:³��eM�Y "�5pC�u�'Iǌ�*����sҥ���C2��.Bʅ����¾��>�f�*��g�"�|P@.� ��2� 5w�:PvtQ������/54�k���&y~��8�6E�H&�z����e�ل��?@d�������m�����q�B�7��=f#��]e�1�#���C�S�F!�7�W~�V�Ou$�:���'frǗ#늁;�����o�-��0��v[��z��]��ͯ��tt�ֲ���e-��e��ײ���e-���č�O��-6.A�)��ύ)^�{nl���b�*@�)��6� x}�eS4J�uhpa�M��H�����(�IAѦW`Z��@��@�v�����u[�\y^BE����"��t��:�@�5~�j��ktf�Z�l�^T7��l-21m��� ��$�D�{�c�Y��$�	FM�����aI$2!;�"$M��:
1;�F̵ql�-����S��xb7���Mw��u��Ip��#�򓟸?��?r_}����?�s������&��e��a�4�lܮ���+�y�Z�@C 9:�<|�n428�U�k��R��"Q!�#L�$%} �,�z��NJ��'@�Ϭ �O�e�9�A]2�f�yR��%;g��n�5��| ���LOq@� �H�M�O���!G�?��Ah��WI�^�U���L � XF�*E�z��7��& �D���H/r=in��e����>�0%A���c^#���f^��2Sb�'F��1�sK���~ѨrG���=C>epH����l6"cs��#2��u��U_��H�{��g� Z|f8��X.��/J���,5b.I#-�A�k�$6J"����Y�� ;��yN�]B�$*�j�c�sA3 Eǟ2nȶX�Ȝ��1�qIˁ����Mw� ��J����(	ؗI�ި�e��y�H���ݥT[I�ؽZ�^�e�//�<��\%e���)�_be_�[_,۽$�J鮒���,�R�.p^o�LA��1�A�8�%����:.���� ��4�/��B�����KC����H��dT��Q�����f��5!vM���g�̚42�$P˾���k.�$�J����)d�R^��5�+$D����Y	�z��u|�=�6>O�<>0Sk������O����V���kf���Yf�+��q"�ȥ�=��Fe�0����p�F�����¼���k��������?f��U���7����'����8}�g�c�`�hx ׍5�jDn��H�d/�WZ���(�-��'�o�H������"���s3k;c��0�L�d���q�L־#1�4�$�$s~`v_��@vגK6U_�\�L%��~��L�I|_N�9����W�����NGf;��1��e<y%D��Yd]In��M�mF	�	J6��NI,�u�6�-��/C\ӌS"AX�*���s��������ݽeSd�b.O�A��:����x�Ǘc���#�z�Rq��վ]�Zֲ�������Zֲ����[)�kV/I��r�Hɣ��n�	v�JP��'&ؓ�m���E���к�'�5����E�� �RXu2�5z�.�`�i��W�H|n�l�h`I�"e��cHQ������� )فE7���j$8��Y�$ˀ�A!,��=#�H���)[%� �� �t�#��I&ցJ~���g&�Uܘ����� 8.����e��e$G�[�kӊ�'Jx�u#Mɒ�wM/}����@9�q�1����w����>�޽;�<���	N����"���~��}~Ff�@I+�`Cd�^4N%* 5�L�a]B��|�\�+�W���xCao'�)#Q)cջa�~��"֨n}����L���;�w��I�lGȼmz1]�	�~	��X��A1LP���'�&A�1��/BM�� t����K5�o��zv�|��OśY��m����
�OaD��~+�@	�7�ԝ�K��wm`�0��F+Xo�����@��ap��� a}af~<P��h&���(3��L�Z���]�~Ѧ1��RF	i��.�,�Y^�ݶK�fvZ֌ љ4(3!���P����/�K."����I��y�^f7��Ȇ�c��\�-�!P��<��Jx@�
�o�g�~H2�Ġ�g �;O%D�3/*cg�'Q��bv�����(�4Y�M����ϫ���r�����q�,���(��:3�H?#$�I��v���k �}�K���z������2� b��^�/��
���z��+�#���ǂ���[vIVn�̬���&���K���=��3Y�2C���r�X�IIR^�����c֮��GJx�e���s]Y��g/�ũ�}W)�S{����Az2����~��࣏�3t�~���#P����S��,�߈a�[H�I�A��A�b�!�����.>��^�پ��q�^�v�����{}���9��_�=���O�������w�|�rj�fy@�l>-n !*�ѷ��:#�O�����Bꙏ�DF-Y���#t�7W���:��J�D���Ϭ5f�6�y�3�8���IKኮ�zfǶ4�X�.!m��\�L��gx�!�E^k���t�r��Ƶ�@-�%2(��\�0E��NdJQ@tɜX]d6�ܐ+�zS ���yJ��ʤ�H��Jt$�P'"�HyS��I�sj�%q���C ֽ8�L�p�Z��p��ؖ7�=��q�/*����X���k����W��~�w~�
�_	���e-k��� Y�Zֲ���#(�h ��N���N��oaxLJ&e3�����م����R�Y/�<rP5<T'_l�f�;��5�!XQ#���@Y*�J��e3+���Z�Ȭxߓ`@���%(� &��=MkF2B�ᆙ���y	Qv ,�mn
y��S�^�]�qv�ܰf#lW#���]��\ɯ� �{�R@��^33BUSw
 FAx���$�v�q���C�V�{f&�)^7t�����o�ֻ������K�[ܽ����4��6ܨS]'��7qc<3BD7�'��P�
�c�v�i$I�6[W#:v����Y��(DDȞp�A�,�j${��ȍW��В�[���X�
���@�B�c��3���A.�ۭ�{���GY�Zt�g�9�G��[`� 8��� ��3���{�}�G�Z�A��A��b#8�V�0���
T�@u��F�it�er��|�LzKs�k�#;��a���w@X�B���7��|F�q�?��l(�һ�"�1��o����$�]|�"����T��Qvn��T�a k��Q�Ԣ�Ŵ[.��#�2�A'�
5�t��5�LL�K�Z꯽�� ��O)�c���G����ٿ��C���R2��D!�U�V
"��q�  1���FPW���� d 嶛]o����@/�q^NjM%s�e�n��A�����4\ �Z�L~X_0r��A��,���z���(��1a�/F��OJ�>{�����%�_�e;�g�r�zI�H�L��&�H���zm|O��S���R\���N��.�����|#}��6��w-{���&���|dYk��U6V�IJ;��%�dc�0+�Dp>�O�CjWk[�$@ګ�&�y�����|��ܿ4���!�7�}��g���������<v��C��O~�>��$�7U�84�/��B��53从��L��8m`L������u�^+���n����%�D"EX��ċD ��,	xU��1~gO�sf?�L�P1S�͢}���F�-)(����&���Yȍr]|_�>�c�r��(2:�`HסY��XQvd8��Q�&��	��E��t�5s"�[%]�>E �(D�6��>�%��E�r�l������2o:�4$���r���a���	[�X���f�����R�G8*l�,���M�L�`Y/QJ��ٌ��ؔ!����؆��@�v���Su�� ���E2Wq�c|v}��Ox�����vkY�Zֲ��NY	���e-kY�?xAd?�zN��m����Bʨ��!���PRD�|Y��0��3Bz��欮��QLj8 ��������j���8 pb��&��Q�����0ى2ZS#�4�̾���9�$��A��dz���%�z�a�QYg n)w2ss�M*6���Xt��6� n`d�H�GNdPrbD��Pt���F�'��|�]ɍ�B`� �r��_R' 
:�l�7�ٸ���G�~�7�͛�}�W�so޼U��� ����O>u?��a�rsχ�l:� n���;7ƾp!�0���_D�<��'浒V"��Nr+�k]�,����t�� >� �F�ϑ8�wA�?�,	  ?�no)%���A���-#$�9����� �c�|���틌�����BÈ�ĵ�<{�8,nSIa����''m~>��88˳Pv��Y���:7l���p�,������=_G�[�,ec��_L�����.Z�$ ��zb c��\$iR�! �8		�U�G�F�h��Rx��c��h_���q}[�M���e� �L�j�.�Ƥ�,ۣs3������z���e � zy��E���Y�m��`�
M���X�j�A�9\�셺�<G� *5R��2#2K�J(����x�����E$��;fA�=Bf/>� ��]'���̐Ў�%W�u٧���ʺ+��}m`��%`��b��}�HglK%��r_i�^�uy=&T3�dI%���kI��]ʵ�}�uR��4����\x��/��=q�%iTJ�����a��J"��ec�>k�o�X���>�L�6�g��(�;e����U}���Pc��ט��l��z������?���'��[��������+��矻�ۻ�>�����O�(�	)���?q-Ȍ���J�ҿ��M�a`��:�)�\�ߺy.D�/�Y�Tj�9Tx�==3���J�����2�mu#�L��2�ZH8��y8�g�d�Fl��\�\�kV�@�r�R�_����ȉ��EB
Ǘ~�gƑ� ��m��8��ϗ�er��~T���~���sri�j�q��t��Գ��ߨ�k����`���(l�;��B�P\=>>1���k=^X4���1�qu��$�_��$Z���E�+}a��u��Gf�n!��LcHt�Sf���78�M���75ﱏm/���꧿�>xu���K���7��|�O�%c��>qkY�Zֲ�_�� kY�Zֲ�o��d���#��6`�"C���e�=^�Q�;�~P=��(&ςM!"޸���` R=���i�f��g�q�|�ty�K A��&�rD�a.����x/Y, L��a�ǥ�&�� �`[�̌���D��y�
�f]�'�͐�)�Ԟ�����~�xຘ���"-�j5���V�� �ɮ �S��^D�����eTp>)��k���	���X��wwn����tp�}�}�����_ߺ����{|z�W�vw�~�wo��7o���{��>������)���Ͽ"p��W_s�N_�؞��S�����g7���0=�!5�n\�[�s�����5�9$]�����{�6��`:���&�E�q�X�CM`����,Ha�7��P�������0z�f��]��T�|��c�'tZ~Ѷ�|�&��#�9`�x"@/�8`���0���(`H񇨯�u� pS��~S�hJ�\����*�e`+�5���~�yH� �G�x"�����I˜ �1�8"u��+�#f��|�80����-�#Ef�����J o(�qo��*�$ϜH��C&εN�d�L��}��u�����x��̙%�&%���G�:���.e�J��~#B����έ��#1h-��<���V���1�g�d��9�(��J����ݰ������Oa�u��4���4g2d�d�kI<6��wWK�6���>�q�����
F@UHU�U���,9c������H��8�R
%9v]��Aپ��k�cua�|ٶ�#dޗ�b�r��~Jr��B�G�qj5lv�wJ2d	WY�se��J|,��t���~�x��4f-J����T��Rެ��/D�!��q���l�ZǕ�����\��/��Kr؞�(֞F��}e��2k��tI ��D�Է{��dq?�_�~��O]�s��|�)̻W��{#�m�����9��g�3�I�a��si�� �v�lT�����TN|�<���C���_M�-+��s�F�%����=���4�Y;O9O��c�,Y����j������RL�/����ͣ��d���
���Yj/0��	_0�0\��� !�5e��[�lg͸���f�����?r]:��"IC0I�p=���H�>�H�$���)���HL�{o^4�(�s߲/����>އ�6Ȥ���~�W��H�������˿������-�O���L�q���G��埸_�g����_����O*�±���H�����;���e-k��,+����e-k�V�q<��L�!m�a4`Ol��@��2?�똤�m��x����t����R�t'��Ih^���O���xllR!�ID�_�6~w����K�H�U���}�PI_��9lU�Ȼ��U���
�y�$�B2��~q[�[ q�I2Sr�y}�*��lF'Q�B���d7���� �&sk!@*��~7�#h�G	hZ�C��ǘ��������h�y:��6^2V�(S��m�>��C�Ŷ�䣏�	p`�M�����|p7�>�����m<~����o��h�o���6��\�X�N̶��=& �؇�)���k��q�<�,���lc���O+�P�
Rg@r�0�vӸn��J���$2?��� �A�}%�P~$J�'&d�w�o������hp�`q��ν[@4�ϝ���v�4b��f�"疣���S��(croOo��/ē�vF`"Z�瘋��Hh�s29gt����m�����QY�|��O�ϩѩ����c3��%)Q�e>Le�E`���� �C�S��@5��&i�1}V�9�v�g5����Y�^ă$�+˸D_9��N�����(3bJ	���r$x�Ab��,��|-�:6	���dmh擳̏L���t���zD;c��� ���q��}��[����T	i�쫾 �p-� c]�� �ΰ�q�ɰ8�wq^�޿�Cn�12����F:
!�Ë\��̟Y�TxONM��~ "� $Rր[�����x�(��k	��/�u\�]��3��CAܼ/��Z��Z���:M�sv�e{8�s�L�H"�1��	��hޫ�|�Kr����H��3�M�{.lk��k5#�^��9X'�#=  ��IDAT�>�II����u]��T�W�_9�l.������\JB�ƫyA�c��gId�� ~]̵r_�mR���v\f��y0t߷�:�����m#Y~�>*�/�������a2��0�D;$�&�z���Xc��H���.�gMZa����t�ϊ�;�<�m+QO� )�y̪�I\/�'�m���C�FI�:Ɇ�������� �r�_,;����>l��ct��;}����f���UXSp����ސ��J�2�g�d�Q���gnnw:^b�C*(��@E��T߼�����5N�8����5��5��:p݂G�x�"O�NN����[���5�Y�:�$���1n;�s����f�$���[��rhA����������ٟ��6�������o�{���s��H�>y-������~�~��~����K�������}����o��?��{x�֭e-kY�Z�{e%@ֲ���e-�(����j����l�j{�ݍ��M�i�6�v���n����$2���(7D���f�x���Q��h��F�a�7� ƿ���h���7�P���nO����I�G���ZӂW�J���}��q�G��%ق��Y�X���� �~��'J����	�aZ�p��&�!n��������� 3l�[%v�w: �]K� d�0�������%��#���o���~����lR�F)Cv��:A�a�&�)n�*�'�hx�x�P�oBs����S���L�����nonb[<��~���⋟�a�����?����,���-͸�7޽�}���ޑ��~���{�����ѽ�t�q{ӻ��w����#��5[G�e@�oZ��P5S1Js��Q<~ ������ܵ߹����D���A����7��:��DB�C��vۻ�-��j�S�PM�!@R�w.~���f�ۇx��_�c|�4����v���yx�lz��_$zf��ȭ ���^b��/Ʊ"�K�q��.AT���"#������%���F��I�J�Wi!��{|~��tAZ��9�3a����k��&8�c�FV����=�D��Xv���DV�I��Y��4���<��l����4 ��z�SK�sx�u�^!�2MBZ�ЪܐW����IB�8�,m8�[��	�JYSd����؅�p	1vb�+�ў$�5d��4���P�`95�tQ���D@S�΍~a��^�N�[�QyB��BB4ef�b	��k�� ���w\���S������oc}l�u��H��/nw+5���+�$[��oi�qzHѼ�QՎsՍ�$y�P�|R�
̛��c��c<��>�7�vv�����nn�)���8�?�]�l$%)��u�L�M�.� 41S������tF���k�.�Ɍ�a	08�L���lu�׎/��g��lO=6�ku��Y�� ��'��c��┼rُ��6N9é���%Z;��9ɻ�27�݂<�p���!� M]B"��[仐f� ���g.��q%�h��O��� ��Y拊��)����̯����H%�	+�Q������q"���Ӡ�p&+@��s���0���Ax%OK��d��a~'�ʞ������<����Yƙ�UzN�n�,�g�%�!�,�PJ�a���A BǙ�%6vh���ߑ���ß��xo��G�だ�R�S������I�Y3�b_��g�e���9�j5�f*@s#X���1�3��MG�s�9�Md�����s�����z�c�L%}���d82H�0�.�s]��e_�%K6�4�v�.����{�2GZFާ�JM3r�`\9�>>��JD0vٮ��/J���8���֭��X�a�;�⚨�m�qC�����5 �v���q��X,�م:G��H���9�.�Z����R�Yq��Ʉ�u��YN�y�;XH�L%�1�!�����ɓ���졏��Al���g?������}�'���~���Zj������$�$�!�<ly���d��v��W����ܿ���α]?����}ׁ�x��������C����e-k� Y�Zֲ��|�eĦ��	�b��@�r��77ƕzNT�<�M6l   �`s��v .��B�n� �?ظ���ع�ݭ{7ɇ�gfl�7�Ň �DKCjH ��x|�sT�!��f�+о�io7�[j)w�q���yOm��#A��n�3A ��_�3u�U�k6�����nZhD�B	�1�M+z���D�(�C�+�����2Ar�P>8 ��n"�����]���1!9���e�#����e����W��* �N�2\����ʟ���I�y�ȇsܨ�k��A= @˨��������0�����w��c]=��e��x�^Ǎ��f����8���D��l��!�(}�v`�޷lQ���ƣ��AL�+'����N#���f��R�r;�O�8�5�F�f�N���꟣Q��JD�b0���R�z�����������5�������zA�S�&�&�B�IwS��c��1�' ,�M�.��I^��E?�\���4ൌ�7��Z�^G;�yK)�2��4*���f89�^i�F���&����xߐ��n�5��I��A�>��s�Y��[}0�}6����f�Q���r��*F]��%�ę&d��>�̑5��,e�Ay���|)D�?��� �ȶ�,m����\m^+?&d&a.kA:�]�(��mA<���njFw�yp\B�-,c����8�3��{΋���Y� �K��}7��@��y8��͙B�v��͝�A��;W��>����J�� t!�Ez��$e�X��BI(+��
��I��^em��l�J���,���قq$�\��n�S�������2X�Z��bj,䉐l�8N�L&�B�_����4�3�|�l���EK�I�1�|v��3$ϵ��ToA�U���d�ʌ����uFL�"������fs�~:�G���Y�U!��]��]6?�2\){��A�X&��C���\���{�uT�X��p�T���o�����M��_s=���6>{�q���x>��o��sv�g9�-�u�lE� ;$��w���8��*��yv��x<�)��%�qH0�q��쿓�XAB��2	[If�8�܁�fzWwB29�ׂHk�3�1 �񼥷��Ka}���![&n�2b�����Qο�n�-ʇ9��Be�\I���"�m������#�~��O�#	 �#[d�8���*�u�m0��u���rMJ�ʧ�W��q��a(�K�O&�˪ğ�DM[��U˶FV�D����3�4�:���=��E�a~G����x�@:�X��p�O���\������O��Oݏ�c���z���>��]�n_ݻ���Yp���)��&~�/�ɊϘ��!mײ���e-߹� kY�Zֲ��u7k�Ў�l���9ܠ5M�K����`b�r���L]�Fe�+���x2j�^��K������f}�ٸ�W��������9Ho����1���ћ��0,^2?@
!�w#�I���g:n��"�x>0����fR�5#�� 0�%��	.��@�M��ОQw�5 ��z���g�F�W��f�!��p�e��^$[&����+%�D^' �JnУ������%#��=�c��3wBXōq�&�x�����OC�
�9�܇�Z`�l���ow������	�����Ͽ�;��7_�!~�xz!P�(BD C�
�s�ݹ�?�X�P)�"�O�G���|!���+�,�(P�I�,˥V� õ��b���B��'�3ZI���Vb|^�X��x��*5����8�H�1F �����P�Mt�7��ff�x���@s�6@��,B�D#2J�����g���5WӨ}E ��6����JY��E|S��Wu��{�dy5�D%��D5�9�jL���QM�̡�B�nY�j�#��S��ْht!k��v7���|�h���^c@�������$�e��A����h_/Q�b�4�^2�(3�%bx�����ͻ�3]C�� �,rct�H���å�ɥ��WPL?�Y�G�J��$������!y;~E`q�-&lx�Lg��߃�m���6��34��@�L� �@2�M''���F�g�tV��@0�*��j�}���̵J�T���:>wb�� }�'W�v��^�v��WO���޴˒�:����r�@+�EjJ���3�A�|��gz$��H$(,�����������$$�,�8M��$�*3�{��f�̎d��t�o����ژ�-#j��t�ʓ.b�	A�[!��#��م>�yXK5�@�ܡZ����c+�|&+�X���������g��Sc@}�^�C�;�4D��Բ�k�e�P�f���J��gs4�¿�ɕ ����fIef�S#�{eLj�xG�wU1����:�Ϗ���T�5��)�Qq���?�5���}D��1O����<���U����7mm�W�����}'�bL��s����ۜ�Ŀ���kw��������fY�)+��.^K��왭�1O�piZ���6Z��B<����_U���QIK.���Mjy�y��)(Y�چ������TAvo⽈D���S�CE:����ގ�˸�s��[�ȷ5ZSye���XBBAm����L��N3ޢ���0c��YnL�g�(����!�f���v{�������X3��H��������5TX,
j8�J��ˡ�O�ܒ���U�ҽ���b��`}Pը��OB��A>q}���J�a��{E�>rZ��e߭�,(j�7��Yf3��}�������K�g|m��mn8��C!��Fv�!w��=ʼ��s��ws})��3�]�1���S�h�"d�A�6��M�ϪM�Ԧ6��M�in�$�Nrf �ߣ���((�0 �q���a'yY���������"�jH��n�U�b��Ve�-:�� ^h�������_`+$�x�ܪ������Xl��77�ib��\�$>���&����$
�Fj��+@\����nÊ
El�slql����4�^�DI�D$�����
���]DD���6%��\�r����\.�/i%������A(򒿷Xئ:Y�Kr$�\4�~*�5�� �fT�;�^�*�-�ʖhE!m{���x����oHtȽ�������@/�/VK�Dj;�{��_U����m�3�^׿�\�S�s�ݖ��<W�l����bIB���&1�Y�󺾾���+)�7LJ, @ Li�i�X�ʫ�*뻨��8��Z��j����}�u������=�*n՞#\s ��T9���ʉ	��~�������Z$Q�F��=A� N��`'�[4ڏC��>�,�x�5�.�c�r��$	+Z]����fPJ�C�Ǌ�q����+s|%���������>@X4�^�Jcd���ګ&Pu���<��$e�xN����RV��Z-uF
E�m�{}X<�5�;�<���G^��+�}�6���n�E��3+x��B+��d/>K	����0�@�c�۪����*�\���b��%[�(�n +�a��3��n��������;R9JP22���p]&��X�Z׷(���\� �j�9%Fj��TIz�E 0�*1N�1R�D�
%j���u*O2Y-S�U�>����Pbuu,��XN�KY�3y������_ׇ*'�^��^תn1*tM��<Ԁ�ګ5�a��_C��+���C�ѯZ�����z�-����Nt�	�@m���q�F�Pf���്S��ꉰ�߭��� !�W���	��+\Ԋ���*�p�$�q�
CSWIx{L�Q�������
����cBۿ�'	@�z�&��x���|����z�Ȱ�k��>��k<O�������q��[�����a��~?�mL�`�B�C�ٮe�杪5�U�m}p��},Ѣ�DU\$���(���
�����M�F׊v���Ϥ'�EI���̦�RV>��F�8��ܚ��5�BA��ٯ	oYg)��a��z���� ��	�a���K�����Q�5\���&�dQO���8��&����Ѽ��v�4{w�;��q��śs�'�U+X��Pť�rPȝ�*6|��lz�H�u�ݸױt@?�l����5B�K!�A�j�y9K�q� �I@vJ���c'c�;���kC
�Qޏ�<��lI��NkX���� @��û?x�@��N��66�^�~)����*_}�%�`��ެe6_�lu���F����l�]��W_~!_~�Lf�+	������'��nL.OmjS����<�D�LmjS��Ծ�v�m��`]���V�N	�V�f�T�]���۴�j�8h�2ø�埲�0BVH
�a�&�� T���&+ޑt ��j6Xfհ��܆�@���Ե�AY��y���m�
���~�y�ԫYMWI&�E�T��b��$�
bۅ
^l^��У�JO�ZͶ��|p��@+щ��)�98�j �)� �� )�c�iXe�������=���#rM�_��^�>xw �����{�@Ff��h �=u=���b\��l0�N�����ɍ�Gl�{���\�X���1��p @@N �|{��/8�{gr�P��zZ�	7��aO@m�!����马�39�w*����Y��i=H��aG�x���F�ƍ9y�kW6��U�"�z��*�*Tѐy1���*<�h奷�aa8�F�(�8�C\��|I�o��x�9'}E5�"�v�{���W{��`���AԸ_8�گ�h��M��^+�� �۰�טV8PZ�׾��խ�^��싮��@��J�߹E�X��z�7T�k����R�TC�۞�Р� ��"�F�7z�*ᘊ��]� a-�b��n~Җ�M�Q5�X͹�l���d.)0f��O p�<�d�!�$+�Y��muh�Sk��+�����ud��Y����CE�2�F��:v�q\��!P�S�*M:U���TJ��$���!P2�t�Um��:���H���`:w�Rן�8�#��ӑ��-��	>:���׷�)�D]kj��� 0��WxSI@TV� |N��d7Gv^֪Q��?���<7/ևڍ[w������Ir���x���l������3��l���Fxp��*x+ ��5v������u��D��:�������׈ї%�t��O
�j��
x��|�<։T'E:�1���� �W@�����G�t�k��𕑮1�^�+$��jپk��夒-��1<&	Ɩyc�o���K8���"ʫ�/P�1�'0�4iX��r�x��/��Tp[��	���n���=Uo��i^�Z�DM�Tin�{,iM�
��EI��`6,�p�(�й�w���̑��+�� '��D8o�/ü+Z��̍�:�p�,�C����+��Dm���$W��M���j*?J�w%�͐��*�����#L�ۨ��)��[ک��mPL&��AO�c����`k��P³�I�h�9��V��P�Ah�^��_Z0b����P�91t����77��R2���yv}5ȼ6�ge�u�{l��3W�kx{>15�Z��bQz�k>~���=3P�,d�4I+�b-Cn]�I�g�:TuN��r����{&[����!����;�+��:*L��wz|̾�����R~���$�����|��O���������e�'��7yQ|�g��/�}*���������'��E�����ǿ��LmjS������D�LmjS�������ȡA�X!�]#�w/$F@9���&8�/4�B��=���\�cV��ݮ��}h�[a�{0ln�i�ͧ�s}�f�66��t���<WP!Q%�����vAQT�!���Z^�~�M��ԉ*<��-m�D+�Y�|La��noy��<��$�i!�q��VW+Dd�tns���tF�����>Wdg ?Ȃ(Ҋے!��tn3e슗�E_��U�17��a�+C+��CxV\2 ���z�P���. %JsN�r�X�ŋ���N�#�i}�������?��?|�>�8GTF��kV,�Tl�2s���6�{�~
^�k7F�AxY*)�aա<~�@�p�f�HZg폼�����A��PiK���ĪJ�ȫ�MP��jku�h	�Oe�7�vu�������\	�������o6V����5�����F%%�Ƀ�
�N|Usb �P	=X �(���?Vكt^��}𽅋o�a���:;���<p[F��|��/B%�<��6(C���/B�=�S�5�p�T��)�69nC��TY��Z���}�t㾯}���ҫZ�0���~ng�6f�����O2x��[�j"}_�E�g�v�|o��/.{��{�+pk���Ǖ�O�j 2r602F�b?�o`����(G�5��ݺ�"7 �7�G�V��Kŭ��a��1�.n=�{���C������L+�-�]�\���g�w��cO�X�[�Df�� Ð%�h�6�����AL"Y�P�R�nw�g����r%O����y����z�1��6�.��3�rlXM���&�q���Ѿ��hߚil��m�������%��㐢�@��� 4�.[#F�?^��꡻6Rc5QO(��D���HT������d|��fwu�����1�J�����o�w~�kV�χ�VqA�{����ր�Ϙ�����-��2��� ���{������w�����"6��0���\ORU6$v�Xd�:ük��$�T�>�j1���l���0e
�C�� �!�-�`���{�G�z.>�	��x�*-�����~��y�~�=a�V���8�hC9�wh�I�~7����U�����ϙ����x<�=��Py���,�tN�׶���$��Wj
"Ñ;�w>�R�0�V���6|��ĳW��q�/������5V�" �q;|��J"f�@�����u����
@����O��)�AY���|����ɽ{�8^�y鮣����4H"Z�\[�D�t������O�����P���Yu?�˿���ӿ���k���u9�?^�z%�������<|�����ó�ӧ'�^0�A�6��M�ϡM�Ԧ6��M��6��j����__]K�6��<����<z�X�YN�9����`o�*8�x=6�P\�_��Ņ����8�"`��3��
�	���-�F���Jv�-�媚ӳ��X�x�៭��~qq�L������TST�ɽ�U�tbi��������p9��_�����1� tlv3�fv�.c�Vv�����Q�P9����Ш8��6��`^��E;���Hn��7V!�X�CM��x�G�m���M�XV�V�f�m�[aq#�p
�d�F0T��%��7�̨Ȁ2��wߕw�yGϲSr�Gù̲H^�~A�3@kn�k�{<��3."U�j���ȍ�[Y��̔@� X�r��(Q��G�(,�d4�����KKK	��;�Z��n��\m|�J��C�+�JK�C�5!�'#ϴ�=�^X��c��9Uk��j��Ū����RJ�,����b��7�*��9�8�-Z A4 �c�hl+�A@�{��	�/�:�	�!�\��1���Jo5�@-�b��?��� �p!ǵ'@|u�ν�����������
m��"�A���k*rH��f?���ط������`!g��5����C?WACO���د����,dބ*x�^�Q ���o�Cq@`JY*��d�~� ����e��.n*�|VT��F�ۀ����Ȳ"����!��=��\�y���F�����n��s����b9KdLq�:�#�jH�L��* �c����Ǎ�ZԺ�/�~����kP�t�/��p�+�s@�1��P��b)�o�:���]���ǲĜs�V�>��.
5� l�hP��v��ӷ�c�?���F��T��ͷ��V8��*��-�+*+1�Eo_���������]2�+�8��F�$��=!�I���*���օ��NwU�	�>�k�4&)�c�1Ys����
��Z��F��~l��5�j�c�?�J��4��>+d�D����:��` �z?#�qߍI�zK�?n�~�Ċ�{!ա ��:+C�b�C��|��Tn�ơ�4$6BU�5 ��p�=��j-l�S����N��u�qڙ"������ޓjg�yd?d��p��q]����ec[,���qȭ��4��8��} �B#I��3�$Z[#���&	��t,�*F`���8Xv�br9w��Y��P���P	,�Ș�rdJl㡳�jCb��B�O���׵�90x�J��S+H�����݃s�"PC%�Z�B���	�8e<k#�~1��~�wϚ�ȉB��E:>w�jԾqL,��������~�0�;d���ޓ?�H>���/v\/����7�y�z �A䩂�S������/����ejS��Ԧ���&djS��Ԧ��6 � a�o������O�����+Ig)A  y�����Pd��2X��{o^�����g���䛯�a����:`��U6#F#I	&MNK�����r`�����m�����tN+,�h�Uk��j{p`{�~g&uW8�I;��ΰ����m�#�%��܂@ p�Z%w�mQ|)a�2�V7��5��2vH 1�Tǈ-V�À����%0�+���Z�O�!7�>�U�4mȇ�r V��#Eh� ���Sڿ�k�� Ti!�6��<��e��ܯ�W<�o�GT�<}�����l�q�[5���qpB�F�L���;~��F7�Rv����;��c��Q�6�n��ݵGf�j1w�-�kn�Z+���t�9��)�p,a��7�jm���F�f�`xd��>"��>�{�#G �G%g���+,���K�	 �� )h�dh �Ν,�BFԝ�@��� dZ�b Y����ŝ):�ϳT����O`����Ѻ�ϯ[��2���� i��b}�՚^��m��7������F�� 彷�8+c�������N��0ݞ��B��c��u���"l̰n���U\:�BO���O&=�KV������L1.p��s���W���~]U���8��`]-����$���[��X��;>��W	M�Z�7$ "�77#��O箟W���Rއ�[�
�H<f���w�YC�n~�@N���S��a��\ؒ�8�w��0�a� *y��c��RU�d�� �~4& u�>��a���]W+�߼��o�I�?���c��w-K8k��#��������m�Y)wA����<o?8����?"@|#��� �����W,�^��=	���	]�����ԉ���t��4|=�`{�+����(0s�����,���׻��u7�B�w ����	�1Y�mꧡz��������뿟��s�|����lG������m��c�?������������z�����Up_�EC.�����f��ם�����5�aG	+�(�H*��/��qh���X|��=�E�)�@��7U�r�/�58������m�N<�>50�Ͳ=�cFQ���;�EI��o��T}�R���<�q�c�u�3���l�5}��G����w�����Cy��[r��9��MT�%�<7S������{ƽ⽶������'g�����w�W�1��Y*�L�D|2�������3Y�3e��e5_�gw}�0�{[*�z�vru}!��s��W�p���ڠ�E�4	�3�z�|��\U,u��{ ���r��<y�<z��̖39�w&�W���o~�+���"�������s��LmjS������D�LmjS������K�ߏ	=��@>��#��������l���k+�2TC��9l�Q����#����u ����M�l6w�X�_��#��;����r)��^担�[�2Cu�bN˧�-Y%Hi?�#� ����C%q:c.	6j :}�2���a'��쨃�P,!�Vi���M"UY�s`�r�7�g�,�eR��;l��Rm/�~.�˵$$j���GO�i�Er}}�?H��^+����	�����G*&��6>��3��l`�p}�<ˇ�{@��, z���l��6�J{�60ŉ�^�Y���
J�F���+;�s����/\�?T  ����J(N5�J ����s��K湜�q������土����v��s(t�N��eu+,!�ʍ�1� \������f�U�t��P� �ƘD�t��������-kê�$�/$ucD��[��C�A�m���[\G�#�d����-�`R2"G�T��?Ȟ�OT6���PhX(�3T :��|�q���$,$~+�+w]҂}� �������U����}� *��_����ὅ^[oC3�#��{ c �����
��:a��r$=؉uăg���o�cb�j��F�H�*b�zI��� �����P1����gAeO'�L	�ؔTh����d`->;
B[2!M���6R�_�liB�)U�^/u�}� �l�{z �J�dP�x�	���'�+��6;7.{k�Z��@u����,�pz�wI�2L:�����º��#v�m�~~��|�䘬n���Aƀ�iҺ���8m�Ƃ��T Y���;�6jX����Ԝ" }q� �`�Y?�B������p�����X�"��%�j��uC�'����sǅ��bY-Ri��r�է����?}GN�y����}~Q�p��1�a�Usm�8W;��T=�D��9l�'?���b�3��Wx�+?����H��+wh�o�nГc"��ê����� z�� T��A(�f���A{D��b_L,�m�)�ZI�JF-�0�=A�`f�d�Z���yzK�1���+���+��Z1(�1�t���}~;�����Xx�_�[�>�yh=qq�Z�.��������{|��q���w�N������o�,�y9�g]��fd_w��d�0����u��?��G�w\�th?7���"IX06��s��* :	o��֍��Nm=�Զ�=��>�=&8ֿ6�ع�u�L/ �s�$�� 񊫖$
�Ǒ�MU� �{c��sL�8��H��A�Ӂ�7����x��<S��9�[���eQq��T�$T�޿w_��o�V���}�-r T����{k�(	����T�^]��չ�=�f�u��!�%P�b��o�0�L��sy|��31�������П3>A���|��sy��g�������G��Ɍ_BM��	���l7�w�ǧ'�����k��g��������;�5!�?q��o���5\����|��{V�.I��M�Ԧ6��M�ϩM�Ԧ6��M��6���Fp]b���/�3�����+��?����~�@�Pu���}O��o�����?��<���^Dk���~?�����{n��@��f��xI`�F��  w����\�lI.
*+z3�+ѡ�H�� 84ʘ�CaU�Q��2-��2���`%��BNVGT���+�e�6G>I���V�߼�O>��|��O����R0LWI ���6ۭ�+�Дj��7�ncx�6�g��>z��I J�7�j@�Ax (�Bs>hg�Ԭ �*ҘU���A���f�U����Z�V g!@�a�lV��:V��T�A..�===���cM�x�u��6��<&����{B�r���=��������U� 鐓� u ��M h�6V n|$��RD���nj�*���	v��Q�{=
��uۃ���C���p �*#� �XE��"��\_�����_̮,I��2n��k�J����zG��^�1Vbp<�u#G<��AC�9�����+H�d˷���z���=���}�G��=�7�����րѺ?���~�쎿�D�^��h	Ya�����;�����=T$��h�cR�&@�Jڅn�i@z��y;>Tw��	�ų/U_�U۫O�u���X�1�&�����ʡ�T�,�D��a�ư�N^�yE��@5�>��CP����S3�F$M!w���}��ӊ-���l:��q�T�0��T��M�W%�ș`�j"6�$�'�VA�&�9D�7��\`�ZD3;�v�s���
W�lO�F�	�,<�V��������zy.�����^H��syvϭSs�G��kX$b����h_�{��ڑ��E��F�#-��`�aa�8��h-�~���n\�F-�t�r���f �i��i^M�s���|j��HYCI�3G��C)�$*���4(�a?"�=N����S"��]J��8w/rߘe'�^��ڷa����pnDEK�jbv��A�1V��U�{c;��fK�����L�~[���|�����Γ-c��s~-�_��6\w���kߦ��Oo�|�*��Rq	 $nz�<T�S���_7V�Q�OBb�᳔?7%,�u��Km����N~��ͦ�"����N3~�\���r��P)Y��9 +[�N�>�l�&�o�$p|�o{m��p9���i����eȷ��7#�C�r��[����;g4�#��EF�("�l�U���ީ<}�]��������fâ����%	�so4SJ�+̬+�g��T��O� sϏ������TH�>��gL�H̒�g��=��I��S�g9$��%�gܵ�Ry�䉼~�)3��lv���=��U� �#�����?���뿖S�����߹1��	�Yw/�d^s�ྼ���_���{�/�����`5�����\�<}"S��Ԧ6�?�6 S��Ԧ6����+�]_��5N�l\ɛ7����{
��U���f<�X�C� N���P�nS��|D���o�����<W ��(�Ǟ�}X����������G��j�� ��=q~~�6����߃-�5��e��T޲���I@�� }vEI�:��d��x��ձ�����L��w_���r�b�.*ٳd�\����z-Ͽ��$��j#�ߜK��� X�Ѓ�A0x".aۓ�]K۫�-��+d=0��G��OZ�8��@�"��V�)�t������bB��V��,�> ��l��\��&���HNώ�d���/�u���>;���H���ؔ# ���\��5���%�%xP` p[iU9������4��,4���J��Jd�?�}�C����էj���WR��	�a(�+a�-�H� @6��I�9!D"J7b���@��U�3捠�䓻��z�34���t�]F�(�1#t�J�����@S�_����'V����ܛ6o����DP
�ld�٨�enEM����+�C��j���d�)0>����v�U��1 m4`>���@�!�ni�(!�����A���þ$��*���z�e]��><6������?i��U1P2d�V��B��Lr� �A�M�DGb$�C��{�F���P��;�R?�t����̢�<ic�|F����=��vYj����Iʮ5RH ��A�����,"I	��X�d �{ưV)��� qs,w�/�Q���N+���
�(dLF��/w*X[}p-*��z�EioG±E3�%4�=�,�7�M��²tO�����:����-N�A� �I�b����kp^xo��E(��J۵���T��zTH~�֤{{	�}`.�w0fAX��m���� xc�-���t�^�w��9-㠠����5���4�-2�#TɄ��ܰ%V�k�U .��Ϭ%2Px��c��ﷶ뭮����vaXsA��$i�	��9�<q���Z�#Z=��΂JP(Pо�: �$Z	 ��l�j��q> �*�,�ȝ�߷wI�[vC#�,}��<���q󠫒ޝ�'+*%0t����_��!������5ɏ�1��+E����y���[��c�,�ZM�	�N�)1��{����|��kԘ �1R��Y�P��.�=R(�j��g6-�i�����g~����%}�F���3��π|��h3s@�ϭ�TY��%�_7���p���W�X�Q�[��x�Ț���<�<���0���%�o���ZrN����������7�2��\�gD|}��J�x�L�P=�JV@��� �-�Dp\�Q$2���a/���[�q��H�D��
���i��%,D�߼�F��x��졽�K5����%Pk��'�Z$jB94[�%�[��ܡx"p�T����~(�=��}�jʣ���0����=�e~�*���$��9�>��%w~���ȴA/���LmjS������D�LmjS��Ծ�V���@l�6lhuy��/�˿��?S�pM�v���!f\���r�ҍv���@e6i�����?��g䷿���P� ���^���m����=��O������%�j3�z��g������/	<>Yqr&��WnSVD���!:�'!��j[,؂���7-�� @����H޿/>t>p�*�yN�!@�O�T�l.Y���z-����@�
�[H0��s�����Cc��@%��R�k)>_ZZFŴRH�I�JYXuT
��
��Ɓ���!߲ Azk#����S�ி2-4�� -"�f��,�ܹ�FĄf7�3�Ưܸ� �ʁ��RN\�%�;��c��˒ �ʽ��}�����V)�].�l�"n�or�~N��pOʄ�����A�'lo�lx|j	�*���X{Uh;�k��ڃ%��i����&""�t�$��w���W�泔Vn�4��h�B�8!�ju�����e<T����R�&l� `С" ���'�b$	�1����qt>6K�����ɇ�r�Pu���$C=����?nڱJ
�j����<M��1�/�$=v��ƀ�N�Q�j~��܎�z_�l��a��� �ao��|t�@Pg��r�c�ً���[��n���0y��������{qF�9�E^{SyX�43�@H�=�^���a�������{�<�-M	B����%V���e��D���ꢊ�/@Ů��3��E�J���`���������r/�� A�j.4�j+v�f ���Bv�lf6HFKݚET��Q�� ���Bw��,�?M�I�TEE�*�3���v��G:��SA�ɃϮ��̹>F6���R׹��l�_K�u}��B�q.����kw}wn�nA�J�,z0����-�.//m�wsg1W��p�򯭢�[�(A�d@U)p>.�mM�*hC�-r*-��<Ќ�����vP\W�j�g�^��<���o�c��qo9Y��^�yI X�)���^Pa�n}��F��V¤} ������P{�|�
����n��o���E~}�Ut���5�z��~>�4���>@}�y�T���0h���nI���!]��=�b�E>kF	�e]���/��~-�M��Y��Eٓ�w�||��D1 l�Fÿ��[$c��$�����q���y�y�g��6Y���@f��wG\G����ζ����l�z�[�?�V�^{�H1\7e��Z2���$/q��1��ojd��\���}��je<�n�Wc�ZZ|����=��(w�[}>�3���p�l4��>�I:q<R��E$����Dڸ�Rd�#�J�s��#|��ί��2��|1'�|�mY���6�-|�i�*���Ə���',���-���yF�NܥN���S�?h>��D�?H�9�l:���_=��MmjS�ڟ_���MmjS��w�P�ՙ(=a�����.��ݧV��Y�Zd2��P��{�n3y�������<򓿒g_|&������"o��Da�b�w}yE �������6���״�������#ƦAǖ��-8��pШB�W�H��G �c��s�Vy�� #-,��T�x��:���X����I�y����m�-ϡ�|u�U��ZEX�t�)��&�C��(jY�4�E+�����Q���|�2o_�Aj�g�G�Zj�D	����V4�V<Z��ڔTA��ve��qH��g_������`?��,rT ������ׯ_���^�;���#w�7���3"T#lY ���'��4��߅��@��
l�Ԛ�}o���=��0p���پX�<�= ���#!TV!�{�Bz�{�]�0̖V�_T�PD
�A���^̈́ >�*P��0� m��ا
 _ZO���HY5� ��P1���>�\To*c��q�3� � t%	e������Qa�i@���A��.H�D�=��@�T�؉:AT��A�6$@\߬-�ZmU �R���F{�Y4M)8G5I(�k�'*�Q��碒�M_I�\��DK�l��^�8���CĥEZGe�ZTR׬@n��*`9��9G��%�`�;�`@�������\�eJ��@�|��� @����-�Z���n�/��'�Tv�8�=Qw�-	X�| Ѻ����eJ��i���-�9�w)2� �r���E˝1کPk4��۴��!gD\��9A'v��1�r�P+�)���Ø�E��lE%m��CQe�)!��c���p�Rjd�Hɼ���9;^J���.>Ty�;%���6���)�ǩT��q��2�9���J�v�Zv�V�����a�ֺ�4�����qo�/򞰌b��em?��}؊f���$�Rc*���#ҽ5����i��h�K(L�-�7k�^I�ui��8�@�$$:2v�~_�y�us��K�=4�5G6��U�1��~��PH�̶*�c��ȷ����C��?OPU���Ǌ'<11��������t���j	�!�>C'
�L��J�p{O����n �_#�3G�9�U.J�ǭ��6���W�$�wQ�f1�n~�ujEj�ĻZ��x��Ŏ��gyM��*�F�T�R�
P�p �{���k��^S�@�DP�֣|�He���ޛHh�'H��G���m,;����mJ��y4�^�(�k��'�{�b���Ǣ'���Ps���ۉ�eU��YmGKS<�"�	�WX� ��J���qP�D�W��f[��<�ܨ�A䚱۳O�⇚wW��u�T�2Uf���d��,��A�J�
�nP��DHe>c�=ț�K����څ䋙,�V��n~'�Ƶ}s��*l�s�L�F��ކ+���m�q���kؚ�x\��^I��\��ʝ���������?�9���S�Y$2��MmjS��o2��MmjS�NZ9���2e>�Y����������[��I���
�g_�؅ʁ�r��<����0�P>��Cy��w��g_���j�0��cl���b%�����y�F^�~!U�0�u����f�~v��%+�NYV�]�����U��3�k�L6�
��2�Pq��@^lv����|�<�� t%���Vh+�+���s�dz�[�w[�_1+�P��mv�����^��Y�߭��%	6�
\�D�2�$[d*�=_��6�X��Z��v�������$��9à+_5	+������8;���ЏPB5���g�˯?�؝�V�{�1mX����)� -yʍ:�XP�&�P-Mڤv��Ƈ�*��ܪ}ۡz3<�UAr�_��AUq0 �%��s��pS�Ϣ��P��lw�,1`#	f�0
���v�vmw�r�`�����d"M��r�t������[�j�e�K�vA$���B���3A��v
��螌�j_�ޯ޲k��Cc�O��q�ǖ���¹��� Q���W�A�)�vz�Ò%Թ�Yj��Żu`���婢�����������
�N34�m��ZDa�Z���y�W%	�]q� n�ɮ��q�*�6r8o�#bЃ��6�ϡ  y냗A���`�U��*��Z���$���h�c�+��}�X�1(� 	�TRI���ʭ?xO�Pu��U�B0\��,7�������#@�PV�CO�v�3�@n��e,"2"���n̈́U����	���D�'"-�B,|[Ǩ �Z1��M��s��	�O�,NJ�#Ŷ���c(�2;���P��ڍ��n��c���6T�d�춀sV�#�%��
���z�A��Y�F$#� ����~����+a�Ē���*��0��'����+^:�E/��g�'��
��6b1-���8�bw�<Z�j��B뫵\�\��hɱ�/usm�8!��p��jW�b��IΊ��F����]UƘ�(˪_#�?}��<���|w�#�]�)0�cL>(1q�s���ס~����� ������s� 	]��;��خ��LBJ����E������J~s΄ �f��m��31m��ͫ�Vx"��?~eM�s��W!��Wa`���zT���i�׈A��+ʈ��h��$�{J])��	��\�[�g��o����C_;d�P1b�cT!���}h��a���մς�*ے�uk8�6�7T}��ʻ�͵\�z)%��p����~]K��rErJ�N� Ï;|>��ۍ�[p:�P�u���X�)���\�dqѾ�S��U�(qX��{�[�K���u���g�
J��d!
l����,�/<��gGF�k!�W��QEB��{��Y:��e����Pع��_~�L���?�������׫�R�6��Mmj�m"@�6��Mmj��V�B���U�����8pUI,~Z���U��w��Ҿ�ZS6�;ryu)�=�L>����T�$���2l����m�6��r�A������q�M�������lݦr��š8.��d/e���a��{䄰j�l9�A����۬�H0�����L������Q��"ʹ�=�d����L-{��F���
ͬS5A�%�R���4�V=�.ry��!=�a}rs�&���> Fm�BbC�h��R�ְaQE�
��,D<���N>���Hػwj7E�Q����X��f����5ɮY���߼yM@v�j�@�N�T��O^�z%/^��Y����G��o 
� H%�m0 �h�a
��VJ1��(1�`J����탴�.$(�v>3b�V̪����� y���Xt�jϘ�����!��^'��h��7����!�lr�UL�jeü�f<�uy+������Z{��!ȴ�������,���x?��������g���qE���@�	D�s�C��а�ʪ�#z�c|)(�A��8�T� ��f^$$,��׃�[S@h��q� ?K7�A�Fp@6�sˇ�3l��hY2?o���T���<#H. B�q順�\i���
����^�y+!�)��d%殷.����'~~���l��Z��V��If�ư.����g X�o�yqy���{����w7.��D�r9[er6s?�ݠ�x���TCP
I��1�CLX$0HZ�E$�bS� S���Ndo,c �<���-�T%|��	J]a��y�@z���2��5{�`vz���*��ܹk���D���q7?="����/�ںq���j&�̭Ӈk��^�k7���>���d�vw@s]WԺœm4���}�Z�y0ʡ�%V�*�,ύ�,���7��	5��P[a��53Yj�vXCqޡu�Wϕ�r�A�J.��'Q�k�'3Y-d9[��m�^�ɘ݀�f �vr�?�	����������-�u���@�3ض1��%Q�9�q�_o�YwI��͑�c�=���H@	�^�$~��������Ϳ�'?p������ǁ*���x��j�JKO#7n�%�pN�����4�at>c�$���[+����2�A=��(UU��@
|Uv����cF	��g�S���F���>��!^���cRV/�Z�T˹���ڊm"�{���U`�;͓����X�C9 ��y�q��OQ�JZ��YcE4��3��C�"�5��y� t��.�x��<oe��L	�A�0(��e��oQ�P�ozL�:4����*�D�����~��{}���N������6��[G� �^u������q_l��g������N����J�$!WQ5��g��\~��W��ц� �}K��ܠ���YP� ����|������|�\�/~�������/����u��?}"�{���{g2��MmjS��o2��MmjS���j$���3- ���$�������}Y������B����|�����#����f���H�@�q�\3�$`���Q Ȋ�%�|��y���b�5ZU�� ���v�=�����#��Ǯ<Ʊ�ܭ՛y�B��\��0��"2@���JX�@) ��B� ��}#��2> �0���̤ J���j��s�C��r���Ǯ� :��7�@2s!�h7�u۬���G�Ջ��g���}~Fp��Q�W�m��>�Ƃ�6d���D�O�`M�\�vP�vn�>K��xE_K2s��T�}`0�( HpL ���\LZt
���MQ��xg���*�P��vE�? �D!Q�$�l��ϕ0�C�{A_���h5ǆ��U���	T4�	�4R�[Y__��P5�����S�z�+��P�$�� �$2������1��n���B *BJi�U���$A &v���A�����z�@�����\����Ҋs ,���!� >�C'i��8ˍ��-e��!A7Ύܘ%h�0�����V�s�'\4 |�r��|�bLm7{���e�/X�
bk��/A��dq�T1e���*�;�&
�B9`>K��rJAʌ�%b�����<�U�b$0*�����c~���TH����]
�HHډ*�`�/u��d٢'V��7<���Q��z<R�*�0/*������@рU�J,�lܜe.оrǻu�]H��T��=��},�n��n�qk��fyB�k�Up�>{ �vW~���p���V������ �]ߴO4��#���0_�ᚥ�,!=�	������=��k̪�A߁Z�u\o�����X��-	�t��x�qk��w�����9\l%��2����틯��ŵ��\6��^��A��ӡ80��6{�,�1�m�:L���4�f���ڍS��3S��߽��XK1�sO���M�����]�v�h������#��Wk�*d&����.��[�*/R%_4^�YHr��+F����/�KY�Ϲ�9a��z�u絓�,u�M�&�z)0�*~�~��߷��"#����<]���++Ƥ�؎h��4�B�I�~��}Op�N�I�K���l�� �Vl�a�l�A��#�[f���-η��0;#og��?>-���kd`�t��UA�?�a���Z��G�f���M˾=g6�8�p_�����lI�;�P2������㯅���%�PY�*�������H�#A��3�{6�@xU�E����R�{J�`�}��"��*�Ð�?@���A��u�yՇ�!UW�Ϗ	�g%�Y�Oh!���n�U����S&�+wOUU��`a`�t}���u�3��[��8�
�R�	* QD�2/�X��vM$X���k.�ɉ�evpϨ������[p��W{��y��b�̂{��4q�[3q����d��-�Ya���'��V��9{�<�{���w|�+��ͳ��g����o��{���X��|;w�>:>�Z�̑����g���pϼ_�O��O$��%y�٥LmjS������D�LmjS��Ծ�F��p��n$�*L�7э�b1g%�v����Ƞ��W6�Vö&�u��pm��&0�zI�^�� �N�������V��WrV������oPC��n���U��̃9q=n��2D�P�v���= ���m"��-���{y1˥+5�c�^�����D���ꇓ#�9�чJ�I�$BVH~��1��4�Y����M��� ���)2�h����	7�������Lr�XQ�>� �:#���.����[a�g�`�h�
�0P�� ���U �
�ۼbc�pW���,a��5�c�����t��x�R�'|�y�ɣ����V]��u 12����4��u!�|�._6��wG���Q�
��pca�*�0��ו��h�*J�P�B����!@�h����\a�0����j�~�V3@:��(��>��K�$]�ղ��q/N%�3�m�^���du*������/ܸ���$͏�  ��&}�Itus#Dx����Y�Vr�o,o9g0�R � ��~@��j� �� �)'�[�#���n�`�m�k�� ��Ƭ���Ȋ�=�PJ�b/=��
���� ��=�YAʊd5�^� a��*�ݼ���?���v$&���VA25ݼ�-	(�"�:��@n�r~��U�
m��"B�'�" 'I�P�>��YTi�tU�ݟX7͆k	���Zס(�h7�s��"G��ۇ�9�eyON��}_5�d�5  v_$B�B��eYP�BD�I��y�ν�7���G,���s������\%�d�@����"pn����#�|�)#*�(k�ah9'�<�9j>��9�ŝ;�<:�E������,�˾�a�ٱ�J�h�L�Vmmi�4�$n�QGp��&9�L��}�*A��8n��u�u��Y�:��b^�V� �~n�<z�Pnڗr��\���"��������R�3i�ڴwG�+5��A��w���x���#:�ɐ����N�^��I���ӹ����\�m��T��y�mw}�A�d�9H�Qq�Br���V�54j5ӂ*�G��D�;��x�
m�TACp����Z�Rʮ���`��־�v+/_~#��G�d�D"���\�%x��'�>�,��3R��#���:V`��L��Eܐ���#���{���O0��{�'C�=oa��%έ�sSá� z|����>�#%30�h�W�mH7\Ci�֡�u��$٫���v�؎K���FdYh
	�g���p���I��,���C�{�����_��iOX�[�P@ �{�y��}-x,Ȫ��@���<��x�@�wg\g�JP�S�Է�9 �𾕛P��@+�C��$�k��Bq�>:������%I8���_F�tw�5����������+^�[����ATc�a.�a�~節k�����|���cY:$<�Cӄ$����Ȁ*׍9��/` ��|4غ�~�g6�����%q��q�v�%��p}@�O���}�<�`�Ƴ4��1r5m:k�����Y����=G.�3B%��n�u�r�֑��sc[���{��u�֗uƢ�(�d�g���H�}�O�}�ײ8:��{grrv�=�ɱ[�gYJ�#���޹5pM5#�0fQ�8η�C9>~ ͡���ٽ�_2_�6��Mmj�s�� ��Ԧ6����[����یx��Z���q'���֘Tv���v�j1K�`��j9g596/Gns���C9;;�����X��N���B^=�F�񝂑�� �hUo ��[�`3qqN�q�Y�B�eذ�r�C���b�I
���Xu�n��XY/�j���-/���[d: l*r�6���{�Ӄ����sn.�e}p�~ �P�* ݻ%7��L 4�}������7�,B%'�Dc �۔",���Wjq���-6�JX���Vv�M�VA�~��nۊ������Vxߊ`R� s��@�p�q��f���M��xx����;W�s<��@���m��y�-����q@��V��R4��}�Z=�B���;��s"��F�c ��~�Ց� ��a������5B�G�ґX�bq�;��!�3�- 
 ���R�C ��3�D,�^�g3ڮ���'o���s~��dk�CY���.���'�� a�����<��� @�#RE�G��꫾i�����d���uUņ����h�j�kD�!P7��YYɾչ�IX�� g�0_}�,ϱ��-A$q}��_��W��_R�k�2 n��c�/4 ��>��K����@���yv�U�+:����&qJpQ�֡[B]���_�a� �O�^y�d�&*�:�/�=�@�Ϭ�h�fsK4���fq���z�� ������k(���P J ��r%���č��E&<}(o?<s����n�����A���?��mm�e1Dd�e��m� �2��ըEW��,����q�Vƣ�h
���N"�Kk�R�TT`�}x5�Df4�����E�X�zM�_�1���!�H�J�YF�e��:�YR�t!?z뱬����o���Z 	&��u�/9�S ���=YW�{֋���l��p�;I�-!C�6��7�s����ϕ�㽮P�/��V;<	��Ώ������=�@h*$���1�0��s��H��Aՙ��އ�c�V�G^as� i�y9�χC�/��q`k�hx7�@�J�Q�ҁ~�6M�/��2K,K ��>�Ưg>`~���?ױ�ٵ�m?�g�������p @
nUҘE~wC��y<APZ)���?�:b I@����5��D�*��GqtK��zs�s�:O�u<��NT�����s�����b�g�x���aN���`.�w�B���r0�Qߩ�&$��*L��$ֈҍ���RIǪ��q����^w[/i�P�ǿ���l�f�
��W�|F�rC-Qݽ���a�gB�^S��E$����S�bϹ�vs���(��X6�x>�,�㒈ϛ��W� �|�V��j�-��s�a�ߔ,:(�����^Y��@F�g#(+}��Z�v=	�Ϫ�z�aH�@�3�����M K(~pǷw�)W79>^��<���G���os� �x�٨��~qN�1qbo����|�Ï��?��\���m��x�6��MmjZm"@�6��Mmj�Ic�c�U��Rb%��vī�cY!�*	����r��]�H.Rۃ#�z��;����<t"l,��-}�����߱"��]�IE�!��76��ރ�����.�4��e.HU�q��1u��n>��F���m����z����Ʀ�6Ke!7W��@����rJ�\�v���y��H�pa�_�����&�����u(�ˣ>��ը�#�@7r?nP)��g6[І�dź���yf�Px�|�CV��Ѧ#R�������t��7J�`��vfyD����!�Lb�{��ݓ{�G�������v�j��}��lnέ_�69���A�$�xt>�wj{������^I�O5� p���Zd�c�2��������E�c�Z!�UҚmQ�� �-��H�ƍ1��QH���^ Ё��E�����Y��B<�/�}��|��kVKXi
+@�<6몐�ƍ�߼���d��OONd���n���hc��4Jn�f;����m�PgTE3 ��XU�3�ϯÖd-�RUM �D	4Xph�t�y$z���Պ
�4��a�
�$�Bd 0d�W}�p�+������.o^��"��.늤�<��I��[Ȗ�yZ�\ԕ*�Pk "���Q��$iV(���Ř�`k�X�Ё�����?������]��fw�
h���Ј�`�Gz����nMPcd��P�Q a���r�?�A�p��Z~Au��0�2������ҝ��,��ݓ���}y|2sﱗ ��-�"%1��΂�[ͩA�6l� �F���s���v���tڿ��Qr�k|@*���3"���u�Щ�$���X�XC�/n�${�Z�Z��J�:#���h�b-���+PB�$H`o�������z�r��F>|p���L��39��c�ػyw��B�YAQ&jUĿ��fj����k\���Zf<H̍��ᚣ��_�M$�`�����1��`��f�@�Wv%�ˬx��)�$OD����f ����D�&󙪙:�rq]�T���R`h�$&	$�{XK1�;�t�%���5׹pP`x��d��<Y�
�Q��>vF�v�
�s����%�݈Thl=�m�����i5<�>Ub$��o�C�}��W������a����\���mZ�Ց���ta�y����)T�z��j[�l����E�'�d8&~���pW�I������v��^��J��U	jξ����=ِ��Ex���L�X-I`ê�)k��scy���Y�O�+�og	^�j��լ�����q��kn�@��q���
��!��	,�B�J����V�0�[U�`m���Y�Pr~�^�r�t���[�`��/�R��g�ڭ�pOR�[^����5�y��>�b�ܣ�.�)j"��P��m�)�3�[���D�������C�놱o6z�q½�|6�r���/��F�fX�sy������?���{W�r�����z��(l ���L�
S9^��h����v����_��\_�q�[�jojS��Ԧ�g�&djS��Ԧ���0R�6���Q�68o?��o��i�f�͛7�\ņl9_�8��,����=$o`(?`�q��R^�x)�ۯ�ٗ_�~�g^�w��Ħiߖ���}x06������ٌ�;-����y� A�����P������f�����²!�Pdx3
B�jE��/���]NO�����>����CA�.���4�
d�Hp\�T�p�[��T>�� 9>>6�"�FH0�4�'8|y��@ZyXy@`pKۆq ������U��~P��c��a�P�y��戄�;_�͢�,)�0T�b�,�;U<q@����nIH���<�Jְ��l������W��T̸�j1&�P�'�C���
��Td�{*������儂	��cE,ªa�Qr�HV��,Q"@�*y �!�ǝ���f��)��[_}-E��+���M�<�e~t$���=�w]^�~E_�����tc�̍7��� ��
�46�ɼ"�Ge��w��C����М�)�~��R�I{��_O?���cz;\��l����k�pѫ�h���l1�Q)ϟ?����/�=���Nq0fδ�Q��ټ�$G:��vĊ����jV��(��6(fm���� ��o�q��U랃����m�g��vQ#y��$�,�z�L�ym�V�3C�^-	8� �Zk�-�&�Yv��9,��.�c����fs9�/ݺ;����&isCU�;����o?�{�v�xؕ�/
�/g$y]�*,"��	�*`:*�Y����)�`{����֑�UT�y�/k�-�͔~l�h!pO���Jr�gTљmQj$֨D�*]O��}�:�͚M�]Hh�/��$�T����6�r4?���H����_~��k�%���a��l�<�`Ym��I��2�"U!E>u��+Ա�c��@�zʭ��nK,f b�sS� ��Vp\a=��s*b�B��u��`2��.�s+WT4Vk�ǽcw��Gdb�\���J0̅�y\%]Ov(9�"����M�O7��������H?�<Q@5X;dt���qօ_��sB3"~<��OI��ʲmtm�]�X 1j�[��|=��d�����I)�������z.�_�$菩�<��;o7�%�I��b�ñ94{�[s9������ֲ߮i�	e�'��j��<F(A=�,�pX����:�g�z��[��g ���T����4���R%k����j����Al��}�c��Y0���P�BŲ��_|��[���r!�*J*
57f���;����x.�%����-XϠ��J�i�t���q��ۭ�s5?��x;=>�b�������XK���(vk���l2�'���Ǹ�G�Ja��i��{���Ԃx�_fv�*?��O��������ޥ�)s�pd����u�[�	��4�*w��d.�f��w��Ka���m���}jS��Ԧ�?e���MmjS��w��c�Mу�#��~(?�����������)�ps�a��Պ�> 3D<VP1����W�駟����嗿��\^\j51��QA����L�:!X�uZ��Z����GGǶQ�j�`�#�#�4�p�����A������b�r_3��;le}������-%B�+��񟿹��@ /��  //߰�� �$�T��kok
T�W5�s״"B�,j��f�8�3Z�T���T�ġ�`��$
��n�V�j�ߧ�uЙ��9���C��Z~�!���i�U+l}��`$��H+��rn���Xd)�!a�!���������0�����C��q2"�}Nm���C��
�@��;O`�$1@p�1� � �c8�z��PՉ@���}���6�A��d�`o��Ag��0�W��*� :НY-s��:���˓w��_��/	�������6��*�p�h�S��$�@�}��o佧����/$�Ϙ��ѿ�����*	Pi�����������w��H�
W"*����O鴯@*8]������:�87k	�DE@�@�@�	�j�už\̗_/ޜ˧�|"�/��%	��\GOu�5n�lv^;�g��QXMݿ��c`?���o�ެG����lu�5<"2raV��,Vqg�������3�@h̋=Σ~��G�� � ���K��ېͥ���5�m�w�w��e��G� �����p7�v�5��|�Z���Xǧ��\�rS;@FH�����~��&�Ӵ�G�,���M)�݊�Trx�d<�u%���q-@B������C���h���ot}�9~O3�ã<f>sy$!�R��n�ҹ3��Zҳ��z~*��>����:/�����]�1 ���Ih�d��;T�Z��R���(N����?���un@��sAbj2ǒt���v\�]_s��R�j6\�,G�5r�p�G����'@�]Y�:^S1�$p��؀VظA�{�95"�;���|t)��� �y���Ne��X��b��� ��N�km����}i:��
 ݒ6�5x�J�؁� *,�7���u:���m�iO���́@q����{����_��eb���,������ǳ�4�s�@�Jm�d�N�����z�o��r���q��1�"��L
�kc��>�q��?�R�R;P��q�l���M�7�s@�w~�Ӯǅ�K���W�t���z������I*ސN��p�
�7��dn��!�z��L�nDi��L�Y^I �p~T�S���2��S��(�u]�|
���ҡL�����T, �	6F�#�B*=�=W9umu��W����x��đ�������B|�uٽ���ݐ�l:"�Ρ��������?88UN�\Ii�-�b�6�2����մ/��t�u����3A�)�D�Y�y=�|���e�<��9�?Q �񶋘�k��sR^�,�{����ˋ��g���+�>����֡�!4���
���l̇���f-�!���ʙ7�g+O�c.���(@��g�m��1U��!u�ǭ�w��7� o���\ܹ���3�I=sw�0{������+t����vKX���c������f�\�:�j
��@�mhC��@��mhC�o���U�&���p���{�������(�<�E �Mg-p��/��W#�������Kݤ���[[!x��h�@�� u�q���N)����p8T! ��bc�Y����x�W������:�A�<y*�}��c#	�*���W�l6��N��lբB+�� .�(O�=6�y1��r�A�͑ph���i��ڃ3ni��Oe2�10�_��yvn�T�4�G�BԈ��� �Dh�ڮ+4�����i+���Y|�T�zM�c�6.�9���ߜՀ)��f����Z��R1�3a�)��?T�S��ȑP��.䚠���@�XA�>FudQ����a��=���K���2�ު�[Y.Rv�u�� 3�d��\���!R[Cd�"(f�$��}��j!�ɌÖX���q&��%��l~
�V6뽼���E05l!��%��\�]#�·˧O���;Y�A|$���o�X:��U��$�Ȯ-%J������D�W%xR�[zxR�,��\�e�����hm��*��d���3�v��'Z@J�^)%�,C��]��F�7Ium��:q��\����^�g֍Ĵi�"n���(:k4�^LV�cNwU�+����2<$��kh�aR�S�_��@U| ���5W;��7��TA�b�	%j7��@�6������3����}����u���U��� g^ȼ��I4��'39�²mC5N2Ѿ�Ff����2a��#a7�b$׊�]k��s>�T&�-0O��a���# B8wJq�-�/k��a��!�\+i��ݭ��-ȃʔw�b@%vϺ��B˺�����;u� ��:p\��f2�׌�	�t%��O�����k_�����/~)�t<�i�Y��@{q/Ya�C�Z�U,���`��dK!W�0SW�����8"S��Gp��0���@��x�x?�˘�c�\�����<J�9����[����9�o)�5��Jh�v�{5�r���e߰��+$(},J(ˀ?�����ª9�:Bͭ!/^�������~-�F�����B��3Eߢ����j�,��k���'��`���;vO�TaM0�+OKGCAI��8�����G��_+�k8�J�I�2���Q��8~�W��0���jAX�8���К$��}n�_�M����@�8��T�B�kڰ#@�i����P��~�r�`�T����޽���~U�F����E2���4���Y6M�B���V&f�%[Dխ��4�s���b���3�Ee2�3��쾚w��4��Yz��UZ�ڤ%9VŔ�#�
��\����uK��9V����yMk��?��%�p�g�y���9�y��1gT$���5�ʹ�Ӿ(}�
�(��"�?�/��Dח�_]���ȗ��2����X����Zn\���}z~z&��\�s.����ɏ~��꭯����j�"�J�6��mh��m @�6��mh��v��T���4��Xŀ0@��Ç�7�H���4�q ��t��?�ˀ���r���ǲэ�{������?��>���� 3�Ҽ��aD����l�lCx�h`|
�Ń(�d��8-��6���d���%+���%�,���5y�/P��Z�p߻wO��O�Ӈ�e�߸��VW���C��##�n� [���6���BH6����%����U*�����bTp���&*��D��& s����_w�PX #��V)��� 0��@s`}6�˯�:�t �����#�Đ]��� z�7� ��,d<��ޣz��l�r����&9�H	�9'�i��g���U�q�*j Ir��f~@��:�J�n>�1��.�*�l�bI �95�� jh����8n�zо�U������=v� �N� A�=sA��@f��D�?FuҶ�2@���
�2�{�'B�d���/S��[o��S��{�]ڎD����2fl��6���/7�����,�{��~�ɭ���&�痏��WR9��h2vVf����=�k�{<_�|Y�o�\�T��h�6���3cy��0$0�*�y�ê��|T��	���sA�����.'Ht@�1�[T�u�������S)�yU�T��g�)���Mgs��U�̇��h��������w�SU����[�K��3�ժ@�c�Ƶ5�(�.�x�������y)���y��
*Z�T66`k�U�X[t�z6�̹n�����G���ښ�`�ε��U��M�����|&Y���"�/~��Y�$����aG��+�]�q���������d�G�Ú����'Ȋ��gö��A� UW'�_��{Ё�m�\�wE�@��xm�n�GV]]�����hh�yE�:��-�"+�1��D9�Sӑ��3����^�.�|z*���_|�H�醶gs�bBz��,������D����,�̈-L�f�C�z����X'��=L�V|>�'@t4X���ik�x�Z�q]8Sok��7�ձ�<�	��,@�udYJ m@�S?0^y��>�$oOI5�#|����vy\���#�g<�h��u?J�ʍ6����,��B�cА���X5�'9��U? ��B�=��?�2�O����^�m=���OZK�l3�ε�*�J;F(!�m=�z��,�[{M��l��$|L]R�?�t~! ^���,��`\�Zf˩+��]�Ԉ nM�=�m1ǣ'K��e���F��F�CI%�e�8`Kc�$��86h�׺��S����L��H뎧#�����1T��N5�g�ƞ1�'����Ŵ´?Ƈ;B��9������O!�P6LQ�R[�<�5(���5�Y�a�����g�|���f+�펪�Z��L�˛k9�s��٩���=�s�6U x~�LgT&��w��жy�ȫ{��R�eW�̹S��T����l2�5 vv��0s'@5dE1�n����!/��∱>��{��r?���|y��dj]�l�$a�./�=m!7�+*=Pd%�t'�X~��~"��ڽ��_y{���uLM2��mhC��o2��mhC�����<�|Fa�@�v����sVu���?�����f�7�O�?���+����
�l����/��?��\]]�a���?e�*6kY�ɾ�Y��"˻����}ed�@@n���7Ӑ.��q�q�F�9�y ��秴�B�?]d3n�.n����C�6����OH�\�����0��1��Lvrw
� �z�>�Mc��? ���ͦIt�z��Fj$6�` �ؔ��ٍ,tܷ�e�5����� ��mm�w��2���J���T?���W��u䇁����є�2H~�Q�����B�3��� ^'�gH���u�iUa�����7k����6!>4�	�N��Gqd	y<�=!X1�2/�^�t��6hhG��� ���H5�@P���HQi��un!���3]%*�UM"�8U: +0��Ь�П���=P%��G��~S0�[�����:����$Z��=fX'��^~����k�<��/��X�xӾ�3xv'۰2B0��F�t��v���ZV�f��V�������j� ��>�ޯv����6��ґ#�&)	�x��`A����(9�B������_5I�C��+�U� s�sO`�V[0,�e�d��zcvu�`k@�5������F����a���IVY�6>m�2��J���Y��'�@��l�h�C�EA�*�01��Uv:_���q�1X�T�mon�OȵO��0���+wo�wnK�����J�|�ܚ��s=Ɇ��Ȯ	��٢�ղ�*�����}Pl�~�B��&b��ӠJ' U$B"c}y^��l|Z��K���H(�pD.>�!��1lϨ����1���\�z�HZ�	s>��"I�y���, �������$�c'����T�҈�L�{��c�S؞�����'�d="����$�@���*��(z�X��k��r��+��P�e��������s�ĕ�_���J�3Q�1>B>V��п���"-۵U�����r�{��{�2��S��R���������+��
���^h�@��J׌������#ľq�@����y{���:B��;#l���7�ZOh��K��D^���'A�ZЯg>˫�r��£�^���'����\������QA���q$p�b�]ˁ���)����j����+;���Eݚ��g�o�^9�v��UO����Rה���������C��>�f��Ӏ�7��Z�����g��YͿ�H(���r�6��k�(f�F��Zl\���Q�P}k�ù��]�p<ZAb�$����\t��P������1�:��J����Ț�s�����z_��g�L{W����"M*@b޻>��#�^���{X;ƺ�`����NY�4�B��^�Ͻ��7���-��o���)�N���~����[�e#*;�>~$���}y������W�s͓gt�^�hz�⎌���������2-
��v��0��6au�o����mhC��~��@�mhC��~c� ?t�#��S����1���@�r>?�[�hɀM%6[Ϟ<%uzkI�V77W���C��<��ε���u3[�FP	�����n&�{<��Ê���Q%��6_�IP6 �-g�������3� P"���
��u�Bv:_ps�A�{�/H�\�9�"�ox�_�����#����`d2��aS���H����V2�Cs�*Gg�1-Lr�N  l �K�/5`�b�M��܍�ʓ���\���*���ڰ�;M�����^�k�l`��
��B0�����c?�8Nu|vvƍ/2`P�M|�*G#*("����v�g�2YH:������Q\K�E
����t>��r�\�T���:.�YiY �p%/���A'3���x��"o����%�~O.��%QW�T���+��%,�V
��R��dd�Z��we�eu�&����${=��𓟐t�EEE	��x$3��?��'�������o���o&�O�Tn�>�k��m�k֗W����-A�:ù�����## ���X���2�u���f���K�.o�#87��o��
�Q��v6-����hǑ��A�r�34���A�I�2K�L����T��J_Z!\��r��ǳ1��/��6�N�ɖ�"���w�kX�F�D�,�;�:J�/�o�͚��jec��RIۄkT+En�����"v9�M]�;,�泙���:�R�FFI�Ǽ��dJe��յ���6G�²�t���x��}yvzNҡҵ���t}���/_�{&ӑ��BF�K��y_S�U����@⊊1^�}��Yqy�k����?:�5=�>p8����q|��|�Щl ,���(tj�hw(���[�!7�z̵�y�T>����;���@�.EYJ҃a���s��0Ȩ
�g��jx_�`-�Z�k��ޅ�z|����p�\��N2}����g7�)j�W̥֟7�߰̡�k�-N��V�� L�Ʃ��J#�+.-�
�a�KH�
To��M3� 	��a�@���am 9���#6��ZSMgS��+�e}I����81k,�$���Hט�8�Cq��~ۭ��n	k��ւ�����q�b�B/[�o��3B�{yPޯ�^]���5�G�{���hjs��ꎇv<��
~��ͣ���e�����؎�G��������~�� �_]�{eJҾB�qkg��վ�:���}�3�3]�v ��޲�/�}�⽋�
��W�[�港b��щÅB�
H
�?��ȱnW.c�g��ˑ<jx��U��3`w�q�%c?�_b�9J

�t����S*�1~{U{��z9��!��{xe	�p�q��okָb��6�s�p�H��ݵ���zE���{Y��98<�^
��P�b]s|K����	��xb��Y*���T�ْ6�X��n��0�11�g�-4Q\��Sj��b6�<fڴFB�b���+�� v։%>ѿA���	�!mjWz��󒷧�"#�*-Le6Y���$����^�7�|S�޽��\�m8���������������;<O�:;�}��5� �?o�o��Q]o�i��}��W�۶~���mhC��~'�@�mhC��~�m[2e�N&2��"d!���ZntC�����X�
�ą����Ź�\]����d!��B�OO	��t���m�ӏ?�珟��e��� zL
l�	<�F�.Cg��*>��������� ~ 6W��z_�)7�D�:2�u��#*�Ξ	Dȇ���F��(�PT/6�ظ��P��6VpB��@�� �'� ���C��ƱN��O�y�"�*w�Ȕ�g�R P����<��o�$3����Y������l3Z�Y�8�tVsW.'"$��*Z!������j�MEOyBbg�QKD�%(0��F�����}nc�?��U���#t��5��1-�x~�FefUwj��%�E%��+B������y��p�W��h ��}x�̈�A��g���3 }��aSG�������$��l��7^��^�V��C�������D�����|��gϮe����O�/������;Q 矻/��F%��Z�����fS`�����E��'~p�������Nd�x��@����^��MГ X�U������tDq��!��M����%��kN� נ-Ma��m2��gY��Ŀ������S��v�B �t�2��m�-�\�w^��LP�8����	����@.^]_w���a��z���	+�A��&]au.@M YTq��O�P{Y59��1����Y��J���T��iۭ9�Py�n�^_��H�1�'g��2Cq��@$&"��$I��ڦ!�EV@�Oק�0�}R��
�f�o i��IX�߇� �z�Y��3���q��fq�y��yE+�G΢��L�C�� I���� �H[r4+ǩ:�q��,Tr�s�����P�Y-�2�iP�˙��ӥ�z�\���u��6�@i\wyH���A%������T�Ԗ��W��/�Y�/ed9�e����.��Ql�XX_IX�%ީE���b�#�.Y}^��ϨIj�����$ �1�����Xis�$ H1~���P,��eO�=*���
~ ��t�����s��<ח�HJ����}��+?K	�W?x���+��ŕ����_~M�?^V����z�G0� ��6(t
9Sڵ�ߞp�E�yFĠ�`v2�]P 0n}�����3��|��k�?r=�,���%�y(�����L�����}9w%p�=/��,uM����������3����*��PM��h���m�����tǉq��u�Z�����������
^cV�a��6����b�L��-D���8^@�u���F¼Ĩ�gW���m���!�"����g�x�c��S����}1&P�3��	�z�i��7%��[(����0��)w��ꀂ���������ͱ���:�Y�j6��� ��L�e<��w�:�=[�>.�����W���,Ӊ�&w�d�'QJ+Ec�9�i���	�4׏���R�͕ު62��mhC��h2��mhC���D�p[����즭�8s�	+��l�[Y�Rr��g���+_���^��Հ��'�0���\]�v�������;�WrC�,��W�^2���ȵ�@��>�� �q3�c�VHe�g�ps��+���o�)	����52F���x ��7��"ȻJGzV�fcP�[�XN�3N���[�% ����f����Voa�d�c_��a^�ش�#B �Q�-�����,X�.��$�����yk��A4V`�l,����fT/Z��B�d�=V"HM��g����	c�~�3=I�u�e1�1�۱�"*�,+;��6b���W����eIE?mT;��ʜr"V�Zդ� P��vw�5�8�ug	�$N\xu�8%�a0 M��a5)* Ԉa3�҇ZQhA� 
�0�� w1�	#�-hֹ3��M�5�j��Y�H< ����%-*ʝ��W[Y]�i�2�������߬�����7�$ay���^�%/7;���!�cč>%`��w�Te�8{�q�f.%�~&Xȴ�"°
iI�����A�#x��Kz�{p��10ժ�A�`�t��[�C���j�8w Ml�":.$w��q�]�Ϻ�j}��\�@~0�D,��1�� jY���<�
}��T���{0�h�p�Ԋ����^a��&�9R1!�6���)�C� �I��ߢ*x�^ɮ(��@u4�y��g����{��9�8��㑞�J�O��n�d1I%KZ�9B�j7K�@@5�|�&l	��<��?"���&�B��2;�����v�,i�D
����V�:T?0"���]9���lC�[���T� U� 1����oT�T6KR6p�ly^��$Lb�*�q_��	H�ş��Ŗ+1�`�s6�"�����z�\���.X�剾u�st�=0��7�����_f���8O�~�Fz���i��� b@�^��T#�����"NCa�Ȧ��.��IH�t3��cQ!�W�J��8E�y � h9-������R�j�*	(��
��JT���*�X0�"p6^Ǭ
��1�Â�_��+*x_s�qBA��t�#����o��n�`|���+F^��J��ȕ��a�SR��#�#-���A�Y
�P8����>���*�9�m����t$�q���$���{�Ȧ>�a=��H1�d�ꠘd���ǚ�a�~�}X׼���	���#@�[_�+=r_ �a���Z˳'��6mr�y|4�=i�&T�sK��e�/T�/�\���V�[fI����5NQҿ��ۂ*�ـBQR�g[{3�W�I2������U+ܵ��"H;r�e��0Smɬ-�5�����Ƽ^�B%0]�yZ�h����
	�s���lּ����5��̼��W���zTRr<����5G�(�����q���\���c�@�;�����������3>�b��Z����/�|򐪎�d�{$�S�#�}s%�X���ú��6���Rm��������R�4��>��mh�#m @�6��mh����14�;wn��W^a��.?0�^���4��999�/|��o|C~��ߒ�������ц��z��������_���37�	�����HMW��<��fݪ-�Ζ�oX�Ŭ~��X�H�X�z˰r���s���*/i� @�������ĳB�@eA	y(���,�����9�''<��"g� ��=\:K`8���#�$��Ђ:�ݬ��I=_D�s ,�W>J}5��"�L��W�U���Zu�U��W��k<�a�޺	5k�6  6˰��u~.�="�ٮu\�4��oU��՚��)<�bd���M�U���z�:ql���	{(�1�Y�o��c�m�B|A}+���~�ˏA@u E�#u���e�u�� X
��#�|�g�V�����d�1� ��ц�ܤ��M�ڙ/�r��t@&�)UR��h)���9�>�¶���ky�/�+�>}(O"����Ʒ�-��L�m(On
�Mļ��V(�EY�M��㋡� .S��jT��W?����#�g��P�=�Νu[��դn���?��jfo�EN��dH��h�9p ��k�� K*�y��b��0��A���dPnŘ�J-�PmTb�\�����$[G��O�����> �GK#�w��@�;*�" �担)H�A ^��Ֆ�S���E��~�M��J�Z���K*��u#s}�k��ʷ2Fu-�uJ�� (�bm�*�1��b|6NYA���Sv�q�MY��K3� �E=�@_:v	)���G9	�r�y�3ty X��{#D$С�u�y�#���[����\@j�7�h�ViD�&M�
�B�a���i�.{��Yڏ�l"����zǪ�3�w�vqKV�ZZ=�q����e��+Z�Hr�%[e�+�ت�]z��o��x���k����U�S���q�v�2��"�y}��\"q �y7�P�-썘��@~�Tp��5����Sb�c۸@�Ɣ� رV�v�B����!o�d��J�z�gF���8���uk��WM�ɉ�=�ļ�����y�':�s��v{^����5������*���yk._h����˭y�Lo����R�,����=���@T#�rT��$�,��#r�</]�RJ����sj�8�-�U�G���cl��&q����+o������l���N�2{�}-N��ϣ�I�Il|�@8�
g����ӈ#�}�=�j��,9��蛑�!o���:�^�]�A�ɇ��u���_�1��4���*�ƣ �X�_��أ��YHξ��;M��{��6g��*�),|ޜY�y2��kk�,��_�5V��#G���!�}�7[<mȹZ�\S��g�4��?Z(��1�?f�E��v�!�cb��#2���p)�5���l��!�xj:%T�x��u%���/��a�����咤�uvf��\AF��D��*9�u2Bۨi<lhC��~Gڰ�mhC��~���+w��'��Ã��7ސ?����ry������=����Ky��97Y_z�m��?�#�Cm�
 g��b�T1��}�[���ݓg���o�`wZ�R�4ے�dF˧�a�!�3<�A\ղ1|���]TÚJ�*0��N�z}��~K�fKO3�~�5�0� L ��A�;-� 2[q^� L{n��^U�m�C� �6�˓7���g��0����Ӂ����o4��9Oxny�w������^`���7�H\��8p�li<8�m�yM�e{�u�r���� �a�B�gW�>������Tf��|�|B���z��w%��}�7���H��#8D�"�5�ΎA��Q4�6۳-+�	�D��>����qs�#�lH	 ���a��x�v�>g
�F�U��2  @��	h��]d����®+�����kv(}n��sVz$1�]T��v��d�'f��1����>�����*g���.���=����x>�l.��R|�+�fSY�-��
��aŽt_ g�����2+BGF�����|�����8�\�Xe�#��~���;�r@~Gr�5 GEYq~�&�-?��S �V�J:�]�+ ��:��	���V0��G�:*�#t`�A����ʐgtb�5F�:��lN�4#`����|iZ�T���$����xX�U��>J�?��ZKLu[��x�ˁ���_�B:w��X�lʹ����@��� x[甅��
�V���D��g$A�\�}�����z�V���M����k�zݔ Q�m���J��'[��?��Z���cާt9C*N��P�兰��;�D�@䴱J��*<S�6��XH~���1�`�cP�FZ�����XS#@�m���B8jer:��jO{��h,'�H�N�#�?L�������-��ZɣǏ���s3��"��g���������� ����j��^��]C���s�{`�sѲ�R��8�%֘���ҿIb��<Ϝ�˪�m�@Rt����ง��&0�q��v�i\6�����Q�n tz��x>FL����X�{O^�m��x]�K�� �%����g����q �~9���Mg��E�{�	�q�W�Pʸ~����rĉ��$����e2��!���X�0v��Է6rBSJ�x��ruO�y2��=y*��Jp�B�����ء���
����PŎt������=F�T$���E(/�h���s�JOT#�z���ґEM`�Iq��C>{jE	_",�󼊵#E��0����<��{�����R\��Ȕn�"�%��1�W�G�,d�ێ���H���j$U� @��}�#��S�Ҫș�k�ڽj(���KS����j�๯u*M�`��f�?���	��̩�1��8^����.�ǘW'�[����%�5U��J�	x���<xFy��|����o~]�nߑ=�^�c����Y|�#����u��-��Ս�����OFK]_�l�!�L�E�gz�8�]��dhC�І�;�dhC�І�iI�EC����=�7���,��������?�M�/��|)���&�'��Aفn�sZ�Z�̀'� ������}]��_�~ �|�1�%¨"^%d�$�U�@:�v���Շ>��+FY��cW�֊W�2v���\<���Au����Ū�P�X�~���F��w���$Md���`n��[���#Z|���F��� ��A���h��`iZG,� `�
��0MG<���sE��< <��j�+h,�)�����Ǐ��U��j� �3�0�ЮkİMq��D�	�G�-�Y�xU�� �����Zd�P-�l5�u9�4P��������X;y�{~�� [_i	�#  ;
�b�c=葄�G�u@�p1�峹��H�m�占j{>_���-	�*@�z}�Lf�!��ՠw|ʺpS�e��Z0�2 �{��X�U/����P�"�=�T����7ߔ��D�iƬ���L��c� Ұ�13���ڲb=~����#��`U�
���p�sG��*[����i�w�� F��D����#��h��0yTG;V+M��I�:�2�\ep��P	 ��.�G�+�r!�Jj|6�;3¨�o�c1;���� ���`\�t@FB���i�G�7���}K�yW�ٷ����������5ձB����F������~�����B����\��<��@���Q�[/�U��f���Hx�̙� ��	2
9�|�F>�Wn��5ŃiU����J{�'�>�UL#,��F��F�t�Vh�	rb�oS�?ɑD��] R� �z?�������_a<�fS���J��Ȓ�)%j�J�,���HIg�'z�:O�������x�țit\/�S�$ f,= 2�� �	LB�� <&�o��="1�ךJ����Ȃ�#��B��Z�~�¸Q&6^v��JB���	�}���01R`z��͕l�W5�B�c�	hL�L���vRSL���V܀~L���Ɉ�$�W
�C�KZ�A?l���<�M�n��~��&�b�)L����Կ��j1��q�-�Ac����N���������m2�� ��wG���Fu�rb��  '�爎��*JJSh�Б���kG����"���*A�x��x��^b�b�l�� ��\F��׶���G0x��=�<���j���V�9�u*Ӯy'K[d�[�}%S۩X���f��;��k��;������Ĩ6	8�=���#��	�B5�c�s �{Y��ƈ�������y/��ilJ�/[]���m�SSj� ��c��i��X�PU����7��o�}�)1<!�W@y��!?���!q�g�Κ�I�td�/�
W�K�s6��o������C*�����F�@q��o[��/���B~��/}�1�c��%w����σc}>�{��:[�3�N�={=z�h��ז_z�;�˳�a�,ehC�І�;�dhC�І�ig�3y��SV�~�_��bA@���������f:�z2[���\'�13`�G���z���2�� �����^{��������H�O'r ����X8#�P��>�����Y�Y.$��Ͷ�B ��h�m@��Ī\�ʅ`��oH hR"���������lYE��� ~�P��	hM���>�!�.Q݆�+��D%�eF��c���"&-Se_��$a��3�Q�@�� 6�f;���$�B�_n�F:�@���R!��
p4TyBM#��Pw� �� Ӏ�e��Fl�.D?C^,o������������'C�����1-J��W_ �	�DJr�]%��}����
�}�	��=q�Z1}�	�rq��~:�2��+�7T�`���@�,���jN�[p�Iޒi�x*Yy@�4NI �=NN'����AI��4Wz8{b��J*Ŧ��������\.�気���U�Kc9�y�J�m0��b%�^Ͻ��qk�-P ��na�Qñ]�>�s����t��0Ղޫ���M�]����+�`�����լT��ۼ�*�)v`ٿ������O ��W*��,a\����%�ގdA�I7��:~��k���o��ݞt�a�:�y��j���NH��������߫�I��x.��w���v�\�C�Be�7�#3�"���Uf��Ծ�*Y�IvA �N�<��F&�>�^�'�߻+g�. f����xI#	�����DEl�*����ozxѣ;r��"B7��֪ȱ��T��%ω6?ȗ(J��p~�8e |I ��Q�C g1GR�P�
�I��{T�;-�p�����i��
e��P���x�Ce	�d�\�G�:OQy0W�'U`�u/��4Q��l��2��d��������+��\B�L$�뾛����\�1�긑}^xgNe��e�Y�(�qA6�ʊ�Emvq�� ��/R����=�:��?Y�$p��l�D��N� �G�9*��N!A�3!� |�s�䘩 ���� �}�D�	�>Y����C[��y,:#�k2�S,8�b��0�^�-���w�U}U�������ͣ-�/���(�H�{���2t��C��y�	�˞u�9�\FIXb����Ѯ�`�̑в��z�:�!�㜌g�� ���O0֩*L9���cNG󣪢6�U�ι\�m�<I��j�1�gF|�]W	�e-�����t��`��IL�^o'�S��t����1��#�g��'������č;;LN#��`����T�Y�IБ�V�����/PpR:��쫐�e�3�G��Z��SY�q.$��*��(b�L��8J3���2�cܷ�L9�uk��x\���,W�:̣��Ύ�s��Ȋ�p��2#<a5(��e�D��J��l钝x,|�fΉ�(����ѣO�G?��>�dyqε_�����ݧ�	J��b��|~v��|��/(�z�K_�{�n#�G>����g���
s=�����������������oޓ�mhC�ou��mhC�o�!��tyK^y��J!-I .`ӌJ���3~�^����`c��{��~�}���e:?���)$�{���rq~�0<g�{n�f��?�F���-<� ��h��7ݭ�ܮ��5�V�E��m�s�:ud@�./����-%��[��������T' �P�p�T7o�?g�l�`�5���  ]X=8O������T���]nClYq��e��zl=h[��J����1���YY�r�j��j�f�_ц«C|C�E�?0N�N̂EM�P ��#�,1o~v�wH����6�;�!1R�ш������b�- �����lZ�9������t���ZW1��#6��B ]
��V)��w ����<l\���v0>_�j:�����3I<�u,��_�k"S�-���^�2`��q��'#��x�N���&���rv~����'cye]�f�Ѿ���u-�˗��-pW!����y���Ou����=I39�/h�TA��v���,�p>^=��f�zL�6`(K���Z����8���\�U��U��n�,����2"Kl-afH��V�9,aJ�jL3h̆XvT#�<��
�X�y����sP���t-���h׺��Z:��#���C�Z��2tV0��/�H%�9O��֬� zb���^���k @�(6�O�k��u��lg#���!��^�w*�t���I������j�pm�z��D�,���L�����4��4���ʎ�@+�XG��\�I�����B�mE"�q )��D�q�ϭ�ݏ,��c�2��TiQ���A�[=o!��r�Z&�H�:ڻ�H*�@Ę�Ŗ�;��l���g��e3["
d1��#���1�o$��P��Iv�ȭ���9�~�8���g�V[Y��e(�͖�4��S�^3�^E�ײ�k	�2|֒�#�����DQJ �kXd��������1��������\���n�'c�˂2,�놶6��ܭ�%�����zN����H�6��}$%��Q��p*q츟�b�C�2 ��))43t^�ג��C$/��{%��O��ߞ��v^}%H���\q����J�τ���똁�H�C���X�Rn�p���<aƘ�mF���Il6+������狄n�y)��$|`�e�s~�mЩ=�bXgG���.�6�u܌f������r�4�w�|�@����@�Q(�\r�`a��1$��kWp��0���D���³�:�p�v9Q;�B�I�;�1X`�*��Y�HL��V��TK:r�[4v���0�������\��5�{[4�@Q9��g�{^e}���ˡq�=Aq��A��{�p'#����y��_U7~A��Q�g��+D��n�x_�ܺu[NO�x�ϯ��z�X�s�'fI�ߡ Co�g�Y���@�.<�!,�e��9��]`6������B����>��O?���7T�|�ߔ���hj���w�\�׾�y��F��3��K_��G�~�9��/��0��(��?������2ӽ�B�-'m�+��mhC�o}��mhCگ����k�_��?׍�-���g�����C��)T
[ɫ�n�s��״$�ϧ�\��s��$��3�?���M���XM�խ۷���_���ߒ��?��ƪ�tӖ$�Q#����ڬ䵦!yQ;p_�����>�s�=�+`���~�����X�2����}T���;V��Z�_l�u��|���x��!�+� �����x�y�����M�'�IC=�
s*2='D� gɄ�#��J�����-�	Fݬ�X%��,4P�iU֬R������Āf� x	؀�y�F������4/j��I�[�,s�; �+R�$�hY�J�����Y2"�G#�A��y�~>�*��}�AzL(����^'ذ�ь@�a{  E� 6z�n�����N�#�]�L7�PecS�0�}2�l��� H ��q�I�P�p��5�ƴ� �0�S�d#	>��;HP���{����X[���^te���v+�lt��l�6��)q�ݮ2�9(�%	�Eŭ�iڷ󳹄�Z���W�znS�����=���{G�Z�	�}�k�?{�]��C��O��?�/}�^OT��V5+�SV��%}p"+�	%��5�B� ���gW���ɼl<bu/�C���$�l8�B\ڶ�} ��ס��̰S��9�7z}i���� �V�A�`���@�+�]X;��ʇj��pC�*��`�+�z�l=̒���~ Xe���i�u��ϼ�"LD~B^aޛ�EL��	��P������v���*�FU�G&��f'愕ݨ�G~�l&����z+�Mn������1� s[מ��N��r!���K N�hd�\\��9�&��ݹ\�֔ �f�P�BG.զ���N _Wܲ�]_?q�%t 尮�u=@E1�T��3�� ~�J��j���"�5;Z�ڧ�O���P���S�s*��%^��.2�� �bEgA�%%.K�e���z�0�2Xt�kN����������4�D4Q�)�璭y�|+��ǭ�L���\�<}�H�g�z�
yr�X�uA;�W��ڮ�Ï�'���B<��aA�ͬ�@lb��t,��M���X/��i�W�[�u�z/�B��Pg �VG�]A�8
ݚ��9AYP�c���ђ��W ��'��1�� 8@�l�T��>o�-w�ix���^�1,a�2c)ҵ���N-��l#;1���2=��2�H~ta��U���m��`�vN�OrDIY�Ni!ϴ�t6]����C�-����N�Ȝ��2;0�.�:x�\Iu�Ѵ������#l#C�XAi��;����(U4�h�թ5P����+���G�Z�H�Hג�liW�2�}5>�+q�qݤZ������Ն��-�Fd�=�HA#Y����oh�Ĭ��2d��B^K��D's�阈Q �T�̆I��ZNI���� \WZj��d��!�j�l�"�/�ǆ�6"}e��(#A}$L@����H*�L��k3��f#>k�`�Ƴ
H1��0н6kS�;q.5֜�J��QjV�$}Q@ؑ�SD�����i�v�����A���[}6Ba�d&ǻͭ�(��|�]6�r�X�㧟�3i�e���j��#	���<�H3��R)ٜ:���~2xp�s��ǲn6$w��gO����Z(ܙ/O�������+]�拥\ܾ��>d���?��}���m}�aΜ��>��{�=�<�����D�z���N�vB�І6�߅6,�C�І6��H�/��?����w��c�J���g ���p��:Y�Fw��g���&m�^���������w���D�?*O�>�۷oI����� �����T���|��*-�կ�9X��g L}&��7�u�q;��cSF���@}2[�F���q�L	�*7Xsma�Ҙ>�s �(ƱbS}uy�Mq3���C7�9�bi���BŸ��5�^:  �e��Z�+4���;�v�؅Ɇ��u�<�q�n"����ُ�z�Ĳ�Ւa�b��g5�i	��r=�W|J� �S������,��X�ru�\���ήxT=&� ��v 9 ´t�VQ�\԰n	s�? ����稸u�� j���r��X�	�!^Z^�Q�PN��.t�w��'��[�LS ϐ2H.���L��|M��BC��:)��8�ס��ر�?�s��,;�l��nS |@�A(*���r
N�g:�3Y�w���g+Y?��G�S�.V�	r�=Ԓ���۽<y�\��o�g}����7p��^���`��8k��Y�6<n';��cɁ�� ������G�RU��pJ��Ug�'�>�U�O�.�h���V��v�'�e��͑������8�TH�}���T������Z1$dH��EI�X��r*�B��[��xF#Z4��3���$W-	�,�*��{��IH��গ�!�BP�~��i�ʩ�%��������F׮=�Y��u�Q	�������;�����u���?Q��P�+�
}���$ �Ԓő#�(]���c��N��t�,����W��_����Z��q�Jj�o�;Z�R�ɍ���[ԥ���C9�z褓��1��y�����o੏�������ȃy)��(������xAmj��BS��g��!�T�K�m�:粀�e���:6���?�����m7;3s�����ܓg��ѓ'z�V.+
U���\�q�@��<�56�Ӯh���tG�5��P�x=߂�ֻ�Sc�.��h3�:[����s(u
�K�1o;T�='r�=�q��u,�z�T���̢'12�<о
�6UZ?���ϲ��<�k�c�K���JO�xu�Ϡ�-�M??�A�pt��Tn��0�)�*������]�{?߄��^w}��������@���N�<�b�T�@ƴ���7�U�j�EU>��W�u�	B�wv[�9��t��БOq�t�I��l���m���c��W^�Z�`G~��`�븽����:��,����VB���y+,?&^�]��[+�8��rCZ^ghHhjĺr$W�y����
C���ϙ'� (>��H^�s����E!s����z&�=����7�4���Γ�h��F��w$��rD_�:����89������lt�疅6�L��G�CJ���}�YqzO)I,�tlC��1��ۀ�j��6���^F$@h�������h-����<~�X���r~qK�����gCMS�]�
�ۧgs�{�-d��ή����������aX����mhC��~��@�mhC��~c�_��?��U-�JF2`�R�].�2gv�!���-~�>A]�`0���jK`�*2+�ql�!3`Q��cX>�Ag��4T,��<�[�rC2�� �ӹnO�/�uK�,�ܲ �T	��Y�66�m�%0T1H3�*CQŎ=��������j�� v7��+�F�a5k�c���<���n�`q�.,<�8�p�/KG���F�BnT*��j-p�U�QH������J�����Z��:�1.t��$��%QiߌuӚx����n�W�w������Lh��c�Wl��J ܁2TwL�Vq��9���<�Y@�
�`k9 �8r�!��(꬚�*e�8�E۔�w����{������B�՛a� ��4�H�W�i��l�~�>L<���%��MX�;�B/�V2Y����b�}�A.f{	�3�?y&�|��<{~#�M!��]�	�ׇ����?}�P�y��)�������|A�&��ˠ#�|%��Ո
�>��>���L�ڝ;���=�o<��2n`3��ƽ]qa䑻F� ����@n ���\C�6�g�c f �j�����zo��j#�H�R��
mkF�20���f��ga\3�lx��^���؜G~T�2M�d&B�Sy���)3RR�W_9��F��߀��?��p�H��H.���B�m�sj��O�c9��d���Z��F,��E�� z՝%֍�:�Y�T0�]��0oK���z#bsW�c��qڐ��-?�⍅,�7|`y�9���E03�vp]��%mz*TfS���鄪~-��)DZw�Ad9'do+����!bD�(m�@F�t-�n�f3Y�]^�C�ms]��J��r	��3�'r��md>�x�Ww�O:PrTC��~�-���L)B�, �3��Hl��*�p �� �˳���!� ��C�=�a!��{p?M��^%��C'c�`�W���B�\��b����Uv@Gǋ���������־��|����\0�'E���Oz��7���},Z�:`�[b�c$��^��+*A��;O��������w��q�L`���,�f��m�����^<
9���^A���+�� ��Rk���I���+L��t��W�0	��2b�.;Ů��,#
[>�y""4�*t�i>
8���Ik_bJ:^���VbA���D~���Of���0<���2ўQ#)��P�Cu|�2]K��`~�N�H[Mfw��x8���#�&����j#�qJP�@M=}���
���\��7Ҕ�]?���/��{��>�mH:�ކ����vxPV/����J*�&�̍��n�(3�əw�S�z��޳���?��ܬ�r�������_���ߺ#q2��y�=P�[����<�㽹���z���[����AX�2��mh�m @�6��mh���Z�P��*���5�9��Q�J��a�$32$r kM ��1=�M)�Pel�)?*	Pb��X����}�1���A��oZN=yv����m*[!p�C-z�W���H�����\�x�*P��{e�C {�U�e[���!���?��єUr$�t���j�jI�˚�l��hƍ*�,�غ
Jy}MxUzr���=�^�x����]d�)Y!uՓ@6�  =ʹ�҈�	�L�zf�c�,��>^'v U�ˀ�������X���gK)�ךv�'#�3&T�D��-<.d��\�����uIR ���Zy�(�6�D���kG�6�ׅ�Lل��1�r2F���y<���O�Pm�lgf��*�A�!��B�r��w��D�ܹ-w���@@��f�|*���T����9���q}������7赱�rŬ��mڄc��c���ƿ#F<��4�=���R�c��@"G\H�nG.�؃N�O�$�Ъie�,��A_
�- �����1���:?~Z�+�`��;�VW-��Mk�d�jw�G?%�b8qc�����jkb�<Ĺ�0��KP! �=���l��r��G��k�[1��f���Gm" ?[�������Y�ɴ	eZ����l%Z�<��O��X}U,��z���&/���Tf�K���yR�Z�.ƺ�v$-��+�و�!X����Pj5&�UU�i���|
�u����,���8���ܧU�1e�����i���Pp<U{��$��RfB�_vo�y,ނ͈��l�Z�J�j��5ilkAY�e]����:w��Bn_o��wߗ�o�k}coe�%fE���V1ׅW_y�c�񣧲EfHe�)�������rQg����K^	N���h�/	c�B(�pOC���ۘ�Ӄ� y	��8����hw��B½�6r4�����_m�r,��
H`�'�T�xl/d7������7��
o��3�Wx��?�e�b��#=��aG�˹#�m��ת��||��ߣq�n�N���������=�Ub��9�#�h��I?$�����:�SĀ���i���X0R�v�g]^��	�Б>[� }c�H�x�M�8DO�3WڞbǙ:[�Qf��ì3R������{�=�
���?�R}�4�����]��g���Z38E�I�&��u�eO5/=3���i�'�c_���aL'\K��s�DP��N5\�g��>KU�Fve���.3ct|�yOz�L�ڔ�7��4�%�������V�����ǴJE� ��x�,�k.��VS�����Z��j�]?*�J#0�r+���w��(���E�δz�.��z�#I�3y�����ܽW�l�1��((�S����fe�W���G��F��?��?���T�6��mh�;m @�6��mh����~$�Tn�駝�� �ͪ�zO@)Err��/��%y��_H�{�������00�d��$�Ec0u:�@���E��O���@ �O>~HK��O/eqr�틀U���R�(�&���������;Yݬ	���OT�~��T���t<��`�L�]e�S�$ZUew�o����1�x?��756��<��>�����Cq���8��PXt��U�����X#,���J��a��l������<A��Ā�3���T'�����T�J�@#�Z�Q�8P�+����k�;�h�~xO�G;�Ȭ*�y�zvae������Y�F =0��n���� �ւ�Ap����?�" ��
QK�&�%U�O��?Gտ�Ok����'��+Ni�e����<���F�w��ɭ�S�grz2�qz#�q��۪��r܌ӄ����}��<Y.x]��9����H�C��2�v@=��@��jɫ;<0T��"��[:k��ɒ�٤ 0���|G�.	��UAP~���!�7�%ٲΙ��I
^SV�-=|���8A��#�W���E���;U�^��l�kZ�ƫ@p���Xi|� ���L.�z� |��J� H���I^�,.9�-��
�F�#<������X�ZT�C�-��qf���F��n+�v-M��K�GevW��D���7�"/�
�Ȁ�Hںނ.�B�64��k�~@/9�Q����14���$��G��#wFX/<)��q�uQ)i��/ 4��d;��WN�jϠs*C��r#�$�X���+��	�-�D�HCS<q!n��Ň*���8�|��<<_N������<�l�gFB��Y �n/�t+aZ�zU���9�9wn���������96��y��]i6gNM��1O ,�S�al�:�f���Y;m.J!�=,|<$AF2F''Ԇ(4��vr̦80�*Ȉ ������°X9�O�: {8䦄���g��\}��y��>`M��3�~���ĆWLxd2�9Zfٚf�k����{c�>u��ǀ�Ʃ-���r�����k�\{����'z<0�϶���S��������*�z�޷��X���5�/��
8����{,���V`h,(���֘Mˢ����>��&p���+�|�x>2U����bx�[��5�� ��Hm~�����g��S��wc�S�f�MX�G��z;���;�uDP�FTHp��N��`a��Z�
���/���s�d��5��0�� �L�3�\=z,9�?���2�n�e锕\>Ϻ��>C��[ޓ̲,��l��Ќ�QV��6����j�D�>�%�g�=k���=4$Up��јc
(�gcqm��@����~����'�~U��|Ku0
�P�5�mm���F���Ս��2;ȏ�mhC�]k2��mhC�����1����ῗ?���k�w�,j��޽{���
����Cx1��o���ߑ�f%Ϟ^��5�L�y��h��HT��2ɠ!(f�c �V�n�9S D�Ɓ�<�: ă�߱������G1���������L�}��ܺ8#V��Y�h���Sy���紮@\c��q�b��ݔǁ*:�_Z�ۆY  �bg�a�T��QwՊ���#����	�~����N��L�QV�	���}�Ё&h7����e�/�e��,� pT]��y@�������UB�w�\�̸a'x��u���a���T�3:2K|�m��ƱR)�����asXj��^�� )�ު.}?�e�L&��< ���K �V�1k�{��@��AϮ
�i��Zg�ǌ �m4J �`hsDˎБw!C֡�2�Th�^`�,v1sV�Z��#����GfE,mO`��$icl�e4�%��TH@��)��f�w��\��8!���ʏ~�c����^c�Y��I3�[ �����T����d�B�u�F�CлPߑUK�7	U�{�����{����hID���`w��@�~�j+�B����!7;-ګب���ǜ(ڂ����SJy�(f� ���8F�Q�� z�t��Eu���,1 ��7t oh�(?&�y�g	@(�@�nV�7{o���u%����}��z�� ���e�	�
K��/�w!Ex&�jR�!�fH�$�n���o��7�[U���'R������o���Ue��$�@�"�w���
���Zc%>�Z3�K6Id
;#>��~�m!K?��R��[3��SC��V��F�ͳ?�t�f{��	����	�ֵT}p�@EP��~��(��\w��QlʼV�z`V�*w�HE_y���H�A�qgW��&������ �G�������gk�/%�:Ĳ�����!�7M83?�Ū�	�kU5�=���NV�k�良���ݓc�r���N� ��j-5\��/�j���;�w̟S�PU�q����Mػ�$$d��VvX���^�b��3ZLAQ%��=\�]���*������6UOY��	J<�3f�����q�ԉX�Q�Z��Y>5�����&R�����w�_�e%��]�K �����������>�<��� |��	����k����|t�SB%�}]�3P���2���f{H��Ix|����!��4�Z%P��p�m�(mVl�\�SP�hksx�Pբ��v�P���?���	]#m��X� ��ͭ��U=���ّJO2�>C�m�Qߊ{��A"�.�}Q�wߒ�j��9�����8&��&Ίj=-�=����*ؖu�FS�H�bIn{��� -l'�_kV
ɪ��!B+O|6�]ߟ(�A�t�uƵ�X�&%��|]UbN�44����#�$�]$�{f�����b��$��L������~������8+~�rD��S�T�c��D��?�\���_|A�Ä�%ӏ� �����������O���R~��Gruy�)�����������O�#2���ml߇6 c���6�?j[]�������O�������vI&+����;!�Y���?����F^�x΀h���ȓ'OX��ƀƃV&Ff}E�U�i�F]�=CK0���:��|��w�&2H�y}}�P׫�K���.�3�o�x�+���O�ʹ��7�<��� @�~ ̢�-��[5<�lP�7ӊ��ο�|�	���,�2��j3,e ��Pl�B���c�mq� ȇkT�l&����@�����|QAY�ȾP��yK;UU��Q�/�����T�q�����$#�|� hX����$��v9��SXA�Z���1�v�:Vˢ�m��H\���P�1��;�a�/�	�����Ȝ��QF���$H�� �|��x��y[
�>��ԇ=+�3�~o!�1A��@:� V4�D+���}vbze���i�HCWDA�� xE��FÚ-��D�dF`!��N�� Ʉ1�s����"�A�G�����#�b̍�r�!�������n��O?�L���=y��M*Z;����#iՎ�@���ծ�����	c�m� ��Ziu��U+�i%�YOa(��ժ~5����@�'�bT<�qn Κ�C�A���M����ev�5}�+# Q���z�(��]<�� ��;��^M�R��;�bF +��\Y�C`-��2�[������b���=PMJ�������ĶQM��E����,C��B�G��¼+0'PqŘo�_���Bu��p؛���u��j8��Ѣ�q������J4ܣMc䐳�[Uq�$���z�H��V�]��uY,�樄*����m��!��;&�  a1�#�r�Ya�����zb�^�{ ��g!���'�s3� uZ�ؾ ����J�'��>�ꀐ{��u�)�nv�%`�_�a�%����[�eTP6j�r ����ׯ��$t��f�1To�*�ks�*L�%��I��
S��&���@ؑpmp�0� �BR�rV�f�+�q���MH���[E�}{� p���	�G������퉆�W��jy����o ��	���k�U����?���	�?��������E��>�הּ��a�J���Dj��7b�W���N�W�̚{��X����u�c����1I��W�R���jJɆ���M��.�5�J��ݺ֝�/�&�%�B���	}�w �~��%ּ���܍��UihY��oe{����ѽ������۞���,��h��g=�[k��@�����v�>*ɚ���@���o�Yr�aɲn|ೖ�#���I�lx�E1X��j����7�6���?2˩���{�O�}�E�� ��h���Pp�@�u8�=���i�FӖ��r9=Y�D���U"#��'��ߑ���O���y���_�_���C�n.�4�2,n�$�}��L�O���_���A^<�Fr���٧��[���̏�ɛo���6������Fdlc����Gi��_���q����Y���grzzW- ���}�������C	A� ���s���>��O��O+��rr|*��?�������[��k"��V��nd�^YeY���=�v���V�r��,�jIT!�t �����U�'�C,��b����	����,fS�s����j_��+��׀āw��
�`X1?� C2����A�_��)��E�Ղ JIpژ7{��,��Dj%�vIY�y9 �D���H���	(�l�[` |��h�j�уH
ZG+��-X��OC�A�tSa����1~vr�l�{���w���|q$��B.��:��`��z��^�Z��U�B���+��|�����6��Gw�k�>����\C���U���5��6�������+�
��N++�=x��G��g)!�7��m����@��ih���ة�*Mq�q-늖>L~��}�~5+�6��&��^̲ H�'�\���+Ѱ�aia�4?�Ln./���_�|%�WT�����:�0R�1�N=�pH+�r�f$���fׁ7
"E�Zv!�%�Uv�-��m�lTʊq�)�����5���� �c�/{?p�����ڙ-�Y����D�h�I�
��$��':W`f�[i���fM�`��Ш��� ���� a�5ױ���j#?2t|>�-�^̦m�2��#��b�1����h��gs�%��LY�ў�'YZ���CA� @�d�>���Tݸ�nW�s��쐐��R�j�'A)�f�5�浌����ޖυ�mu	�#�Ǉ
iY�;�	+�}��I�֪A6l����Y��jU����)�P�}�-N�@@.�dK@�EJ2.Qռ���b��\�����U�ګE�r1��k�z#�gZ�\3ç�r�@� ==9�ߩ1}Kb�P,�@�ٿl6Xw萕������)�� �Lt,�\B>�9�' �1�p�������)j�U ߙ�U6Te����MJt��C��0�n��D��?���o�w�y7Ѱo�ߩ:	�x}PB��%�K{]�-%@�d|oG8ۭ4�T!��3��*�U��R�A�`��\A� ���"?�z�.���,hj5����*�DVLB�{L�Ժ�be~�ߝ)	�u���M�?��E�1�?6iov�z�ラ���\,7u�5��v�Wk��p8�ne�4��������S�u�mIx� �I��t���k��~�PUJ���0n�FµJ����}�p\����K����+���XZ/�=�L����+T]��]?`�A�qrr�~U�O�Z�)�wvz�����P4`�U7=��R��������}����t���0��'�����?���_�wT��~�_]_ɯ~��T~�O��F�U�D��pa"���]��?���������C9::��>������?�8?yG6~�}�ɓ[�7���mlc���Fdlc����o��������+�h<{��� ;_L�p�Y�*�) ~�A���Z&��ܽ{� X��\X.�i�u���a��~��'���+��j_ؽtV@V���πF��?4"��m��^B�,, �������[)���_���%4��ʂ���ె������Y�V/�s��� '��u� ���Ё�Z�	�s� xM� dˋ/̎k��R��>���k�Q9� ��J�T����ٜi�����K�F 4/# 7����|(�o+?�fX驵�|�4���a ��B*S�����y���|�����?�<Fe*Cx�=���	U��f��3����3��!	�V $+Y�LW!aR�Ԩh��~J�b*M����M�������$���.�J_�@�)hs��(Ҭ��DBd!�m�Q+�����ㆊ���T���h �����#� `fش��Z��L1��������c(i�d���g�Æ.>(����	���KT�s,��V�?���<x�c\#�4T"������SJ�����?u]w�!�y Ab�y3�c�������o���ܿ���H��dÊ� ���g|����6K2D��� F=A%2l�U ��������5�P|g� �X�W+��JTUT�Պ���\!777��{p����iKP�������P��b��d@���y�!�+?�ְb����V���.n���Gw�I|�8?��~�]�k��ɰy�`�Cm Rv��?pӘ<�_gK�җmB/ȊHX�Yq�u2Sb*4�����|kVn�_�kZ�T��X�$�P-����q��,��p�M2?��ܺ�(�J&�l��g�|� ���y� ��T�� HQ��9�s[�aV�\?��X�� ���ofS�����la���rk���F�N�AP��^�eG�R�����<~-�XG��
�u|�)j�')���P'��������X�t�:�s�1 �*�5&�5Jh�bn:�����.��Mp�Q�KE�����V8��iu������װ�ʮ/@tf��� x���8���{�rQv��cľ������� ����?��a�׉��[v놂�mg���H���A �C�>�{
�* ܠ���B��{� Zm��̾?k�3�u�x���@
A�י���YC�ŎW$0T���$p����w�pr��P ߉sS�>��2��!����NP�;�ĸB�����\�`EW����}�������נ�#���'��Sl�U ��v��*�W����ةR䝡&�l�{�~6�kWnJ>LZ��+6���5�WgD����,o�_�k�"js�rM�h%�8z�X�h���)�h�$1�%1�ߨ�!�*v^�nLև��N�D	�d���qXJ�r�~(`�6�ȴ�{��s(�_��c&�VܢykY<������r�{�l�`q�*��>~|��u����u�68X�<�����;39�����*L�ӟ�9���O���J�ǽ�$��?)�ܹ�����o�9����i����p�(�@���ə��9��љ?��rys%���s���6��}��H��mlc���୸\K�&�����o��oD��_�+5�@
ūH�~�H䈿�jX������?ܯ�ן}"����:�m�0b(+�81CU�U�MD��*жT@F�{����nf���n���7?��l)��\�#�g9~+��<X.��� �?���C<���)�IU����r���8_��u��n 9@�����T�~D����F<�`�ࡹ%@u zc�1Ɋ�6b�̯�� ���5����c��F(7@��g�ܽwO<x ��?�S��C��|�_��:u��5���@iU@P*�h퓐O�L��PPG+�����þ��Z�c�R ɠ`�v�d��V[�]����j��#��SU�l�C8@��va˺Ө���=j{�u�o�::�w���םT�:}e4�8 x�����Vm�X�N �}��)-wV<�xVЪ�� � �{[��dJ �4:���
�@������\]]����̐�TX�TF!��[ɑFU[,����pJ�Pmr(���c9�LD�s}Wr-��� �a���X��0�)�܇ؑpe�1*�����}��j�R�شYoIN��*�h]�q��e��jKˢ�f+��n�zpvJ�
�b�����(�ڒ�s.[��4T� ��zUXζ(���b}����E!����ORG�>L<���;����N Np�U��.��� �@'�������TS�>����<Q��@B�
���׉f��������
U�*��N1µ��k���*	ӂy+�}6~{8V�C�V�"R�c�c~ �#�c	*@ߧ�l&���,W��(�k�B��A�	�ӵ�:�6Cj��)&��]!$?���SК*���~��4
��Ǳ,	�&\ױ*��EPAr��Mt���0Ň�G%a��s��~Y�BsNB�f8�<(����B2����41�a;!y�5c��Z`�+���0�EH�:�_/n���a�����eOt;3c�ȋ�s/��bȿ�zX�X�0��$��^��D"]�C =����߶[K��N����eGԧC�HP��`�K?7[���3ڌ1�'��k^�Fj����-!׳هl)�<�h��S�
+>&`����:	�x�L�855f�B���N�Ե��R��`Qt;'$��捘����Y�y5�0��JJ�xR���`�W����{����F����s^�\�q�$W{�%N�N�mڙ�����Dӭk.�#�T��b -��:ťڡ)I�E.N�CC�1��� ��k�@		%�f��!X�p���M�}:X��� �"��taV|���A�M?n�T�}�w������= l���r��k`{���ޕ?���\���I���m��W����Dj����֬B�ɂ$��f#�痲�Y�t�da����w�~x�����6��}�H��mlc���8��K�7�<����꓏�@%�h��D9Q)����Y����++�݁vVϟ?������~��O��?�_���A	��\��|Q�� �c�����o�K��-�H�� ���W�3�#�!_�aP}� ��d�
�8��sY-%N�b/C�+�>P;�,��"QՈ�q��(�۵�K�P�MR���_%��5����Hf�#I�)��<X���?>2�BiaÅc�ë�� �H�R�
91�:V[� ���V��V��H��h���C�!���,,S�R�����m >|% ������Z��?��v'Hhk���xp�]d�A��� �@�6�3!�mi����< X�:d.QO��V�k�{�܄<к��tavJz�]��NC�@gg BD��,9ZG/m%;�3���D	Fl@I2P)�w�*�p���6��޵��\|���o����6mC)1��.��"v� ��j��8����^ C�t8��a�뛚�N�Հ�-�=Vw���k@RNT��/����ꐲ󮰪\T�����%f�UѺ�"�ǵ�̏���V[jU��c5"�-Hm����zBA+��e��R�d�W+�hGG:0/@�싒!�Q\Y���J�f����w��,��X��q�+��fdA���S�A4!�,!?�/�?�D泉_�b��9�Cj��hA��"9�GY�XH<}�D!Ǩ#K0f�VU6��T���l� �����T<��6� ���1Ob*fx9�#	 �T�3��qS��qoc�ʶJ�9`';�2��}�_�ux\jAN�z�5 D�a��|^H\��l��_��z% �a�d(���G�ώ@z�O @� Q+Ĺ�=����Ѷ��+��lf�!�kV̵M�I�t�q�Q�{����p�� �w�T ,m�VW�Q��ת������+�*�`Y	uN��8�eq�1,	c{"�)���-�Ⱦ*J��[�}�6q��������{�!C�\�FM��@>	�@��C����	��+^�PI�� �C"��}M_w��Ĵ�**��$]H��^a͋㐥�?õQ��γ�p�Z���DQ�v]�j��T��-R�iXת@r��C�H)L�b���@�G0<KiY�e�$bd���Ъ���"��ά�b����z����*��eP~Pa)TCQ�5k�!����T�	�_v��C���`f���p���ɔm�t$R �UiGb��"-JQ����a$�Z#��Ѣ �L����}o_n$��Dҏg��"�|"O�?Xu➐����iy�\�sJ�uX�����S�`�s>��T6�Y�B��f�KiW�Mg�8�里�ͮ�%������K�Y���]�G?����P��_�^x�����+��7�=ס�B<ĵ*؟^�z%��۟�������k�w���ɭeylc�����i#2���mlc��7��L�!x��x/�y&����lnV�������Qَ��  �R�P��?��\�|!�؄�ǿ�H�o����_����7�u�(  ��IDATn���j��d�`��	U�Z9�݃bd�X��ޜ��@�ły��j��ڛP~���w���O���\��g mՙh��;�������hB���a�J��yN�������Vv��̏rv���T��P}��R��{a���[�M� �����@$*8��6�iV�) ��L��%�e�}x���ڪ���� �ڑ���T-V���4���' �j6H
L�:�����ԭ����*U�dE$��+H]b�� 
�vu�V���@���
��� `�~_�{|�ã�����q̰�ȚT��s�� c
yY]�^���u
r���0��t���҇�G�߈���j{Я����[���R�W��8�n / ��n#�}�L���$����$�qp�K��A��WPk��f��H�>�<����X�= ��N� |���F�4��.oUSӣw�
mG�%�������W(��R���_8����
s���ȟ=s �c�ȥm�`Z��z��V`�Jd_�2
�f��P��H���J�yv�I*1�V����@���hF5���A����y˃���}���s�l���NA�J��p< �A��و�yܩ_J��$H�
�Ɣ[PJ9������e���)���������扰/�o��J�A*��Z��xO�� 5��^[Wt�8[QPٴ�r�����f�J��u�������wFV�w��6�������H<���k���ȪD$�@Ed���a�:-�p�8\O���w��<y�m9~uI�����q��-���vN��.�x��|b�J-�������Ņ�\�d��{2cP��ø&��H���@��XB:�� ��q >mM�M��_��J���js����'ȮaV��c�~�/�푪�꬛g� T�v�����ǎ��\룾J>�C�d�4	�C�3���}�0�;�(b�Z��ĵ���=s��4$P:;D	�S���Sρk��6^�}�5�尶��������� (C�����MT���/ʚʱ�t�פ��q��4�c� ���Ȍ��1����H�֔����gYm,��	�\.@�{ �}�ܬ��֢X+AbZ9�-��1��Zd��w'����z�>��5h�����וPP'T!@>�����j�2W��}�����$��T��x'�`myÆyL�8�l���������Kb���п�2s��,��q�X�-Ov�y6��bʟ/,�< ��s�V�x��S2a��"��Rm)Ԇ I�ON�������-��|�������Q~����=��3���a��=����ל���������w@������hл�Nelc���������6�����]����\���K999���l���lw;� @~���}�e��ዧ_���)k��@�!�<�mn�h�1�OYy��ت��&p+h��!������k /�S�7p�U�����e�� �%�D�<�B�B>`q��1�&��A�ǽ{�d1�K�?ȵ��rOK���+�J�����<�1�;N+�,��I�
��S���,;���M-L� ���B�8��@���V ��#����ܒ�B3��<
�"ө�=2;�\��*�셤�y�(&��J�!�$} 
Y�7le����\�p똺^�-y��:�$�bݓ,&�Ǎ��~�}hvVqb�nb�H
�����J���z0��A8�[��d�@��(�p��j��Hm�ұ�vX�n��9Cڳ�MB��)���4�zO��:R�	��p�)7[�Ҹȶ��\^_��N|W�H /Ě� ����J�{�@��9|�1>q�k?�כ���Y��<P R�Wx��4�;�t,���@�4�T����" Q�P�_���-�s��T$�Ԋw�@�GǴ����f����{�-lZ�����n�מ�J����q��	�0� s&���c�"��C��GQt��˓c�j#���}f�l��_]_�a������%ͪ��c�����
�����:��a� J[�6~�8@�9�����?�!��֬�ڎ�Pb8n5��cj��LE�x��7X�S˲	$U���̑��u�
U�
�R)��\�����2 �U �C�R�BE^2aurN�H�k��Г5G �'���S���
�*lyK)+�#*k�^!�O��B%���d.w�O���o���=��Ս��;+�>�YJF0C*R`�֔�T���ȭB�� ��?��U���B.����s��<��U�Ka�1'�p���b�Tx�ڐՖ���^��
��-wS�ք�d�����`衴9���P�����5cK�-`�����̧��n�a����N��1�[X���0,=(>p@�KCL$3�g`���P%He�){���l����0��S��[����`}�y����8��l5�$�+�|4�v����,�Ǒ�rvOe�;
U��-��-�5o�Xpn�U���*�spn��X��s��Ty�Q�>�#D�h�V-�p\��� <��1���bv����s��Y;1����V�D������
��G�
�
��m���\�>��k�P��uPE�xb����B�o���tc=�>p��m����=�����(D!��ߌ{S\��=�d��@@9�*����{'�,��`�B�&�H�N���d��K��2ω�u$�5�F�<>�����y�{/�����������K�`}=�{W��я�ѣ7�x^��?�[��ݗ/��O?�������78�q�.�>?�U9�sGD��I���mlc����H��mlc���hM޵�͡
���ճ�r��sZV9{N�* "·�=��j#�a�Rh)�������-X��ݨE���<�}�^��l.@�(8���[���5� �E��lp� � ��[�?� l��M�����q�?�0AS[ �\*���E �[V�!���ɔy(���=�3k��^���hb��!+��PUZӷ;<���i���<Z����m� ���{ 	T�T0��kM����J"O�<�7�|$�wΨHy��״9 N蟌�P��^9��`�@���u���\�E�8bx�T�����Tu���t�^��9�`��'' x)I��J���}�:�9 ���TCvcװ�Q��체L��#��#�xiP�;w��R�6T �
�|q�b׏�F�|��{�ɬ62]��'��pZ Cp�I~�
H31 -�)2�-Q ]��Z�#h�*����L������fS�ߣ�����s�,�nn������k��P�Ō��ZE�Xem??��P͊�`>��QK�~1]���s8f�*̌�-2��r9Aeu.��
8B���`����� � H��jx �e�~�� X�V�s��7���
���j N�1����F,�������Y�9��9��A���ӛ��L��CH��S�?����Rp��B.O�F�������,���z	��5�V�
�J���MQY����
��Ip���l�v}}pе��v�UsX; �
��q�t�6���ErJA���Ob+뮻q��h�: ҃��k�9�u��ص��ev���D�p��X!���}�R�V��?n�~��c����e�1�R�LJ�J��YM���� @�V~=Z��	�?E��LĢ�l��v�kf>�Պ��r`�3��c���������M�gX��Wc�-{E��4� �%2��p�Anp�Y����<������
�x҇���'��6����ZI����u���Q����@����@`�w)	�j���{��pde�_ 8����$��k���H��@�T�^��|�^���e5
X-�zR�:�|�Ha�Ҧ��%Tڪ�
H�������?��>�$r��KzNqG*5F$`�H��~���h��PͿ\F�@�pG�~��Z�Y���=_��2+���۾�21����mU�Y�k����8��t�wD��u�ﱂMf�4��Q���j�}���"
�>kvl��H=�n��vj�=�suvSƹ?Z�*�����:6�9�}��np/�
�O�iK
;���s��~�A}�O�lw*:��V�^ܿ/��_+�z �x��|/N��Z�>���+>���oM"�������?�?�PV7�\�����{��;��//_�h"���/?>�	���mlc�������6�����
�ċ��Q��k�&l7+٬�8��<=���Ъ:�1��zLG9�4<0����u�V����Ȍ�S�� k�X+�gX�G���-k�A��#r[�i��x��=��U�[��� `��� �N�����g>7p^+���i�r��H/���	�A���r�ʩ�G��a����9ɓ`/�8QaN;L+���-A���u��%P�*p��=��5p�
ʾ1�*��s��x�?:YҢ
�k�EBS�cK ךDG�P=���h	��Ω2k,�����>q�8����[�U;*������vC �m 
���Y�,�,CB�Yj�^|E�y��D�V�i�k���f�F�T�E�!��,B�����v�\g��z�]	�&ɿF�Xe���L�%�Bj��s�ZM[�FFG tX	lvM���C%s]'��UӾ���{�ND�o���Pe�*�UJ���xJ��'q�C�4Ta(%���J��b�����Tc�9����Gݸ��
D�Z%Aq����8���t,��^��f�'AF�m�$?C�>��1��	�c��`�d@?�MUR9�|m��du�&µ `=I�L��9`̭��gwN���)s^B�TZ^G%�j ��������5j~�sT�cnW��Ȑ��kk�\3ѧ��V�a)+�k��8�&
rӖ�d Pj�`���ñᏯ.��P���6�j�$q��4�&�k�)���ۓ��An��*� �"(ĥ�X
��s�� 46T kˎ��q���H��Y#���χ��Q��`�!_��	2'������U����pfL�7��q<������+��4����;���<�������w��LpH��� ��\G�e`��a���VMP,�-�`�8?'1]P�4$2+ˋ�M�ѵؾ��B�6д��\����Xw(��m���� P��L/�
��$��{ �A��-J"�ۯ�kw�sӯ1a	ڶ����@�ɍ�פ@������B��{��I�@������*1��*SL�c��Zw�ܠ��Z���;X��E�ܚ9�"�|ҭ�Mg�ݺà����UY���}t$3�+������B���سK��Z�!�}�>$��sӫ)Zf���������6���V��߁�bpm��T��-�|D�G)�eo�j�X��y0�u�����4W�VJ��pߦ�w��Ӛ��j�xP���$Sͬ
���J����=��0�&�w2��㍄����2?N����;w:�2�x�ĝ%�)�ꎅ8���Z2��o��5�c� �y؃�p��D��=PY��:�O�"���sŋ�lժ͆v��呼��;��;?䟦:�����/>�/�����Un�kQT�*��}r�L._]���6������Fdlc����o��K�曏� ���5m:�8�	���M�XUe�,	����� z~y.��d�9 ��f�����P������b�2%p�PM<};Z!��%"���<�	�P��=[.�Z �������0�L�İȦ$A 6��d���������N)��FLi�R��e>�I���W�_-���	R��Zu����f�U0���4�~_����V䣲��H1P=n�@��`9-�LI"R Pk-4��ZN���[���j%��� ���~���Ӊ�=;Q���FUsx�'Yg)�\N�*��: 8�a�o�ce�w�0Ę�����P��&H%Zy���H�*X@P�zf���ov��^��$xOC�B��f�C`9H%\�Aёe{DfoA�dL�5!򡕳M�Wi4w!$#D���' 0��H	�nm�a�:8B?�;a%ҘMm�`�TMŀ��j�`y4���U�3T��N�Q;��([�m��]J��- %�m � <��8~~��R���>z�T��Lv�׬J���pԂ�ܭ*���|�a�I���*��:nC�u��f9���ӳX�з`0<�wP��/�)	�A2��*����ah -8����I�1P�:,C��:m�[�������b���˻�UR`��a.	Ȼ�~&���6H�ǃ���/�I���w'~�ͨ�qАѶ���?�)���X�N%�f��*��K4H>(6����ʨ� �����jFC�*]o��RkB������z�j"�>H@ �u�A]����d�~߰��s�,�ڈJ� �Ee����i�ua�_�R����	����њ�d�0�$|�z��
�v.-����KST\�&�[K~��
9�+y��e���S�.���Kz�ףȟ�ե��n�h���(�5�k�9��9��n{ q�ĲX��ჇT��G�(6��鬘����*D�>���,&��V[6��lH|��:0�c �u )q������,�j���k>��',h锥�	�
����b�S+5D[w�R����Hu�Z��[��qj�
:�ju��U��@ԇ5��$�c�FÌ�p<x�/� ��B�3:"RK�ڬ��k?P�D�q�R��2�N�]�<�H|*�P��	��L$�jr�֤-�?��G\���,�vLr�7��P���2� ^��?*֌&�J�#F�����W��b�����l�p��b!DE�2e���Sg�r�P�����8aؚ0N�.�F�Ќlb�ɡ�1��&qw�~֢��`I�N��O����y����~�2�����=+l� ��wJ�##��ub�{�����2W�χp�������c���԰P�l��z�+Mf�#��6�y3x��fU�i�u$Ҽ3(�A���۵b�h�+X�j^�ޯMP��δ��"�c����������'��2my|,=�=\ӎ�N��'����z���/l�.#+%�� ��#l᭜�9���mlc�������6����� l�"`��a� 6 �g-E��\����x�*撀X�J���x!p��իBV���@�F��n+��D�Gr�� XQ�wd�����o�_��ͪ)��?)*���,�wv����J����_�|/p���2ͦ��K��V�ú �*L��l��j"{�8X�2������j�� �lb%�N��A~ �Q��A�E��Ӏ�#bN󈁴	9���?���z�P���m)QY 1*;+�1W;+���J�J����Os����^���K�y��>���%֝�Y���V7��n�����\�7��ic��k��f���~A��n����}��N�I*��̆(a���q^C�Q��TBG���5ϣ����h%��S~����A�#0�	0lZ�zq�J�=?��P����D�Ng���p��q�F�>XYKS���Ɣ ���,�Ā�87p׳*�r����Aj�r2Z��`�pӒB�T�>��I(��Z$~�gȢ���&Mfǌ
���穓�o�j�jL@>���|͊L�����X��}u��߯P���'Xm����2I܁Z�Ҁ���6�?� h� ��H��܋��� ��wǄ�Z�5j�7�qVT{Z���!��"i3:��aG�@: ��,>�.# ��r���\��9]�9�U��l����F�n�٭yL��� �	�SI��r��5jO����DQ 3�����W�d��# �`�E�ɮ��fՅ?z�P��<8�'Ϟ}#����T��5;l|���9���bV�� �1dE�b��4oǬuH�vŏ�'k"~���MN�k�cM��V�0��u:NAl�H	E�	�s�����Qkn�k{�
�����}������i�5Q�kI}	�|uk0��.�n�۽�[a=W�<ؒI�*�A@�ސʋ�g:�p�i���Q�2ϭ���������>�z�J>��W�����RM�?::���u���{�����~�q�� �w��Z,��3�~ �w�'Ӊ��)T\� ͻw���SΩ���8����-�z�&?�A~t<�3��D(����(UU����?��6ҕ�p��LQU ��x���|/o������+���^L}��=�X��h:�F�l�Z�xmJ.z��N��e1�'8N���<���������6�7���p�HɥN�`��M��r��X��\v�\�����>�5M-�4;
�����;Am���*��=V�>������e<F���#I�0�L����W��9,�R��r���.�<m�vQԺ�j=�G�@ޔ��l(t}�o6ײ�l}�C%��e�����jH�b�Ĝ�L���c-�I���l�[~Z�j�YlG�8�?�������Z����)���+8:��X:�i[��c��;B"U�m�5 ������3�d�ڍ�>���O$n`	e�&���I�.�����4�f�h������PK��q�5׿gyt�u*�|��9��p�9KR�{c�l�~�+��ld�>��N,�ݪ�ƕ~�d���;��,�9�{��q?��+3��:{��XX_pO���������j���H��1�c��O��ז���2?��Odw����~]\ʇ?���t��Oϸ�_]]��O��?�/���Ƒ�����~�ƞ2���ZV�����޻�mlc�ؾ?m$@�6���ml�\�/�������*�w��Co��U�j�fD)> T<�_�.��lxD��h���2l�G�+c�?<�>�B����d������R�}�s�BA2��
�,�>��U�M�t����М�X n���S���'S>d�E���Z��hУLj�����Ã  Ɣ���w�l�yg�� �ݖV��B�H�H��2�*$�V��6UE4�X��
��Z�c����:`3�T�-���Uh�v[>�޽{�?�Nx\����1���گ	h��u�PU*��b�<@�HA/(��KK�01��b}A��"��5�W _�Z�z����S�� ���>且T���1Fe`��ե�<!��Nv��N�Y���}R�z;�u� A��vT��
��j�����X�[���� �^g&���Uڒ)�C��P�J�F�e�k��Q���D�k��Yn����0�c�;��KsJ�����A�B�5���1���PUS�%0��jT�O���9y���!�E�냗>����^2$ �TEw�jlL ��C,���YB���ڙhշV�6�o�}*�������$\8��K�5��6�h?g!�rX�A3�1Pv������%����!?��}P��l���4�z~��}�A����K�V�3�z;D�q]����P�ܹ{,�cX�٪UM52E��͕�Kr
��$�Q�C�3��:FC�/Zb
7�m�{*���JG�٘-�&�K�0�o�����z� #���4��
M��J-��$�9��r�"�5�(�q��.Uq��1�!;���5�0j��i�QA���y�3�;S\�k�=p���n�-9�  �`I�X������L's��e���^��hy���H�ݑ�K��uz��<���g��aú�ۭ�ߦ�q�E�#���P��HraN�ED����2��Wr~~��8T���is�:�CȽ��h�5��8�r�!��5�;6���F�փ��@
�J'�;�$.`�_�o�1!��2St$�\��ܮ�$�9�BH3ZG�3��{h�E�,p}���~�zޝS�k���F�{Qo54̢	��0s$���`8\��?Tu��kP͂�!���筢? ��u`�ǒ�}�P�F,2�$!ek���Akd+����?�?~튠�PJ�Ǹx�#��qxφ~�9'���;�
T!�ɢB��C��"�1�og��	�U���ڞ�����k�gP$Q��XؽYM3]���5F�����	��k�'M�Eh!Dq;i�o�5�S��jնӾ��uUdp($*:����m���7����|&gggrz焖��Xc�c�����Z����@��u�_D����[�k�=�E ��؏%��L�}������	I%�p���U/
��i�`�m�'����6i@���Y#�9�bF�"�݆����C��u`����7e�����{�_���1�}�]��Ή��ޕw~�#y������7�p��Jn��囧/xi_�|.��?���mlc�������6�����47R��hmC�g�>-�rZ�����C}(�#a�����%��HZ웣���A��Ā�V%���v��� � v�;��� ����$�OQ�e�h���B�����ğ��5A��?�pD)l%�> B��\}b!�)�fPn��~%�� �ż�	��z��y� S�
�=A%T��n��R�W�+`Z�o�j IaO� �p}�j#E��1k+	@�e0tT-�Pb�@EJ�*V�,L"��n�ti,��A����m����Jb�Y''KY.�Y�X�_:m�� !��J��N���[�o�j�+�@y��7[��b/�<�y���/�R&���Cΰ��� ��DT P\��K�y��� n@x�I��޶9N VeY�*#��:���V��"@�,�4��? �M�a�qr�R��Vb�]J����iԖ��o��4t7��[�ho�SU3ѡډ8F`K{�+����d�`a @2�oX�AY�
q����F?��i	��$�,np�:��%���S��)�<�u� ��w4�E�.����F�#��p��8ٯ�]h<R��&�A>b+ �p��" ���'��.J;gp�Z�t>�%�V[V𫽐_�{�I�0���D`�6���H�����,�OW�(�����@�Tsmj�����h���m1�ʉ�ܳ�c9Z�8���ر|p�$\PAo9㎕��+��@���vZi�s���b(y�5�S�;Ɔ3"��#�ǲT7��I���I����'2�$~U������?}jyM�EC�	^��S�(�\����`5���fD@�VȎpi-��v�7p<�5׃�� ����C �s���}�PA���J��x!�_k��u���L�>�j"�����g��~-��`��XL��
6n�ϴ"Q�]��)͞
ʀ=?O-�Z�f���rYoV~<��.�m�n��E��G��
?��윭8�W�Tm�
�řY	EJL��W��Q��@� Dn���*�cQG*�����TIs<�:j&S{+��T]uQu,�+ޏ9_�}�D Y��7�	���A}��279$��	z��p���p�97Q��N�2�Z�Q$
t�L�����%q�\����yXj��hR[�6B����\N��}F;K�"��'��f�9��mk
]�!(8%ĔV�m}��&��6��t�����V��`�bw����4��/���Xc���W6�c��hl���BՋJ�1��^��m���`K�E��muoGFTEu��}ԆPyŰ�kx�;��;p���s��HPA�.�3���� 	��,X�@%����o�`�'�[���#	�TZԐ�LU1�3@Xc-��b�u��]&����<c�+�W�k��l�q�`�T��w����� �'ȃ������|���rv���{pߊ5ڜ��?`�c\����ϰ�v����]�����T�� ��z��Z�7O��g������ˋ��Ç�dlc�ؾm$@�6���ml�� Uh
TD��X��l��
��u$Ev�l*�z�5�0OH���<�'>�2�V�	G+����e��_���?8�"
�G��\�v@�S�o�6�v�����l' ����������Cu)�¤Q�����Sw	�J�^�T#P��A�Qґ!�5T��bySf8S7�UFd�p��S�� ���;� T�>�3�|t=ٴh�sf������JqP/eT1�  \ �7�7r���77��9�����oT/� f���ߍ*�ʎ������7��H�i&|��5��9�6 �#��M�� 9	9+͓�v��⠙I���E�*n�_��5��]N6�	B-�@��� 0�%q�t�W�l��s1�u*��-*� l�U%�y&�7
�ӿA�Qb ��L�F��bl���������	d�� l�p�u���)I��I:�O��[�H�� 8��
 �P�u� ��;Ѽ "��25H�;��CI �9YF@	��H��������S�d����C"���mfK2*�JQ�Fɑ���r���U�(q�si�{�t���_�`����r_�Jh�כ�rA U	#�Z�y=Q�
��Ə�bg!�YL��j�4cp7�������nV �\�y�r�� U�T���vBX��bZ@%| �:��s������#Y&���[/d]�h	�۬_p�up�W3~=�F�ѩ�]�_~C���NTI�Z ��h��g����H+�L⺜��H<V�cݴ�y�uj�WJ��Q�͠ǯ����Ѓ��|�G�8�~Bw�ZUx`�Tv���C I�*TS��U� 5Hx@�_�ON��(�>�B���|_MV[٬�8����`��=���9*Ϟ=���uE��Ν�V���|��2Os��ܹ����ե�WW$)A`'~mX�Dv��u�l�y������N*�Ϲ�6�b	�[��'��s
�9�CQc�߸�$C�����,d�hߖ�H��gw��f6܃��C����AR_����~셩�f����N�܉�\�W�B�)<�'E�'�ׅL�0���1����I������	�ё�����6rD�H?f����ʸT�6���a�p����C�wc�K��"2<�H-�4KJs`@���oy|*����gZ*��9m�Z��C�������Iw�
+��%�
J2�o�;�;��1�\��������Xгل�	ɔ�k�y��T�{����n�`�������1�}�+�hHJb�C>�j��v{�"fPC�U���KDs�b�GA�^$:IjOk<�dAe�^�ؔ��e�p�Xf�{z��ZI9�w�\ߴ{�����4�4��Y�	�Ub�3K��O�[Ұ@�8
��`��`jv�����kJ�6Aa��f��ڏ��}Ϟ>�����
�����v���T�����縯���rv"�5$�`�
�3m$���O>���K���w����s���6����o#2���mlc��5>��g(�>(A.E�, ��L3X(��A�j�������-3��^�\���y	�*/�����X����\_��ڔ�9�^����t6����"6B#< 6@��A	<d�3/��B���^��?��
'�lqG���y� UK�Y[!]��Ɵ�Z����<u����7����U��r�V+sYew �S�
� �	
|s���Ń>��k��I�>X����dV ��� c�Z*�@� /����9��_��ѯ��ҏ�HN�x�}$G'wYq�$RK�X���zb,����u�ʮ���A^�<gFF�������ޡޓ#�0�X+�벖��^��jt�rv`��6�L���gG�Ǳ�r@�<�ߋ%->ڶ)h��uڮeI� 4�{P׮����!@c�ĝ?��{�(��~�>.���v�VeG��jڒ�.����(&�(���A�*+�\��z��X���H��g���J/�֡�M�H/
��JN�zAp�UI�v��: �]���� ��f�<�@�D�]�浱�߲����Z镚��ɜTò�ߴ5�������I��`�U�t����?�� ��0�X�`ߥ���Q�:�� j�-�s��Ϧs�1�%��&�RZk9�U��"D��ՔD$�@�n�4�<����D-א�R4R�w�Z�%F��Uc�qڹ�N*?�B�#%(H�DJ0 �CA]a0-�Pf��aU�d���x����5�g�m^����׶T��������a�N	���9�2�ASVZMm�0>Qɋ��"�w �����+�A�����U�1"+(/R����?�c@~��*J4K*�¤!�z���ǉ� �6A#uyu)W�-�� ����`������R[F �T`�����\5ײ��� 2�
�\�g��=��o�KH� ���p*|�H!9s:��j$f���1��?ǹ��P�`H�+-h��w��N��@\r_J���j�I����0�<�ɂn�N׏>L\m�JSR�u��S��"
�ɒ���^9'=��A]�֯QQ���,���W�u��5	kY�����ٺ	�[ �{0%1pO��?�{�I�1�+(�H���L(`����$D�ڂ�w��m�+���-l��*?/v��kaE�_e��� �ǒ(����k��!D,�M�ԘG�C{�UQE�*��`eK-�E�[�<Ry��ם��`/���닿��ŷ�8�vi�����a�'G�ȧ�,��2%�c���j��l[͠�U�[*�S��IU5����m�I
Ls�'��7�����D3-��CQ	�J�I{��5_�{Ydt�[��b�`��{݃��b�`�T!E�!�/iM�G��V��T����;�ju������Z~���䫯��m�c�����3���*�����q"���ȓw�V�a�
�y>c�9�X�w��S~�&3Z�9s�"ک��9��|��_H��<��~������dlc�����h#2���mlc�/�UUm�=�x҇p<������������K�|��IT�o�
��ԇV�^xD-iU�P��\ʣ7���$uxp-�j�4����Ml��aZ���a]�(��'F�h�g G����U���N�w���YË������1�Zx&9ɛ��Կ7cE9"8
�1\@�hW����SV�J(���� �f�ᕰ�(��_�qpT�I��J��^ⱅ�Z��6	Ε�W�?�uΰk�Tų�l3�������[�Ƚ;�e��z��g��b� x�ϖ���ڨ���y�`+ R � X�\^�۾�mi���<:^�/�=�����A�e9��=��JC�� K��7
�L�܏�S�{|7���� )��w�,d
^�1o7�?�7�;�z�s+S�5t�!��� v�ʱ��

�n�U6�2�!���0�(T���
�
���ֵ>��%@H�e��-��Ѩ��0�Q�2��)5"�Z7V*�܎����}x0[� ��:B$|�y���`��Q"b��i;��X���"I����SU�ea��]Q�d�x�5iE,�$��f�p���X���9MK��o�r�[����G�9�87 5I��t���+M��V�s�ܙ5�0$;Δ���P ?�TQ4U2�`�Ѫ-�w��Ș��L�e��l*�GK���kZ���әԫ!bwP��U�X����a�=`=HHb�cWI���dHn؛� Yj��a�0f����4
��a8�(�>�f���`��#6r"( `��b����@eՀ�m�S+�و����3��*TD��
 (ǋ�����3�x��j�ֽ��0����_��o/����yuq-�ٱ�~� �nv����a���߷�NN�����®^����q�� H�"�|rb}i��	�}�s&�	���sX�����vM2$�f$��@ kE�hHĶQ���S�����-�j�?)�KPy�,��u��0�yY.�����
�Y b���C�s���7�� ��k:��d��)T]�R����ǂ~�h �C6X '��#�cPs�1ĵ�>?�y�#��1��RR$�e��C���.	�|󱨅]X����(a�ŽFe��^�V��&���B��1q=P� ����ڔ��7�5K	��(i�����1��'M3�z�*(\�@R���u���{�t�֐O���re�j���@l��sZ�5J�[��-K�<��;�����UV�ϡW��=��[fm����R{���%�1'yO+ǹ����ʃ��\����a��$��1�B��=?ٍ+����B.//y/��@^
���0E+�R���W��+�I0L�3�Qp�ƽש�V��������s\+�����3��o+�ݞ�#~5!I�@Q�"&��\����mhU�o���o=��o>�{���7k�}�� ϟ��gO��urOR��ÇT �{1���{�O>�������C����6����{�Fdlc����o���,"k��-JQ��I��̳mX)�|���+h�Z��'��L�E�62L��cx4��G3���j(ч 2� �W�{�浨�6��"����D)l(>���`��=��ǿ���
�Dw{�Ǻ�b��b@���b�ʎ��n�$[�k�����<}����b5�& ���1U ����;#<��)����K���Y����(L�qW�����M7mH��nY?Њ���m���4<10F�>�=�����ڃ�C�#2��
 �/�/��W�o&�}�>7�����;i�*��X���յ�ۧ�i�������yk5-�P*%_�J���,��*����ܫ�{ -���b3��ci8F���J�H�:���j �jc%���Vm,�9Ig�%�4�N����QR�A��onjݵP�l�����X�	"1��Ȉx���AΕ{�h�e}�P1�c�,b<��)tr��,�b���6�����&���1����hc�� �v>�ݸ г;�	�᭑���9�Ѭcڭ���S�#Y# 3#��U����������˟���Ԗ��GT:T����\d3+�^�ʌ�#n;�q�>��ֈ���bI �5׵Og�C�t�v�{��ZP�5T+g��F�b/������7h"�iK�H+�c7��b����Rx��yԼ	��!��v19L("`��T%��֌��
9�f!o'�&�E�?��tYv,ʮ��%�:@%3g^������W�!�qľ��&�L�q_]U?IIאd��!�v��h)���u��NE���&|z��/��e����މ��&</���b�*�V�7� ?x���Ϟ?����[j�T]���d�^ӄs*���A|��ם��V6ֵ�}i�1_�0���얅�k��h��RqP1gʯ����k�b-(�d��%�������4��J�^Ɗ��`g�t��̸d�6z� !�<�ڪ f�
��-�+|oP�{��1�e�� �� �a��c����;�p� ���*���#�@��
R�kiv*ݟ����I���Ug��K#"j�1U��-i]�1��@lc��-��[�,��tj�WX�9) wV`��$X�﷕�&������+�Ü�MBYZ����� ��֓���6�1l�Il�	�l����ׄ���$&�xM�		W;@��=�5  ��=� !��G��/,�ש���]���_�����m�p�H1�)nnV�G�����"�K��߽����CK,m�m"9����,�jX�m��� �Q|tt|D�O|�
<�z`��JnL�	����Zd�UT�ą�9��,�^#q��_?�Z���9=9�7��!��<���=���?$yv}y-�}������JNNO������W�c�&G~/=�R>���>�\���ȯ�_�޴W�-��6��p�^�|Y�tu��N�@��_� !�B�!����@����. Ǫ�2��|v�9k��="�P��2Q���7#����f��9fg�����O�?����g����u?��MmjS�Ck2��MmjS��4�n��Y�b~��f��V�2
�+ �8p��n$>�!r}sͷ��Z��V�Ϡ����C-�{�����cشm52lİyҴ
��k�
��x6n��Y]�fCS��I���k@�vǲX�Jy��~��ܰ4H����MR�fƆ���_�C�D6L�5냰Y���d>��/?+���"!���O��X!1 n{�^\��f^F�a��~�.`c� ��q���*_= hn՞���٫WR���O��@|����!����N~���3�c ��UKЗ ��X�i����V��	����X �5�"�,E���CXW�Bkw"�����/=�Q!�hzi��P ���eRt�
T��V�i�$��a�H�R�M�u���(��ԎA�>��������ԮEgW��GP�$�h�NdQ��p	D�R�D�Uo��h��1�����YX!;�M�q��@��+��aw�,��5�"��O��)�*i����+�A�8��̂��V�:X��U�����'K*@И2ѓ��S���e��#ȨP�-�6�� ���lEum_;��`T0w��ܙ�^��Ú�Jx��!O4kE׊�T1��W�����[�C�2��
�|.��6��O��w�@�\��FA�z�!�H;�p����e~{'��LN۔VW+x�����`��J#����۫
 1H�èn��g�F����o��(��k4��_�a��悸z����U�qdY84q����i��&iH��F�Ǟ�1��c���3ʦ���=d�: D�c�]�=�a~�Vu�$X��!�e�\��E2�|�Z�Q憄��������{��|��]ON��A5~�+T�Iϡ�I~����QU��$���K���ϵB=�W��DU�:d���� :lY�>�$mA�������%� 'b#�l�{J��|M���a�{��5>�"�s�@�fڧ�9�=�8�{��Ěp4��'\�?}�p{=��s��3��+k0G1����t�\w�s�d��]Z`9��V~���K�ßoP�롿�W����R)�,$�0�x�?~�����=74����U1Br��q�������_�3ܧA`b��A�y��#�!Vr�����2�D��~f��{x*úVAx��;qd�1��m����l��DW��s^C�(#8FRS���YwV�^��=���)�5m��~�����������:�;#Sy��t-i�ЭI�'F&'Cd�3���b<�P�{3I�D���͇�|�o���c�����5c����/@��cc��2�(��3�5��g����K>R������>�#-�Θ��W��~�o<.c��TC@�
s���U���c�\���4����Pl�v���ۻ+�9�����xC3�@��v���|�՗���k��O~�k�y|�_���}�&�}P��ɛ7od�%�~x˱�'��\��y��[yz�gG ?��IdjS��Ԧ���&djS��Ԧ��o�n����;�@�h�"#�7g0�h���N+���䇏uU���3�[�4c�a�Ñ }�0H�r��8�|lTJ���/����� 3�	���p�=�����(3�y� �'fO��>� �5�w ���zu�CR�>���"��Ԭ�/s�{�:*�Pu	Y?@= �ؤ>==����<^�!V�W
f�ʾ�/������<m���Z��dX5���D�@���1�� ��r�o�^%;`�D��j#��v���u�sW���f�b}���4�)+���O��4�I��$b�����VN ,˥��G?��B��(��dG�u�Lh���2G�u*�k��v�y=���! E��ꦧ��`P��`�U�Y͏���#2D�Z�3��̌��� ���6�p�����{�.B�H<h|�W~D��N+i� ��b�,��c��:���BC�3Zc1�;��CSUcq�,~��������H�#̟��J�5�L���-L]H���S�=�tv�l���4@N��Q勊^�/�m���E�C�������s������@$\󕂖U�j���Jc�ϗ$�8��?����ްb��u��� d��1�8
�% NAD��V����IU!�h(���QNZ9K�60t��Z���pM��I��(+�0�GB�FnGR�0�?���4z�1���g0;+�� ��ã�H��-��W{'�υπ5\[W���Y��R�b>	kQX/�-�$A� �p͘��XT��)��'�`�qЊ� �z��Ѱ�d����Dk�ILX>��,t��O���Ģm FTV�U_��T�P�,�sZ�2f �T����D 6MG�wMhCf+�d;C�m���*u|&�4�$/� `4�Y��Ǚ�b,8>F��n̖�Z���	�"a�A���w��N���[iP�@�!�jц�~T���q�u��wE�����ߏ���"�5������ ���߯�w{��u�~����#���a�F{!�_� �y������<f�Q�(��w���~��	_��[�f9�Rаn:��@}6�,��l)ϕ�g���X�=kd�[[����!bSu�5�E
P�PyV������Y��ſOa�na�j�V���Ѿ�Um��g+���g]�c���h��OG��%8g����l��g�Gag�k\����������,	k̒�L�`P*Da� /�GHR�~P�"�kY��	P���h@��X��~f�&�FP�`�,��y	�����7'U
v�ط��c}o��E#���Z��(�	�����k��� V���K�G��a|����o�Y}J5G�5�52%�5�g��y����M*��Qb�N�V�b��$,��0o�����>�[̩0V�f��~��x̩�A1�쑙WS��1�^ƽI%��U��56%�:k P��Du�j�@\	�c����mB&m
A��E&I�)	�$G��*��\�$QN�ܤ�X���'�����|.������e�[��)\�J������[�{X�v����������Yf����8�g�0/�&����A�p����_����LmjS����8�D�LmjS���~��!�4���D��W t�8�K��61�����jr�u_xO�(����Q6CGT�Ug��훷�~Z�v�'J��yF�G�h�M��'�2�"���8�3�3 `�mOZȍʻ���b���Gu_��2^�G�jc�+6�e6�9s�fΈy3�r���C�<�æ����s���e���|��+�? ��"�U��UMZX�U9�=$�   <�A�qD�bi$6Ŵj�  ��6��0��EAN��	dO���y�o������I헋9�Qm���{i{9�M���u��p�i��t �ł�C�V״y�f�C:O��$iD�O��C�<������r�}@e�2�`��/��.b6:mtZ�~%�g$�`Q��
�0^q۞�� 	��r@�R9[�(���d�.%5�% �$����>b��8*"^i9�|���4'�ώ��Ƒ���P'�{��@�@��V�����Mk������
v�y���{����r ���]��VX "�Wj#s}}����̚�r8���f3c�0b@ao��]COR%sSa�ZJ�X��b'\ׂ$mL��d]$5i-GEPL��cH�P)��u
T����̆V���>��[G�5l��
�������U�'�먎�	>V( ��>�Mk��Q��A��B�X�� 0���$s�6�%�����ϥ��VRu`[8/�lZ�4�Qa1�ƫU���f��գ*�����xmE��� 0��@�S��$��\.��i��j5uo�A���wk�-��v0���������H��
�dΠB��NHj ��	p���C�9&��U�m��8�K@��$�-������ȃp�>�y#Cxoؗ�U��j.�j�p��z�{ֻw�8������`���3A.sA@���*UV)Mp6��v���N���͵fN�y�X?Hr���X5:��ҁ�y!����s/� %�U�Mը�6ICZ��n_�Z���܅������p��9���_� �A��HW��z��\�ӲdWB��lT~\���"���&F���ߥ����9�������VL��K���t'F.�"�S)TA;5�#��~�P V�Kcu��߀@l@7a���
X���	���%��Hs*1v��M��k]�����T�H���}�R��k�^<w�}�jB�������.��L}��o����@���mwVz\6U����g,��@�$�[��Vb�Yz�:��V~�Y��3��j��k����7�����2�����۫�
]P�=�qӎ� ���@x߇%nS�_�&�O��I�h�D85�OB�s鰎¸jU;b���P,�����nu��)O�T�e�!��j�!����U��� ��Q�����JKU{�'Q=��LU�$ʻ��"��RX~	(!e�x��MmjS��O���MmjS�����=+o	TK�2�AЯ�����N�IF�jM����-�
Q�dA� ���
+� �j��6�mZ�5�u����p������!@9�,'��	*Q��7OgSK _���Cţ��+�������krQ�������lȩli��`~��?�/<�5�R���җ��#9���� ��4c��̪`�����|�9 P��,B�$�-��^�D�bƍ3@�H�`%UУ 	���j��-"n��(��vg�~X�t�U�9Gq�js�KV@��R>�y+����H��}�=��D[X�<��u:њ�Ҹ�M��ga8�����a�du[�]B��Xҟ�	@=/�0n�O���YQP�"��; �b� d�P�[��a�^�d4c�@)T���(�	ԋ[�� �@�����&�Z����@��m�����C�x��`+fZ&b�e�= ����įsb�[
2���ߢ��ā�O=�|V�j�R�H������圩@ρ+��i� #�㼪�O.���׼�Wm����e� 1P��Y:��a�~�l��HՄY�e����x��&E��|��Ym��f~kZ��5$���¤�\	(��6e�&Z��k�J�<5�/]�<�9��y9���˹$Ǆ�����T�h��u�h�a���"����R^�5�e�s��W����)L��#�A���,�x�X�Lk�8o��'��caNLF
�`��c�ӱE����$�b��u�V��pɓ�Y)�qa"Jk�q��"��W�cu �uU�&iu�EC�����=�Ц�# ����2�+$�.b*G�YIR�����cX�@M��Z6I���Y��������*,��<�-��?|�H�_�ku}}%��9�����q0zGbdf�!����9�1�����F�Z��[a6R�U���e!�#6 �>��VA�E8X;rx��c���$F���t�`�&n�j�8'Sо
�,����4`�]�Q��ظ���[d�]z{V�Z���J�|��1�C�{z��Ա��{yV��&J~���>>��3/	���L<���T�@�z���������L������g�F>봐BlgF��@L��]�L9UoT��-��%,����/i1�}�� �*WR����LcU��B1R��<TuC�b�
㼝���g	׬,�W�S�L4^{��A=�yfΐq��#�hh9��`/�U��,��soNؑ��u",��؁��ɀvKQ�ګ�k�����QH�yC=���Zl@���N[�l�Rd�c�湌O }8ڵu|6�"��UI��1�Y����)�gO���#'�_Pi�9�����L��,�\�A4TD/���$�Zڢ�$���/�'P-�z=�R�}%�X4@�}�����EZ̆��Gޗ{%��(2k�pu�=	��$f��A-(�����զў���"�pNP%'-_���W��̯W2��MmjS��o2��MmjS�����^nn���:aU��h�@۰�9����=HX�ܿ����,mSV&ϗ�h�� +9˙Ta����J����>֐Վ� i+I5 0[�M�V��Z)$(;xE�ٳ`����f>l(qd"��
��Qb!��֯Y!�'��'z*wGYo�����f�pL���7�	f��F�����{�\��������2# �U��V������^��dQd
Z;ts�g@s���ߴ�)b�;@�l��Vl�;���P���<m6�<m7r}w+/_��*�#����\�>l�-��3D�\��� ��\��B\P���Q���g� ����� ;1l���c�}A�wD(�L����@�� ɩB�=E2��>l�������E��`�<�1ǌ�I�g����	�x�p�����o78��J�~�ͧ>=�jm�*Org�m��o��h�H&8�� "���p�X��h��@���x�4-搏`61n�9!z1G�;r��w�`�hK�w�¤��6&Ѱ��3�~T����ꪮ���@t�*ޅ�{�v�RK�x�F�$��a��^ёX��@�N�. 4[Xf�'
$*��[�������ź�JC�q^ Aq]hÆsITA B�v��i�_YjV_q#-����>o�j�D�1��q�Kàa�bv]�(�`j�:�"7s� ��@f���@I�����4N���4@`�H�+	N��Ǭ���
�i���f�3�q���U5����p>P����#-�x8��F�TYê�X�N�w^d�ك�w��A�8�p�$ՠ4H��q�܇���蛰f�m8�|��h�$ԠB
 ~��$=a=��EsU���������G?��A�h�m�%	�Y�Z-��剨�ЩR����>��7��u�EI�{h�j��6A��8�n pm��~�CNa�⪕�W���Z�(�����p�E�9FV�I\�ػ��b^���
J��xp���J�p�Ϊ	� [Sl(��D����:k�o?��(��둬�'6��8N�������
��\I	�}�-�FBŀ�$������T>E#�=����A���>OI>�b���'�ъ�Y�����
��
k��:��2R :1>�OR�}\Ŏ��1r�>�=W����Zv�vT��{�y�`�RG���Q��#��T��x,^�A��=�hl���-� K�Yo+M����u=-�b��ҹn��'�ۃ�z-Z#��ޅ�����<[���}:Zb*�1+r�"{HӞ<P�¢��s�q�o��y��1;�$�S����|?SS��$�@~,ºCEO���Tm8���ah$P����q��
��P��.1����Z�ʪ�����8?�/���x��Y��� �T�&6Jx�/A�X�*MY\R����N�R�$��+��s��^�ks�X�P*�1��N��ejS��Ԧ���&djS��Ԧ�;o�8�R�@�ݎv2=���r}��&�+��*ljӊ �,/�,�ju��W� ���$	��fV��V.2\�7�a}�mCd�MRq3�?Z�lh3)E��zn�5�Wx����-�*�s�%�f�2�ۡ���.��ɋ胎@KZ�%���G��ZzC�qj�c):�� �}��$m�����v��_}�k3H��fG�dB g��d�'*��D��kz����HGlP]��j��A����ln+��A7YZ�D���zOd��q������~�3���ߓ|^��n%˫��>�	��7��XS��U���S#?`����C��z��`���ǉ�۪w�C߭w�0n2�7+�a1�/���2��1�O� ���ڰ%�ޫ��0K�HP����U1����P��Q���x#H �����J� ,O�+��4�Ӝ��W�_�(b�)�Gƫ�JrXդ���b�������>��Xq������o�٢�JCm�x��V0/A<-v�N;��b�G�����̈'Rh�w:�؃�\�cUs�2�q�c��d��cw�q�w��e�n&f�h`���DN��sk����JV]�J�V�U�9�PT����C��X���U?5��Pd
�.���ҧ���8� ��#+$���f#�B�?�}m�eZ�3R��8է����z9��P�5eX���t�HKb�]�D(�q���vl0B�*�U@c�g��k��Up9"	�u�e��<���Z��Y@�*5R�/�;T�*lS�8`��F��k�@9�L'ta}��/0��׵�w1�}��Ы}��J�F��O�j�; `�u���*T�p����A�Y=Z$�4K!�����>��۵�|W˕��p�쪣�N�0�#��NR���臆��<��t���˗�3D��A�m��]������׻O�攘mX��ev����y<h�?| q\�T�`��`�A�V��M��(4X�a<���:�T ����h�9�V-IRVŷ�Y3�_XL]�<�U�H,�:�VN�d�@q[$"�ETx�� Ƞʬ��\�9s�X����gA�d�1���1{���/W�`M�zuuŵ�s�Bi�k��H"*4T��5�vz���1�U]�t-��>�������? ߉#o��̊E8/�Y;f1Ŵ��c:��3�Ӄ<�W<�g�grsu'�r��N�y<����U5���q��b�����n�; ��Q���h�F�@��E|vJ��DQY®L	I15�Z�}�.�4�Ϛo�U�H��� �����<j��r�dT� �I��MX+�V�����X��t����X�萭��^,��~B
�YH!�vA>T����pBZ����,�*��y���I�!�&ePX�����L&j��\Mk$�(���D	�ek��k�m����qۭ�����6mS�W(x�s��j�����>��t܏Ev�Ԃ��	�HU��&�R�Ǿ�N����H��Z�6��Mmj�m"@�6��Mmj��V!��$2=��V<"f?_�7��;�@6�M��=+�Wa��V!�v{Z1@$�n�PA��2<���CAQ��!���� �{���&����-7駺�u�2����<<��؁@��R	�iN�H�Bk�.3�ݨ��-��a}�M�c6�i�%���=7���@�#ÃV$���JT���گ�<A� ����_(knno0T��j	x��Pi�u��9٨����U�E��8�A���*�B�/�����[�UB�����N>l���;�õ}��|��g�ipb!U��h8�<+B.�~xE$P
Vk�jg�vY�k��!�q�#^W Y.H'�[f�zc��v�؍���"�5H�~���(h=9%?�0
 �m�\��3�Β��� 5C'A�?�19���� ��WL/"���pNt������A�,UB(y���c��j�9��8��js��G:��G!�$�,H�kE]��D9a�MIn8&�$��ni�{��][r�X�,��FL��9f	5��J�n�.�m� �W��r(n��G �gF�S	 m �H�6��!ad�����)��Zc6]X^�UM�E��#���Q��3~�IYm߆�!�
YF)	�n�s��PI���p��RJ5�v�0� H�Y��3���>"���#s��P��z�G<�A)�빋U�CA��6�f�$��p6u��E��SKW1�ʋj��!�Ο/2~u�J��&0:�A:�|A0ֿ
`_�����~�|��nN�NV%S��^��{ ��˼�BT�E�o�>�����r��3y���f�uD���1|=��\Y.��K�>{5�*��l���l
As��L�� �5�B�,K��f������Nfw��92'�oxLm�$�fL!k�c&�އ�4 ��A�������Q��U�X���(_'|����	|91��ȥ��� �5�$9��F��]�z5�Y�6r�u�+I<������b_���_�U<���>.׿�����-f&�[>R��)Qq:��VgK-���u�!
F�����/�-]���� <\�u<�g+�{���������3�`G��Y��z0$j�c^�q�bx8`��cd,eь�a�9��A��ww��8��8'�)Jt_���Rʩh�3���"�ݘ��'�!O~�&Ӫk�W���
����9�{}_䗘J�$<�oC���Uf���(G*x�7�2���c0�Ԧ6�xf��y7�[��u�%}qc�Z_$�N���Y;Ju���*G?�Ȕر��QXsϋ7 �(�<�~�Bh}˜�T���W���7�g���Z,����
S�T�LXh~��Tg�3Ě6C�G��Y-�`�]b�`>�mScfQ����h#��(�)�B�6��Mmj|m"@�6��Mmj��h������� �)���oG;���k�Vn�A��*��@�氧����YO`gנ�����P����Ii�bs�K>����Vs#���"�p���*�Sm�

l���J�}H�gj$L~�Yq;�%A�D-�H$Z��1d׬��^R�ymh�Ԫ��]�ib�l�v��i�A6۵ǫ5G+�V�^ ��\�u���7�P���5p��M�V��I����[���@�έ~�9�Rs9i��ݝ�^iW>�q��}�p��ϟ���!,��R `�%���*?���{��$W���ٰ��d#�9 ��p��ׇJ�UG�<5��@UsSw�?��~d����ջ��f�0�%	��S��jtf��Ѯ+�>R�z~,���Br����X�Ƞ�6\ E�NL� ��Q�v!�:�V1�..?粲����r�mRR�5ȩ���ȴ*{���Jmdf��H��Vw��p��$�W5��)�"*@ ��6��>ZI|D�a������}ҩ�;�����^�LP�����2l\tB��1.�ܥ^��U�T�D� �	ަf�2DAka�P;U=0[�@��:��u����k�- �A� ��N�uIDp����A�fGb�e�}$Yt\����i��k.�F��xP"�&Ҽ�[��q�v>_HsR�v�
3��j*��j��-����=<�^���,?���@u�s�yQ�v7/,���3Zz��:v�|#\I�|��ɠ&Q@QǍ޴����P�X�Ϊpc�
 1�/������f���#a����yYȢ-yLT�u������od��������\ɟt����~F��ᖚ��)髿	�?�e7׫0n"��h�e�Օz壟�T:t��n�d��js����ڡ3; ^0
t
clb���r�;I��r}���;׋� ���@:���1^������6y~���"W�a�3����p0��$Pjj�#��3�N�\摸=��[b���	_���}���]��V�����0Z�yȻ[��;�zi�Š��l|n��qK4��9�4K,̑7߾�{,B?��x��^��5�?(�@��݄y��R� ��q��`�cku�q���vn��#��@T����a&(S;n�"UP�p�:H�`Lk���D��XR��ҡ���߹]����NS�|��\���=����F�[5���h}�Q}l)5UL!�\i4�շa�]w0�J�cXojf:eE�w���P�5�
�L ��Ϲ=s7jP���}#�g$F���Dm
;��s:����Ֆ~���l��7b֍YB�.C�s������t^��M�hD��݉�(��D�y(�h�&ܓz�A�����x66{��8�)�!Q���P�Ҷ23�p���gU,����ujS��Ԧ���&djS��Ԧ�;o�|6<ۏ���<���M)�X5Z��w��@��L���G�}��a���/�0Ax*p�SK�x�hv'^��O1�R"j�Le�]�Ű3:U�(��	ll2���j������q>+��@-=~^_0Y�0Y��* �`o��̹q�X�֓�o46�eVҪ	>�PDMG+U��a�16���« ��ǩZL��q͖�Y]3'���#��|�n`���V9&uG"��BHx�n!j�d��y���&�l�}�R���W�+��҃z���Q���Jv�������@0�'T�^��֥ј_2p��� ���	�ac��"��Le�SM{f,����{|���7��$�j*�joz�g�p�%���\T'G�*Q���1�^�՗TA�Y�L4P��'�����_C071�^<��e���5H���$�}�P�a��0�m��ʭ�qܜ���j��#�,�-�~��v�D�tpB���}��C�;`x��nw`���D���ܶDAF*5z��X�[U������(��Ųj�5�9��Fn��� %�1��줄ծ�R͇ I�zp+�����k�2@���̴29Ҿ���b�!����6��̡�~��q=f�BI*Tv���3Y0�t��O��V�b-��H���26��4z�/ʹ�����1�/���ĩQ���׉�<Tk�Ҙ�W'%F�|SK5z��<���Ɠ♁ֵ)���lj%${��Z΁(��H��
�f�G��lc62 �\	�A]�,�̀B>ֈ<I�fG-�4`Z-cX�m� �M�(1�)1Gg �*J#�J5�c��@�#|>S�C��k��z*��� 6-�r.�>{A���w�r��L������ߟe�E�e�<��NL�R���ڏfQ���{o�Pl�� {��"����_�֓����k�p���$�ݳ;��^����c̡S���9��5/s�Ұ�2ǫ=IDvI�	����9R���8l�P��?P� ��q]���,���i<�N��n8w��R>nZ����$\+�����+~�g��Z*���<�G���vb¿��
W�\�;IT��*��*p� �H�<�ːv�=�����j�8�8�5k#��$�b�s��z'߽�V�-R��/�s����������*���v�5�	����#��0�W�$��~oA�)rk0ohEF�P$}@��KUw5j5��m8����W�����<���%�Zڧ������1�����92�G�s�*��|�4Ϧ�5&��.b�"��pE�+FI8�"��C��I��IH-�(�N��[��𽣚�J�g�2�;�U^�	�͗�]]������b"%Uxz�9�$Q�kz�g>]B����F}��9����|��=���3�9�#�â)��2�j��Fx��z�1�JĜ�p'ڟd3���!�b:�sm+�h�b�&�eV���E�Tb�B=j�co�������˿��MmjS��v���MmjS����Ⅴ�\�^��Oa�x� ��z�M��DO���aX�6� 9�g�q_ ;����O���Z �  �D`�C�Z�C�xl�h;�N��4�dY.���Y����j1V^gYG��2~�D#Ȇ�k���<4?��T)��B}�ۢ	�ݐ\@�$�Eld�x��w�L�lN� �Usd�a���%��O���(��0�`z���yA �A�y�d?�y�N�o�˹eA4�N���H�%X^P����R�$o�,���b����MBivG��_4���r�p6�G�d��b�Ԁ��ym8/��<-��j)��P(��6 :N�? 
�?>�SS�����%� �ڰ�>lK�j>�e�y�ʡg�g��\ήh;R�Z#�#��XKM� �&�a騈�
�҄��l����+y����a�]]��#����D�_o�"�yN��jŴ$ @U�N �ڈ��1�f�=�V*�]V�+���|���`�4����� ��A�ȟ~'��@YO>'�d&��}�,�I����g�C1�~ٮB?�	P�Z��FvV���C�U�������v`u�Jp����(� ֫�1p\���&����p�ق�p��9�* #�O��\�eV���c�R�J�p��&\_����<~x�������f���7�;�L#{ a��D3?@��{��;���k^�a\�q<?<=8�\#��{��ai�O�d�9}��TP +�9K��=�	��w;��jV��5s~5���i�N-iP-OrM��A;���Չ�����D93	0ܲl�M������K�R�?����%����bN�; �$0Ü�b'�O���N��e������)�3΅C� ���盐x�+��w�1l8�>[�I�枑Rc�T� �^��UTKV5��bM�5U{��~�)� ,�%/o��o��W��R���Ǉ�V��S�W2[]��ۗ��w�t~�������@�q-�}"����y��U��P�̊�k�*�ˊy��.�cJ�\��FKd/]d|�0l�ŋ�]��ǧ�0��Z�m�~$��#X)����-߳n{�}H�����2TJU�d �*��G�F��v��zǋ��~���"�:s��ՎX5 RdֈZ<��c�D�}�`9
 �;Y�0y��`}ҍcǉ���4�o1/F4((�Sĵ�U�Y�8�����2���9�*BUh��9�쨔NI����*�Z5j����i֚7d�U��y{A���)Q)��.V+*�Ne�S�p,�m͹x}{%�>��o��Fv�p�
��O�ZV�?Q�9��5��/��p��uo�,G�E~,�"|I��N�
�/�����c6��
��IR�,������|��䛯�u��Z��>���$��be�ι6��﨣�@m��ఀ��� Vҽ�-+"�}���C�Xw�G�vFe���a
�6Y�C�2����ta�u��s5K�%�:���i]��]R�k0ߏ���>�ș��{gD,�@��g;F����ߟ���{ .ਇ?�U�g�V*nkz���R�ς�DB�L���|�:��9�U6���Pq�f<0����;
�pьFr-�G�d�|��u>v=�j��jX�.����'�~�cS��Ԧ6�?�6 S��Ԧ6��}ÞM����,
�ǉ�
�� GP16���q�n�a���<��Ša��nP�ϗ��Ff9�/���AF%�	�	�G-�E$K�N����e�ESѢ��)�O�JP�M_�V%Țs�Z��+q�F�!b�@M"�� `��ĭ�tT5��>��W��j<W�_���1�z�]/��K	ؘ��������T �+9]��6���ÊE���ϭ�u0 �fMQ4ھP���Q����V3�l����J�-۸�����n>�1=��h ����o��o���Q����o=Q�,����,��wPy��$:p�-�r�h�Lg�zp#� -� �죁f�����?|֑ Noc�bE,Jȫ�����|���hG0�����;�	���hX�c���$ �ǈ� ��;! �L�F� �T@�tY�LUP�!fUs;H�ȍԧp���Cu}���F��[�����K�֪*�ج>H왚�ן��fU�+A�{.�[fg ��:�zvO?w=�Qi��"@U�(𥯋-��cд{�+@���0o��
�y9�e((�~�Bp��$���3T�O�5��di���T����#��A�8@Gd����j%W�=��ØU�9Xc�Dk�[��jVPm��=�զ�>��g�J�g��7�J��$�,(��(L �q&}XGd�`��,�{� �Sk6V���$&E~�J���9��X#��,�F	���:I,h�hB��kP��*����V���}
0�޼�x�:�����*�rXz{ik�uD�$	��UQ�2�(\)��� V �2������~F7Xx�e�t�p�U�����W�k�?��f�F�3�,Ws�VD�y��?�둱_Q1��6�@��P�1N����B�F{zz�YY0��䂔�B�o�~T��.�w4�c�Z-���e�5	cz�P��&i�8���ǧĀ��2�ven�%��c1����"a� �Z�7�Z�Z�܏�.b�te����b����v�x����g9����f��:�n�Զ�h���g�ВD`)��a��{>�����+.T)����\���,��5���.���<
̓�I�Ũ�T��
�?���>���M�Q}:�1w#��C3Zga~cB�b�[o׼�K�99���g̜:�*5��P���'���.��J���.H��=0���W�al��o-*A`�,/
�򪚓@�þ�4c�!�ZK5��$T	�R��ed*1ǔ����.��J�\�8�;�E%�N./�b������|ߖ�6׸�b]��F�B��>r�_��m���?��n���U�"��e������Yv��m��������XN�5Y��Fb���7��zU��ch�g<N������â��=d%��--�E��3>����k�g�*�X��c�bnWO���r1G�hQ9��MmjS��h2��MmjS�����XY�ب2 <+� 2�1Qˑ���Й>�o60 ���j�J l}F[����6���g'�l����
���'�! �~ؤ�3�7^��J4�|�����Zꀪk�,�����H�"�	_f2 l� ;#x�F.��w &@c�(������#���>�p�U �jQ�M�����VB&�]�j�Hٶ��
�k�4 ���b��V�8lc�1�ˣZ�����J�ĽT�(g�#���m���h;[u��	Q�߱B�א�+V�w�J��A���Z޼~'�_�?���-\3Xg�s%�Я�W��6�m�q��^��ղ){�����7�Y�\�B ���IaQ%Ab�P<�\�m�cf/sT���z`P�/~����_��/�����7�8TR���Џ��`�D[ ͉����B%��p�a��$��D�/��a�C��R�V:�8��h�e�C�O<O4�<c�χ�6>�Җ�̭0R�X)����=��٢�c���܌�����@f%k��e *�"*��O��I6ZeTŵ���H����{��w�{2������x8Z@:*���c
c̃�>����5�|B���t��z��~�s�cd�g
P'�
��pCV�S;�_�3X��Yp��=��j���y�j%��'	�(�9��c%5T!�9F�N�g����ڐ�j��VmI\h����B�R�k��$�h�L8N��z*���f'����KI�5�J|!�-�I�IU�jn�[F�U̰��^��jX'nq���C��U�r;�?�c��d`Auj�!S���XDR��
�(��i�z�����Ȫ�������a��^h��YF�I�0�g.�0��X�ؘ�YG�U���;(������j��W������K#�X���GJWB�_��^?@f�~�f�0��8@�8 �`� jdIF"U:�U��b�𙽁� J��)l��U��h��y^n#��gxo�|r�@Ò�1ܝ*����3�<��s')ܚ����N x���,��r��I�ʸ����Uns����&�׹�r�T��uF�eX���P������=$ݭ����lI����݉�c��Yǵ�l#A����^]q��ɌY5E
�f�y@m��sX�Mb��0�%<��k=l a'$�6�y|Zs��P���J�}��m�?�c�K\@Qj��ڐ����V���j�I�NO4�-	w�?���@�uB�V������XH�ne��<�|��~��x>��H����P�X���T]��6�6_�m����_���D���.uT�����Vx>g���'Ci�A7�.ԕ"�XފYf�����l�KPU��=��1��<�㙡p�j�NL��ּ�D����?���Ԧ6���� ��Ԧ6����[.�n�R�Ԅ���\=��F�~��
/�D"� z��p�u�}g�TǊU�-�� �l��(l��+�;I]eu}-����^�Y����ݩ%���DU
���k�^��w [dW|t�s�L��q	mPE�<@�A#P�Y�B+ �
Z�  ��7or�z(*%�5&��qG��ڬ� �	R�߿��,�gw�2/3y*s�� �`�jq#/����l,����+��Nh��`@v��+	$G��Z���G|=�*@�� x ��M
�e�kq77��U>՝��"�}�����)��_#?��OG��.��A޾}#����<pLm�"*68K	̣!'դ��{��&@C& @\�,ͥD�<�x�G�t�Qz)����{��.�j������ʐ�ާ�Z��o�o������J� 0T <96k�����,�m+I��6��
�c��m4�ǀ�`I�u�㨋u�@�l��P	�����t�0���{7@e�K�i�zo���c��Z��J�3�A�B���QVrd�( �hv@�pAj����f���!��a���!��q���p�����W�J��q�RE����E8�L����D��`'���--�Q%|��Q�cdT� �����<�ԲB�'�����''��A����c����M2���F3�f�C�i/�h�?� ��;�)�*+�~%<�`���NP]�ju���A&ttGd�^[��u�� �L�XCvI�B��DDۣ���u�=�1����$��%��1-��sd��0V�c�X.�\t�bA��G�$�! ������!�M�J�N���Z��r�@�65��	+3'Dx^���^=}�RZ�Ea�B�p��@�<�=��ZI�q.f!��>:�0;��>�h����G��}UdF����W_�{GE�������U�����#���jV�����d�q��Y����H@�$@�?��T�ı��}l�BO[�|3�g����e�r,���:B ����9uAN`}�߹���w�cTDXN����hn���=� ?���\p��39X�.�w9����*�'J��������������jeN�Or^Ou�G��c���2��i���~��s���a��x&����Y��æ
�V Z�:������1�3��V��ғ��F�n��E�{���cn�V�SQ�yҀ8���T�W������.��<IP�θ���gϗ��u��ُ�k�������W�a��T��"�Pu�w�>��tu�l9��:��ik���`4�*�.�C�q�M~;9���o|�F�/�����{Z�$��O-��ĞK- ~0�C4�L�����+����=��*��JMF�A�N3e�ն��ITfa�,F;\|Za(Vf�A=~
ύ�7:@,��Ԧ6��M��M�Ԧ6��M��� �`����>�4`8ljf�U�O����la76TU���f�Ǭ��k�6gw�W�|�?��7T3V�◑�p@��ʱ,n�`�Ѷ�pU��p�U�!�H	.���V�� ���P�<uL�.KFob�����la�n�`*���6s���pd[s�`��SG����h�
<���y�{ɋg�r�\���=���ǘ��P]|�Wr}}'�_���n�Y	K���S�D�y׏�s�I4��o�:��=Aā�7�Fes8�t�Rv(P��4�G�q�e�q���q#��%o�{C@�?��7o�u@O�Dɨ�����@��TK�Z��d�7������lTyw���؈w�Z�x5��O=���߳yN`�K�=T���w{��V sR�bEM����'�����E��^^���܄�oe�����!�/_>���O��ϛǝ�y�� <䡠����AU?x��<<<��$e�x�1�VK���(0����'�����������KB����;%�o�y��Z!�9�v�Z+�q��A|�p�bM�U[�9p�1ÝFZI}�<{���m��w�,����лf�&'�,F����%�����T�Î�$T�k��Nx=�Y�:�B��ZUPLe��_��"�P��:8!�� �$3�6\�V � >��P�����IIjA�f
h��X�H%练�ާ
,�u y���Jȶ�G~X�)d��p�CcP���)�G��8�g������us*\�o[�M��� �AV�UYsN�~)��5�>[1	p1����_��1�^��q��"�O�Z[;C��iIOU�d�`1�nқ��V|�R�k�9⍴B��f�H<�ʫ�
Z���D��sC�ǡs�� -��x��ڵ���IP�q�H��%P������}��)��p�ȏ��=AU�l!9��mX/߼���/(�
�F�Jl��꼡� @I4�T�(I�s|O��a�#K��-�(���&dgd�e�Hv�2c�|R�Tm�:����,$ ��P��Tޅ���X�s8ɉ�s7�2ω�׺*�m�\}qiq�Q��'����+#�]-矅����뎌D�%��Y�����{��z�FI�+�w�+)�g��T�vX�)�Q_(Y��K��Û[pq�E�W�cj�D���3�J�1����N���3�^�)Z��ߩ�5|��Y�OS�<!)ƱH�p�[�âj���")�)��U�$�p�}����b<�x.@uBe#�:�1,/�����r�W�pϦM)	G�.l�3�"{-��W�1���5OG��K�~�,�0t�ĦB`��5���5(�S����+
�e#���>�D��kI�ą���gG=�OH�����%��z�~���-��O�L�s��c�g��VT[a�L�Ɯ-t}q�֑�բ{fǱ%)�١ԁd�$֝Wٌ��Ȳjq���"\��A	���/�3W77�0\�6��Mmjm"@�6��Mmj��ƪ鞁��X��i�����~���7��Օ�˰a��`8����ʙ֙��
jl�E��}��+�f�l�bT.�ծ	Y �I�`��nw���i�16��Y.�d�O��;q�U� ���
WW6�Kl梈���,��*����|�� G�	��3L��%5_-h's����+��l�^P �2d��H�,���J�V�,	0}-��V4��- �6��2	�)n���w6(y�kX�VMD�|�Q���}P�י��{�	|�gs��{F��� ?�ƀ f��{�^��K}:�b~%Y��u��4�H@�{�y�@r9/�%_v[c����5W�y�=|�A^����kJl��Z�gT�[�	��rJ㞶�U"�� �<��B�P�*륤EJ;��ъ[XxE�=7۝�<|=�?ɗ��JWK**`���ˬL��?�B�����˗��}����wo��_���`{j��˱�^��$��n�;s{��ʗ�$	�)X�9BEAϾI������wo�5_�M��U,E �Ľ�7���kS~^2Z�Y5�Uo�M |8�D��.�JǁB�7�>v����Jp q=3y �l6K'����A^�wQ�5�0�$�7�Tϐ�J�,�eI�#���@9T���X�Z0�yX �*i��~����p<q^`-�U��Sox�rvma��نKC:8�@� LüC'��_M�F����1�A�w�mP!��hF�c���B��b�����Y[>�2�e�z��f<H޳ �v$�9ǲ Q1_B�$�F���뫃�<�ReK�w���!��j�H��]��V���dr�Rmݩb��Q_��r��z�-	,'x`�}dMC�X���h���vH��O�rt
�6���4��)� ��V��3�x=^��z�#M�������#�SXw�2��A���}�, ���n�$��w&����E-U'�y�.�ӕf�6>c�=��-	�7 �ێ��u�lI�]恠!}�R�&�n��9��������r���_�7<�e��u��J
��X�����ҳ=z���|��ұ��Ҩ��"q�S���X��p��R�vT���'�gx=޻c�D���dqk,'S�}.	Y_ۜ(�\�>%'=��*�8��u�2��SۿĂ�1��Y~���<���Cz|U@ �u������G� ��ǹ�����*W�W�u�<�� ���NzM1��2��R]�®�,J�iqb7�*���۾;�v�၃�J	R�;�~8���ex&)��U�k�k�-��׿��"��6�/�81KFU}TUL�0�$U�C^'�D�Ԃ�+�,N��x�͠][]4T=X'�o.�������o#3~�[�ZQIR���g)&��0�۔�����c�d���1��8�?��
3�!�mkE=朧����h<��-�y�V��,��:v��b.c}Q���K���w/S��Ԧ6�?�6 S��Ԧ6��[Cu'U�Co�(��'sw6�jkp{{G b�����w$ ���ՑaS�~z��Fm�6�$����:%�9��	���Ҫ����d��]6�x� ".�J{�����Y�,�����\Å����-��VIp�����+�Q����?|j՜ؤC�"�M�n@��}Ͱ\4�g�/�-`�6������}8��,��X^>���՜��o�{M ���oe�������4|��h&K�ҫ��h2C9>q��Z���X;S[, ����ک��������F���62O��,;vG�A-xB#ܔ63�$P=T"�Ӟ��P�@�
q��t���l�L��
́y�=� �r7IԒB��n�4�%��m�պg�
PqY��(;���J�� ��,5�Z�al�j��3���;�C�~�^6��!x�&���P(������ߒ<��Lڞzy��{�o��cMB���ZJNP@�p0����y���U�������<w��Zu[��-f�GeR�P+���<�����t`A�x(�a�ey:���a�2P���t`�+׻0�AI_�Ndʠ ���������B���S���<|�'�:���p�9�Mj��g%o�<
�ꟌpM�������V�"w�kIư��=���j ���q�jE��=�ow�Yr
�5X�rZ�dc�; &`��;9�.�?�zSm1�٬�0	���c�v8��YC��ù=b�G\z�� �@�����!��?Tds��P_!��"T('BO���$#+A�~,�y*��:�.�I�� {��B�ԫ4���h�6���A@�P�Ʀz�6�
�V�^��6ŝ��0e^IGj�#0�hlJ��a�(��8���Dm� �5�$�v#�WBI�N�;�o�R�0����1�5Y8�!AH�a�e v�����Nm�u�AtV'��_����$�>�9l����$w|�k��>�X����~�q��c��v���f��N7k�I_b���J
ƫ�Z�����h���ȝL���Ә�3�bn�X��u%kq/V�-���HL�fOI�/=[L����Xr�)Wm�9�6N\����'/܂����x���E�q�	W��̕i���܆���U�E�jĕ)N�:�j6'z���I�Y',n��	�6�m�|n���R�3�'Xsƣ�0����p������xC1ɫ�}�`t�qAW�*Ts=��f1��N�h�
yA�Ʋ6�+�Ə�� ��?�}��9-1{؞�sH�RoB+԰�����N:�g�߉��jk��<���U^��|�0�bKʆ�	�C:�X����*��������U3���������>�S�h�-��:���G����O�G�D������U���g���ʱ(F�hV��X�a�{ӛ�+�����Y��)s�V�\�bП�\_t���+�D���\~�O(?���i�A����/x7�wa߇��2��MmjS��o2��MmjS��4V�%,�V�B���Qظ_�>��O�LV�+��'�l�a��
Ƞ* Hu<���^˯���|x�V޿+����U�e��r1�w�ҷ;s�$�PEZh%?+ Q�'J*t��5+r�f3�3^`���VW+�Zp��k 86�$aP]�U�DS���+K��p�&��k5��)
РB�����Y��ӊ*lH�wk9����Z����o����+��|��(Y����� �� �6G��<p}@b�i��< '�T�4j%U�2Iz�#��Иy�~�ݠ��xrü�K�����P���x�9������D�yި��U����r!��A��so�ބe�6Jڷ�s�*!V�7�V��p�2QhcƸ�W�"�7�<�9��8G�m@e���YHE�o�ya�2�aI^K�`cV��E\v��:���a}!d�4u�G�UVƳ0N���GU��>-M� C�i'��9��W��-��@a ,��a�T-��$^�;0�7Q���>S�8bH�rZ����P}>��������Pеǵ��f%y�@��f�%i�?�Ք�?�s�}}/�.�����'j]�dA�0� �X�˲]����D�v�㸁r׮�j�$FFH�*E���3+����۫��ƒh��*�z��p�n:��� �����Ų�gi_A�p.�f�ͭ�*�4(]��h���$ c � �SS?l����0���E>����:p��:�M$��12)r��a<�������:I�� a1_J{�����pR۫pL]t��<Bԩ�
�2�
�CR���EJIp�8DJ����B	�;�h�r�v}8~X�A����:�9��@5P�y���3j��gfɠ$#�Z���r��#�t�阁�q�Fb�XI�����VV�k��z��W/>'9z�+f]u�^	�P�|��5m� �������n¼��vL��� ��!Ӽ��g[���A}|/�ߛC�]\ʜ���5>Vz �o/��$���~��X�w�-��f9��de磊���(���5S8��0N�x�xK�3)p��i�]݁���w���2X�X������$��nau�@�F�։�r��#�����:Z��k��2|���v�,?�s�ZiAi��uJ���~�C��X���Ȕ�ɨ�� �J�!��/{c~�k���3Y����0�T܃=R��av�,�s�Z�kU�����u$-:S%�e��u� ��_2�0����Z9�"E�x�5w��Z���"����=�)��D
�2D�ķ�J�Х��cx��:Z��{���T"8�����,�	��7�;L�`5+,���s�6����g���;���W��urIo8������3'��b��c�,,�SMH4���z�ѵWW�������?��\Ӳ/e6�53h�i���`s��t|~�x�Ǻ�ύ�|��ߗ�������G���C���/?�`��싗2��MmjS��o2��MmjS����j$F�86��ą����3�7���ȟ�ٟ�_|�M��+�R�M��o�PX!�}@x�#ӁDț��'���)������:�(�$����!�=����O�Pq�PiT$��h�������sTs�}��@��,(���,�%���vhԖ!��U�E,��g���\��ƪ@�xK��D ���II����Uz��{6������*;l��sK�8~��B������ǵ��D���heuu�iF��x8�Hӊ�,θEq䁢mXEzuf���<6�{�^��Ч�}��kzӓ|ǳ����^CK1�.������Z(��C���/3*��H����}� oT#Gm�υ�9�^��D � ����y
��@v�
, ���	�6]M� �Gd�����������@e����QP�n���q;C g��r^���pܩJ�u,��)�oi>��͖R�u�̨4+R.��x29��6���Ӻ?\J�E8ׂU��F3o��U��da\@o���?�Y͋��&�E�ϩn��'@�)x�67��n�r����i]�~�&8c�6��Q�#{ח���	͜׭�c���㼗n��A����\mM`���0�[ߑ
gJ�*��8/���~3X<�L3�q�O�<�Ir �3xf9+�1�A����{ڴ����b~1�#/�ʀ�DU�p����E��ʬ+�1G��`-Z.2U������!��0>��`$)��b�A����}�ipzv��@㶗mx*�# ��&��/��2��rv;�|���Uٰ�B��l��%���0/{�6�_Ԃ|��TO̓��Uy��
�vך�3fq}�5��5���y��q�`'Eo%�?�~��O�|ꨰ�%9�~4����
�}ǪX�"zP@pm�4��%�jf�w��aQҞ)E��a��n-oØZ�:̱m8�j�I���J���?>>�59�E�8`��@����f����j�%1ķ �6�"�����o��n�y�$���wޅ��E ]W�Wr}u#�YI��û{���j���h�8�y�$���e���F�?����{��I�,9��H�ɒ]-���mb�����_��F�$�0��5��FuOOkUU]U�J:x�Ͻ�YM�łF����ݭ��ODF�U���i���W��d�r{�%��8~6��3^%�l��K���ރH��H������*t�v5���;��Z��2�,�� c>�_C�z���$����<�b
��a��h\���	���������LD�����a�еsL_g~O���$D[��"Ň�{r����nCr�#Y�����B�Y$K��	X�ZU�������*/ا�0����nCU8YL��b�&��yFM��e��(fp���s��q��ס���+}&��hl���"c��J�Ǯ?5;Ad �#���{D����`o�� �Ջ�����xb��)�	�I�qm-ã6k'�E���ȓT(�~筝Y�uk:�A��qؓ*����Aڞ��2��c߂��o��E�?�9� y!��}��Ro��S�l��}�z#�5Ϥ�?]�`�	�^�[�]�L���5��B���@���D���wߑ����m�6�©���������D�N��=�?ǎ���V�oߖ��zK�}�>Ӣ�?��]G'�������І6��폿�І6����ߨW_�R��er4���|G~����7ޔ��sY�X�$��ڪ.ONN�<:u��-�Ve�c?���)_��>}*?��Y��������vJ �oݽͪ���UsV�D��3V�VQE+(<�"�!: obR�����ێ�7�R��A��.�	�nĔ# *W����z̋��@CͱX�I  |[���\��)|�)E�.���bJаП_mVzG�]��B7��}K0 *�N�� �wTd��{�b ���sP�o�i4�mJ,C�U�Ph���͏�n���sU�Ib��:�J}�в@��Q`��X�
�F���(�7R�qN����6/z���^�{ ��ip��h�u^i�3���󥎡|�v-���giHP�cp{i�ٖ��-6<���u!%*��B��v6(���m`*f%XJ(n���4*��(� ���]��}��$
1�`�4re�A&X�&�����*6U��f�Ī);翭c�n3z�ӵ�e}䰭%D���0V�y��3 �c�=P\� ���:C�B�Bx�ޯ���?M`zk,_}���1s F9��J<�����
%^M�~��4���k�}�`@&����,��H���P�-1��ަ�c��2��UÔ��o\��z���걽f���d��.��t��f%��$-�5��/�G-C�u��S��%,܂�Y���moXH�m�B���:�uN���KT�c|�����p�d2�X�Xסh�焹�$E2�o�,�e]�3'�I�8�I���>��z�#W�)�`=Gr�4;�v�Wi�\"؆!�Elm�CB8��]����V�٘^�3[ �	�<��c�s�t�� 4�B�T"P�Vm�_7Ki����ߊm�������dA�q��Z�y�kd�������2=���[������\�����Ug�#(&a����j��y �9�KB+Ō�����d 3{���;2� a䬲��������O�y�������B��W�����ȸ�¦v��7�|N�� ���q�.l���T]^�8��+���b�(ą���^�qH��q��?cYQOBxŇ���!��@�~~Go9u@��s��g��m��˓*�\��W�{�'c<��m��+��A���h��&J�$�x�!�ep��:v���i��d�3,�đ� �Cg��s+&0n���E�;�?W���\d����Xr֊�]l�Yṡa�"���i�yf�&.�Y2�
}U�9�㱻_\U���[Z9��aT�"G�PM�0��y����FɌ����r���W�g|����P{��#��Ae>O���ş�Z��M��r�BS�:*������Ԟ
{9װ>=0�$��9���{��������s���G��h�#�F�_�s�$G�{��W<��M�P(B�D���������s���dhC�І���dhC�І�{o��c�݇���#T�����-y��+�3}����}Y��/���h���6 ��)���B}�/��v��wL��W^}]��я�x����H�K5� ;��y�֪ЃJ�мܛʬ�<�Aa�0?J-�t����a�B/Kg�3"(oAэ���	���Y��di-��q������w<�x�҈��vU��2�Wk�._�݋5@h ���,��rI��l/侒5��I��X�'r�����U���w�d��˵A��DC�]���$>��6v/i+F ��>����$Mr���A�&�;J��پ�=&0K�LV~����=�+�;ȩ�'@@|յI/ݘ��5,@z`�!	q<��aǪ�
��f����R��� P�$�U�����¯z�?%x
|h����Z���*��N	bM ,E�8����l�`�/�ϵv��q�H�e�`�K x�8�L��q�۸���B�P���Mfb�c�1@�.�+d?�̚@��p�N�����J��)3�I�:��no�BE����(�If���˺ Q����	�{~��$&�f���[1o��<E{ȱ�t�}Je�'�a ���Mf��1Y�$?v�]MMb�'_����I �,��G�D��� e��S	V��o#S� �{�sПǜ����#�����z��uW&fU�6ژ ������.�=��V���f����Wv_�-h3A����~�_L��I���pMǝ�}���t#;Q�D�� Ɲ·�
?ڮ�h�z�[aRs�$���V"��έ� �1r�U �1�c怄�W	�.���@?�eu��ȘQй�����*��!+�#��Z��$Z��U��Q�5{�vļ�J�Py(4�\o�_k�ݏ@��lfp6�E������q�5��.�!s�>b�&�}��ݘcXOA��67�/�)�GT�c� ��hL��8���F�ֺׁ�OXĘ���d>_ؘ�\sYz�X�h�f�I����^�>$
 ���\v�h��xU�u<
{�u�|���Ox"���~m����I^^-q��W}���d�!��s?@�ZX�zj�.H��y���@v��l�5}��.�ss��t�#�-k�7O��y
d<�9�GF:��Ơko�ՔUo���Z���Y��\�Y(Pl�Z�s�Y ^�I�=#�����S{v����~SA����'P�F�rIB�Nz~x���-�+�n�[�C�����xB�Y?��s�����k��Y'�'ngk�I�r����`�5�}�G�.V1N�أ���Bm�G{�'x� !jYs��{A��@(�B�<���|����	2����~G����YD��V��o����Mg�h�3W��STd2���N�(�CW���2c��}��/kf�a�&r��9==5E������==�?׹"F����%lP]Q�oP|���dhC�І���dhC�І���v~~K~��Q�~������C��|�\^]�n�!���^^^ʳ痬�|��9>6P���L~��?��/�s�ݧ���>�=�3��k�n7�٬��s5�y���Ji���lP�j�*��}�h����P�
ߙ�?3�h4R2Lڈ  r�Np�V-33����V-׎:����A�e��"� B5:^N�������fI�j�����'O�Һ���X��	�/�[����J&��A�9C&:�e  @>Yn�k3�f�{kAt�������E@�=� ����*�$�=����UM�ρ�O�����0i�V�F�l�  �w���Ug�?�&�>��!�s�C��f��V&�����P�t�S�4��� cO8�"2k2�ȯ��d@$Um���!
��5����S�v�&��@�`\�����樑��p-:�J�%I'�F�y��01 ��x��VR h�����,Ce-��nK����Lbc@m���
b�!�1v�>�� ��h�WJ��� �^� ;�я�Y�x/~|md�勁�!�V��X��rۃ�ޒ�
.���)hX����ݎU�;��2J����A�7|�1n9~����E流�)p-��c���5S��kѢ[��@�e�$��Põ�ޫcb�H�f<.e[����*ǈ����5�z/���A�Nז�1��L�C�T��	��P���7�\�qb
 ��}b�<"�GC��Vh������]�L�j�J�����#(AR(tm=N �$hj�W����\�Ǉ%W[�����F���S�o���[(���H?3�{E��dbפ�2���i-�����1C5�Y[��C�A��Vu����Y\�8�$��F��,|����Y*��kY�X����[�R�}�^mx� ��d�|��g�㹎Ǖ�|��lz@Dp,YC�z��Hu�>���&4X%a���r�s�zŹ��;q!�����7�8�=逆s�����;��c�z>=�� ��P�@��Ƹ'j�ldĶ_C�5`�t��?�@�^�e[F=��?8�6x��!��� �ǯ��?�i�7p��_�x~9!��� �'0��?�W���#�+�*½�k�'A| �||�'D�ߓw.�{t?ݹ�#C�; ~mm�M�Ŝ1wo�A���H¶������a����OS��Z2�����\�b�/�˃9�`٘r|�0���$�C���'T�H�E�A��[�n��E�D�\ϸ�@��<7}Ngsi`�E(�������ҭ�FNwޙ�e��S&8匷��@�X�J���l��Z_C�Lk>#˿���g׸4�cGv47�S`x�$����+����:R��e���+"�3�|��q~����K�Ŵ�TF��4(*h�g����t�<�����,K�+UG�a��a5AV|@%�gIO�umۏ������~Lu��ye� z�8'�o��n���󏑮x�����_���`]�І6���q�� �І6���Aڻ?�����_�>�}�Uq��ŋ��Jj}9ެ���Y���y��;�.W|a�{����3y��S�͏��ޓ����ܿ��/��@��ɷ�������x����p�+�j��gq�v
�.$�4T��ڲ�Y��P��Z�37@Ħ�,|�$��a煪�в( �bʩ9�uA��4�r�-A�PQ`�2����1���b���D��c� >~�\Vˍ�G����d@��bxqy��ͳ� `��%A\:������;��s-"�~Ҡ?	 �j_�ڠk���t��pU�Gh��e'�x���H��΅��h�-d�*;�7�AD~V���e�o�<�}ɛ<�Yi
�>����W��9x�_�	r����Z�4`��1 

�Vu%�e�(���|�؂1�~g�/�^�C�U���?_��z���s|åm*z�;�RͪF���X�� ���T� 7U����``.>�4��:6��Vn � �1������N�>�u	A]S��F�z��1��J�I��a5��A�8+(�;�@[��4!t�Jf ���O�&�4�X�Vj���|0��t�
�;l.X�l8kcfy��c<b5�e*Բ��w��X�Odc�%@.z��Vъ�u�Rg#�g	��I�U�~s�+ �F��0��GN�v�@x�p���K����� P�<	�R���z��Q8�D��h��N�:���*�3��:�wUi�h��m�� *���U!q��P�z�
"���T��:M;N}�H�>�L�,B�ǝ����-쳄r�`o�1�G;�4& ��3X}��5t�CY,��L&e�x�׉PmXD�6ES�W0����2�-]�_ϑ����4t�9V�c�YiL�N ���$C;��S"��F�e�u�'�3L�ƅ��X���Lt=�NgR�5����d6�@o|[v=�����U]�P�G�_]�벑x�o�b��ʲ������5bY�^�"�k�U��pvz*���ܬ��ڬ�f���)�犱O5��תb&�\�c���O4����IodVJX���.��A"ɩr������O5����l��'�����a��:����hɩ�H��X���������	o��W��T����}�g��bΙ��Aު���a�2����o_P�x�L�=A����U-���Ʃ��� ���%-�����c�bl�$��(s� 6gq�����e{,��������T��b�ܟGTtDV�����)���<p����}��鸞-H����"�,�>�wv6&H�����8�
$O�3�'L�V�e���Ĉ�^�X�אa�5�0,ݩ��nM�j���"�΅�	�?J]ҰB�|�[�:��U��oH���c���s�qd2Ԑ#��-rr4��Ŝ�텮������9s]�`_�qh*X�C�yW�Z3v�h����$ޡ�Ø�b탚�J��sa���#Y���_S����F��8���k;o��xP`��Y�i��3�{&Lb{NA������_�}}Gx�w���mhC�i2��mhC��7��0M'�7 y��Ӟ&J�݊��J���S�����ן&�O���Q��D�!l	\���W_ʷO����뿖�^}C&S�?yU�g���Nf�BN��,����1��C��)��t �V�@����m2 ��'F� ^��B�[�&��e��ZDfZ��%@�>��� X�\_\>��1޷7�-�͈���`<E�4,�ZS>𚒈��ȑll/� î�/d�4���J�z�� ��D?z*��F_l'��\���@�i�# ��A������
S֦��
�D�ڷ�s�O�ڮ	Z�O�>��n�F��h��b�;Z�5�Y`X�
�Zt ��o����`$���{��N����7�߅3�����K*S���V��C�
��uXU%����8�#2�ʑ:t���Ѭ����e��8%�H_�6�7O�X�0�+}E���9>d�#�:*��x,E(���O���J:�dYȶ�GV�L��Y>
!���=���d�<�yt�߬��|�lc?����)	\��E@�i�7A7�C� ���9�? _��@!�Y���,w$fujT@l9>P�w�U��'Ͳ)A^T�o�ҍ��V[�}��v�bn B�+�8�#��7� ��%������'1���>s#r� o�B��U�Z�rL�~n���Mo��?ü��#�}}}C��V�
���T��JZ�EF��˧!�[�/�8�!pA�� �`c<���iǘ�J��+ײ}/צ�Y�$��c���]&]\S-�Ҳ��*Bhj0�2�J�1��Ɣ,��Hw4��UT�����\��cY�X��;f�̴z�"�]d%��6�y�d��#�R�d������|���׸C�?\�������^8[�p��DB؅.�}�*Gb�w��Z�_^蚸�X��3�Iص�h��M�q��lu���ֈ�$1�*)��z\%�
k����أ f��T+��I+G�G��+��X���xP[b\����8v��E�����m���I ��b�D˒)o1e[D��U��Tad���oK��R��w���~��z�s��D_M�=Pث7�/���I��x�ï�������%A��>K�s���/�?������xh��!p�D���q��^5��,�^�f�#qܫ[�Bm����60[G�^�"��n˝�_�"o$��g�Z��Ϡ��8.S��AM��dR�lMc�E{�#�+ e;��D�\7�~&��PE�$6|_�Yc:���~�3����ux~�,��"�?�by�C<��=��ԓ�[�j��b�Y�v���dDz�<��F�XPia��"�H8�u=0�
<�����4�-C�˲��'P�g��֌|$)k>���龫ϋ(T��d:!)�g��Z���u�����麊J/(q�X[��{����9v�<*M����r���u��1�>��
!./�Q	<�=n:��s(Z����H�(X�>����}��ߗ!dhC���t�@�mhC�������Y}ָ L����ꫯ�o��o�>��� �		�j�8����@�@�=.�~���������t>����C�ce��bq$�t��^��M<N����Ƌ�y�����{l�����q�� `gŚ?}����B�Y,�� p*���8l| ��^��H ��>ɔ-*��(%�[��_F�
G	�46EF�0I�λ�|��l2�:�YIyqu-���/�P�eIK���Xn7[�^����ժ�� ��
�� �֑9� A�H-���PqZ5�>"$���Q���̮ t���hY��t��;}�*	G^�z�EX�9hΞI̧��M�X u��p>��pT����R�����@��'ŋ�D�/�̀���q2a�vK&��6�f�CyJ�/���GV�ѫb��t����o����<xp_N'�.0R��bޔ?/�����^SPr$5e��D��,�"����Z.&Hh�-�P � &�4 ��F������~A�U��I��<�[W��}�H�,�i�{౨��1�����o ˃��3A��H��L T#ϥ1A��R]��a��db���|̳���9�
tV[�2�����T9V�;b��$�e 9����=�Tf�W	2@~Y�L�v� V�:�/��TV1 �u�����ɑ�����j�$�6/�R<D�D&p�	��nyLX�����ϜE	���˂��l4�*g�t���d�|Ap��1��Z�CM7B�,~֮�b����6~(�0�AJ�	+�+RpPe4��1�d�X�f>�H�������A��Q6�\?��
��XY ��G�s]K-�$���_e8�~~����
��3*4l����ga��}�`�Y�H��0�1l|Ȳ����������\��	����F��I��A�22P�	�qe���,��77+�]gyD˼�i�T"�kӺ�*Aj�L�����B�=��/5z�Wr~:�ѓr-3�@zb�^]_�<@�B1������:T%�8*)����Ĝ�^)E�-�l�	i��g�T~=�ρ �����ȓ�Y�y���uH���==��������\F��l�7֧��r��_�Ҙ
��q�U�#Hj����Ω"�n�|ks3�\�F��uHW����][П-̲1m�<�Sso8_A���/����a�,�J����ň{ ����,Nz5��_B�Pyӑ(�\?�Te	SۋH���a1�a��:��(�0�f,a�X�8�_�̆,��F2��hN[5�@B��=�$��UT��s'	$��0g~���-�(ړG$�t?���e1q�.��Z�h]���Ʋ�J�J�k#7���#Z3d����
6�S��C?��S�1՘ ,��}(�`7L�P����oY�Yp����dA�d�3q?hn9s6N۪0�de��j����dA�PLә�$�����z\UI��S�Ж}xy�\>�����cZ㞜����}��g��1�n�M$սn<�8U�kF��3������mhCڟ^��mhC���f �_���� �1^���[��/~)_���K̩��0`��$���-ְ� pEO���W������۴�B="|����/S�68],��j �_�C{	c����A�T�0N�+k����U�\��a㨄�:T�]�\J�/x�����hd�^��f�S�{��P����r�ǳ�j!��5�����E P���q�G���*���|~kTA߃=��o-�<͂�#U��G[_����_�	Gv	_b��o��j�*nc����
vZ;z�B%'����	�#w�e  �P��c��1��g���	�`W+�
��J��YY0k����5RG.��1@�`DdJ�rTE���e�c�E��ↁ�z��R�&��	�$�K�G���ү������bt.VX�E-�|�H>�Ϭ�^��f����_��o�YP�v��|lX5m F�L��L���J��Id�����S��j��8�@��·�J̬!�iY01�QM�/�B�M�P��JY\�� %�����wĹ���P�4�#�B:վ ��D15�y��^�P�� /���F�*m�rJ������Q�ܑ�B�*�e�g��u�}r6��,q��;���܈���?�A��|�;ֵkڑ��>B^K�,�ЬF��F��8`4uA��r9�I�n8�����dS#Jv�S\�S�� ��	��ˮ�> ��2"�!�(�=���̧h�9�9�Jn=.�J`cuCm# ,d��<A����Ӷ����?3���juЭ`���JX���Jt|\��-7[�����^�&�b$��|!��u����:U����*��oP	�N�o���,�"S�խ����w6K:62w��r�ݮ�Vѯ��(��1�Z�gK����j�M`E�d��n	&�j0վ)J�וe(�.�T�#���R��z0�2y����a����!W	럳����4m���Pw�Jz4�}u��V����9�$�Z���a��yN��#k
��%����cͮ��r<yB��8n-�+[�Y����]O�xb��� @�U�';��߷��V^9�m��q�E���C{���r# 6��_���!bkW�5=y�grԦ�C�u��>��P�a�A,��g��$hZ��e
-{�
>
S$U�n��{�@���+�Z��j$����r�L�hP�=�I�M�S	Bm���$w@��Iխ����lvGAh��X��ن����ώP��Y�q��`��VL���Z������8v$J��R[ˍ �����7T�:�%h������p!�9R��u��I�䠉�s����#��Q��w
��2�R����F���@P|�=4�mo�&:>t}��k�.�9w�-��9�J�������vL�.-�Յ�h��i Gǋ����0������y��s�����2r=����)���:#���5��ry%���C��������N.�_��>;?���Ux��y�Ϻ�;Q|�k���w������ݣ����/��+��І6���O��І6����^{�a�ߨzhA��3�L�/����)ִ�<ċ1���^ܾ��k���������ـ�  ŨRm�F����x�"0�j�|K`/�qY�_�-�ݴo(�TzL������驜���x>sUkS�u��������WWW�]������-�fTa|�����ݿ������D�����,W+i:x�/�EoB�'�md����LPl�wO_R'��k��*,� ��H6�r$�"�h&��J���(��jl6�  ��
o��.-'E�A�q�*Q��m	� [�P�!�h��5�`WW�P���fI`���&}�Mb�3i|�R���J�W,� u�u�,��g?��V��Uģ���WFz5���)+��3���e� D'���2C�}<�b��d٘����[/�ZcdES#+F���B7�b#U��:v#BRX� ��6�]JD����+��|�EL���O?������� f��Bo�A{��Я�����k۝�q������35P��a-�,c~�R�T�#�d3Y����s��z�Z��\��`x*�Rm�!9�O�޽�d~|X��Z�so�oFiP�$��=x���E���?R 2�'�YX��Jڂ�Y�x�(c&�̈ �h@�@O�����~�އͶ�ƑB��/��(v����}�f�/ޙ��B��l�k�}����s��*��u�[%�)  ��)u�ԭ��!\k˔�Vv���#��s ;P���;<֓'OH:�T�9�f�9��]�s�,�n�-]$�ٔ�.�X&�D��ڮ|س^�����SZ��Ph��"틢�nC �f14
"Gd�Q����cӦJ>fk�7+��'���L���,�MA���򏜒��7��nF���|�#źp��bBo*Ġ�⚤} t��e����z�5���k��SA�ǻA~�a��T�E������6M�9'����$��y��:��w'��/r��ҭ[����,&�KS���~�L�R#PZ���R��̎%�}��*��Syp���C,W���7�d���d`��tI���r=��RAT�4DVF;�X˲D�޽�c��ujI ��"� �vW�y�>u\�IC@�������g�����d|��Hz�`� !���!�ucU�T?�>�uOp���ГX�Ŏ�!(�'g:V�{rf��-�y/���͒�G!��|6����]?��g�͎s�=I2�F�|ݺ� �%�o+e�c�V��Z!r�Iۓ h���H�Af�4�|�H��K폎�s�$�{a'ɬ�瓐H���M�	K � q���9�f�Pg�$h�d'���l�u�[e��w.d�8(���V�n��q�똭e9I8o��PXx���R^~�}n���QKKq����5uX�	�^ƌ�wP��T�敵1�����A���ϐ����Z 10!9�:��s��R���G���	��A��(��g@�k���c��h�U�^��l6C*b��d �f�f�3�:8&��u��t6��\�b��s�x�7����3�6Ts�z a��A�85�812���&tJl�M�	��V��mf�[Ŕ$x��#�ɒ2��#��!�޿��J�<�	��y��</,$^??/M&�������*���4('��Ho��}>�1�����n��~(�A���&E��7�5b:3��ju-~�k�/�r��=���>�L��/!��\<y���뵮t�l�>m:�X`zb�Ou�}��鏾�B>��S�5��{�<��mhCڟF��mhC��M���F_�Q�W9[�荅��Y5�/� T�J_��#����y��˘�J"N����ˇ(���WB��v$-	�������
�\0��VO�I�]��('b �d�����R����f�~>@�㓅,}!���|1f��]}�;>�%��1����
�M������ų�|A��q�/ɛ�J��W���+�R&(���u��
]5+^�aI�#Z�Ja@avR-)�x�����b�n1�"�/�U��$?RGB�7�۫=B��$�`t�G��;�\#m���J��� ���<���Pu���J�H�A	�nD��	�=go�jː�2@��Z��Aظ^H ZE��0�%�|.�e\ $����,�l.w��ɧ�/]���z�WG �٬V4v�zAϖ ��Q�%�qß<�j�6�Hx�G����ۖky���6�:o��]Gd�
��d�|x-6<*?Yl
 #q�c*Ψ��y7:��6fE�����y��d�Z�7�|I���o�_vڟ��`%�VQ�t4�7>�UW 9`c�
�ƅX7�Y�p~�ne]�"?uJ��R�� rh =Y���x��12�g	\8	�m^���y ~q|�����?���>1�l^V��$g���n
�D��
 ��JȚ�-���Cq�BV�5B��5�*�誳���l�W�o@d8���j,�*�y�r�M��K���
a�����teEлq�c��_�Q�S�!혀�t<�><�=��H��;�=�Ŏ�� �<p�,��,ި�	�

D�.-W#��V�O�.�������sL��^�J�1�I�<,�`_�@ƺ�U�t5��k= �QF��܈$ ]7���ju��E�
��Qm��	�@�ҁw���D?����OPW�YĦ�K�3��F�k'5l� ��1������rC6L� �t���h!���}����s�*�T��
fJ���UL����If�1JJ�T���%ԏ Fνi7\'N�n�b��b�3k3��J��� ��c}�s]*Za|%�H 1�	'& ��X�u,q���ʏn2e.F��8Q���w�[y����ņY&�ٔJ��z`(v�|��[���x	E{����/��o�9�������?�*���<ogd�������{�%�"�2K]�tC2�,w���d�?���v�m䂿�{�Sh����*�x�k ������p=�_�(�yY��c$�U�,��4ퟁ�46%�t:�g�S��(��t\"�,��b���^U�Ό��gY�DЯSx�j�s��$�%_؄��oUo��R������Rʻ�SKٚaa� �� ��1��g<���r�綹�	�n�$�p���ku�T������7*niw�r�maE���ʲ��3Н���CI'��*S�d����Y7bO��J{��i��5������xv|<��!��}��=a��8����I��<w^�dl*��u��j
�x�o>����	gX&B-�1��ubŘ>�����NCG����=�Vƣ��V觝�( ������'�Fθw��)���"f~U�ge�G$��{�g�"ח����6�$��mhC�����@�mhC��~�m�.Y��
R�R�0Eo׀C�4�u>��Y���QT1�EE�蝾dn��L�1UǓ������ޏ~ ��U� �G����֔ ���	�@ .�Y���*HX�l�\��6Q��Jiؠd<�L�󉜜�P�ċ�Ї�\T������2���7=:��ba7 VW�o�O��gr���fu-�������I�*@�aЇH�AO;�!�/�EI �� |�|/-�V��S(:��,s��@8'��81��� b�6*���@�$P��	I%4�����.�0�֓&:{�`�څ$��M���~@'���#�(�a�^@�/ʲ� ���\������M��v�!��p0�!�>A�*^����=�>Ķ! B�	 ��u
�G�3<��N�ߒ��L��LV����XV@��0���tBK&x| G _�H�Y�?���B	�4��؍R̔U���~\�\��8g
w���@#id�G6�d<�9*�C�nr��B ����#-�V[W��*c�ozO��1����{ �_zI�~��he��<���������}(ϟ}K���|����sy�7�/��ʻ?��P,A]���U�>�����^���ޒƪ�X4`Ҫ�M��`�4kg3��ֺ5r��iҐ��*�9,Q��}�,3X�
"b��u�m�qb!��=��,�p\do8p*6�IG�%�	�l�;�� 0��e6��g�X�
���7�hh�Jv1�줂�Ȇ���JX�13#��m�-׆�2R SŠ�ڂ��w�z�}��M��*1s^��$�o��d1�}Pi6'f��9k �����#���q�rj���l-��<��e,4n�� �eX��;�{��Q���Ղ�Aϭܖ\Ǚ�2���׶ٺ���&$���2#
��Q���-I��;�5��{�	�����9X,ci���(�tM�{v,��Ļ�����ȗK�O���E���qgz_F��m�sw�oEݚ��[Q��8qKB�w�m-����a�9�{����m�Lto�B#�0&}�6����@�˝�}	IWe�S���r��|��[ހ�Z�㬗6'��ry�*k�yUZ�"���z^N�'�;+���?Pj?��?���� p�	Fj�Mf|�-��k,�(ry��0���c�����R��"v�Z{�B\��>�����z�œ*}��o=w�M-���Ն�����	�B�� �I6� ҜH�,��	�ޱs�D\;�օ����֊��k��TL���O���l���������o(y�|��Çrv~���nWp�Ş�)q�
;=���2>�q�ca]��_�@X{~�[�1��*����2G�	L�g��̇0�ٳ��k ɠ~�55\��_
,��c�hq�B
("B*^l�!�X���{b,
���&tKg������\���hyE"+��1eR�,��_IH��zeGd��?pŕ}5�-�#r{��U��G#'@�`�[�'�,��nߊ���N�oZ��.��}.�;,�J��jK�
Ea�����l1�[�FGG|���Dt�� 9��Wrus#덎�nc�ץ�����u������/>��?����}�P�!�+T޴f���B�����%�������G����d�}��o��}�%�:l_$��6��mh�m @�6��mh�������u/�hxɾ{�����rs}��TX� �{2��P+����[r��}9�u[������`�gid�H_��;)����%9�B�L�g�=G6Z�f�6@�F7���јvG.�Ã�ݚ�FC�;�˚�z��m�JK����bx{�����ɻ?H�_��!������_����%c�jT������B�D�?}��Oy}��#���dbU�̀ ȝ$}�i�<���A����{���	����57olx]'���R��$N��>�.������w�� �񺻖`-��-��#�<���ūwƕ��L�x��ڪ�y�[��7���\(r��[��e �X�a@�K	�*��,Z�x~-O�<�#� �����B�s[�b��MH ��T-3�8��B��&�8l�h6�[ggR-r��:���@[�QHp#ٙJ��Í�%��O�����ǡ'9��A��������6k�i�f]��?�{�@hX�T��jzq4�;���k������oX��2�i�L>��m����#�~���V7$:�~���{?$�x��Kr~~� ]��\nB�G]$�����8�
�Ћ߃��}.�܇�c� 4��#g9��xg����	:O��4�e~�Z�{�؅�V��w�!��� ���s�q�~,�3,8~	$�
o�#��>e�yFm h"�7�Z����|��'3Z?���.�Fx���|),�:1u,�u�X&��r� �_��U�cdƌ���ۉ��n�
m�eN�2(���t�5���	%3�t}��_����)t@��{�����<HY*q"#X`�U��C��lM6;"�� �	�f�¶�
�� �� p���W�(�V�ul9%�p�R����Jv덩;t�m�+��� uk�1�MA�U����pF8ܬ���J����1���:������l.�INPU皮��I� �1o����G��j�c���"K7�d��/�li��{�9�.j}sC����kC������;/|�xl69�l&�9	��)�*��a�T���1��^�F��Y�qP�fl��X�w̫��3t�@��*q��1?�[6�Ƽ�;]�cG0�iE���)�(+��Fhz��cs ��`J��[/�~��D	�8t�Fay(y������U�u���'�#?l.n��c���}�z��#8#��i�Iw}��?���ײ�h�+V�}@����W�/K^3�o_�O�@}JB������,+&���vOΆ����ɉ��/�l~�y(rHy!Bԫ��X��1���A%*�*3+���ГH���V�AL����%\{�3;F<X�aLdY@{���{��Ϟ��$���3�R�{I밐k��"�Q���+R�
 n���w ��� u��AA�}������WI��q�Tn����찔�F��}���bz�4���6uM�F�@�ZM�����t��ji*��YE<w�ܑs]��5�c�n�l6'v��� G.��'�����W�Z��z%c؏6�@���Ϧ2]����Z�/.i�WT-�E��f>Mˠz�O����`_8m�F������Ib�(�gn]_p�@�v2˦\'w�-3��>��y�֛2��mhC��i2��mhC��5x4�U^��Ϩ�m
�.�e�޽{�ӟ���,��V�F���I,G��rr~��S�{:?"Ț�0��� X}X�-���[�PuT�zf���B%YD��>�~җ���3��'��jy�QP����#\�/����_@Q=rrd�G��\��DA�7�zK�ώ�ڎ�X��~)O//�+��;H��K�	b�� �C����I
���!�W��ys}㈎�VhE��v� �z�=X�*%�s���b�j\عU`"ׁ���a �,j 䡢�Ӻ���ٜ ��ײ�2��N�Z#�+�+����(*�> 5`�#ɅJ?���{���@��_��oj	�1��>I�R��Q�)����_~����w��B��٬�H''�r糧r��mZ�Ay��^V�׭�*̧��X���K2����BK��6 o��P��6��J�ոV-�v��-�]��ua�d�$tV(!�6��G� ������,@��g�r|tJ�d�+��� �~�g�˃�_�G���\]]��x��7��÷d2�Һ�``����r�
��|"p�1��١��BL�����-�J�#?j�V��}���@�K�U��q��/>�����1mQ3��t�����Z�V����ȭ�� i"+��d ���>�@��)���fWt]l@rQJ��SǠk���
�������@��ӱ�����γ6b�)`0��21�sǁy9�L.t�S���1I�����Ɍ�����y[�|������=֩�vq�LƦʃ~�\ X��Y��5֛�T��k��&�~d#c��E��	{�زyb����ZɃ�������3�����[Xnt>��l����7K(�`S3�H�d�N������d<���z��>��T!#�XיB��A��^�&5�E��C��\B�7��|2�騗L�a���GO�˵���GӅ�u^�a½/�Vl�cAVZ`tI� ����:��fA�'ֱ����i�q3�Z6r.�?Nq�U0n`;*�4/o���R��+�V=�݂�[9uΈ��w0}9�1Ƨ�Ǵ�D.�) �5T-s>X�llnq/cվ+PpĘYF�t�(I�y�)�8�y��2��Ĉ�]_�`ꦲ'I<��sA�Z�Iڞ�p��X�m��ZĈ��)�#��r�q>�VN�Y^N0��� �\�����W�x���Y�;�i�#s}��Eum@w�v�
9Y:_���:PB���iC��?Pq2Oj�}�����n�z�G����s_f~O�ӵ�����0	�$�\�����?8���e��I`�+��3����M��qbc�X�[G,Nm��Qd��Y�+.H,ǣ���!-�:�j�s�A�=_d���L�}k�O�a:.�q!��=��\_H��X�#�e���T��GXߨȤ�4R ��*$��W��`�r,a�L���+���
%3���\rvv���w��W_��^{M�+�r?d�9
3Ĕ�-	�Щ�wrss%_}��|��G������_���s�F
X���2ئ�����X��s����|iWT[�#<�`���m)��l<��k�
j�w�Ĝ!�� (&ia��8�T�xu&�+��-�hQvsuMS O��Z�?xE�6��mh�m @�6��mh��ݣ'r�;��d7)��Pa������|1c���v����X��3 � |�w����2p֝�3�+_�����xo��pN4(>�M ��(d%�t�0�(M a/� F���U�����c��2�z�r�r��p����xy��_2���B�{�m������o�{�p�#�z�/�w�ܢw���I�Q<�7^yU�x�E_}E/q\ 5&)���5=������b���(�F��1��� c���k2P�<�Y�)��;tU���f �H2 6;�����r<��<>σR#��6$-|3K��j	#H:�S!�e�'�V͒Â�wRn� �	�[,���WN:{!g偏��Z˯���^��^od�/��xC����ᛯ�k��,��� ��K�79�1�xc"�7�+�sy��)� ���A�1�M�WF p.d{��[� �Ep.-O���}�[�n*u�
]�tb���9+菏T�NE,����?TWN�A~�-j	Խ��^뫯r,�MF��IV���:ߚ��\W�=[S�ތ1+�SzV����Ə z�LJz�����k�;�p�B�a��<��M(���*x1��ܪ�Q�>�M�τ<�=B��� P�W�s�u9�ή%m`c�s`q���1r}�sAleT�`��G��1������A��q�M��yܣ��VK���<� �h� -Tr#��	����P�?{.��,���]��H{ �a��uǸu�\����Rj6b��^� �n	>��of}����7 �@�²eg�ՓiF�7�Lea$V�ߩCp-���H�Y�H!(Y�<ُ�����)!�}�/Mfc�K�g���Z� ���u{����G���sSUM��l��H���[�t^�Z��Q^I�t��}FJ��Y����\�f�W�=��~���Ȟ4&0�����f˜ ����5�&���2�<��ʡ��{�l�Hΰ��HB�Hn*�q��;a|�Q�`��a� � �{k=��uc~�)K[c���^=�X��F��"�����nKf����Z�a�U;�S�c�JG��b���So�g���u�[Z������	I|n{U���@px���[]����T��e'�ˡ]��<�娙��4	w*��mN��ī5<���q���?۫	��E�*�^g�W�xK�(j��uk����  ��IDATI�V�{�af'Բ��ۇa4z�Ȣ��ֽ�tO2֕ȅ��$jz��Wι���7̘��Щz]�݃�T(:���n�,�m]��^��s����x����x�"����Շ�;=�CŶ'ͨ�h��$��"�sA|HkIn\uf����Օ/������%�EZ� ٛ�a��<Ӧ���IbjP��{Tz4�!���b��ƍ͈���[�z�̏�w�h��7��3T���ݿ{��iIx8XF����GL���ѿ�����O.ޗ�>�X~��/��o���O��'���gٜ�3ҽ5s�!���b��R辰����n %f�}�6fa�sŭE_C�g�۳#*���8^����"B�'IF)�@��>PD�����?�L}�5��_��%������3]�ndhC�І���dhC�І�o���3��Az������٩�t���.0v�A�)����v�|�� �2�����a�{vBg(%@A}���j2  �D�P�];����NH ��@	�����P���Up I�b��F_Ʋ�`�^o.V���w��y��m9=>��˧���c���ohp���z~�ӹ��?���j.�ϟ�v���my����͇��wO����3}�$�}M�D�,�}Ȥ�.{���Ug6�������k-
��8:���w����]H߷���t��U���:��Aoe�@Q[�z/'#` h�+u�c�/���T\�T�����*U�e7.p�9_*x�(��?����w����d�q���;��ʏ�C9�[�{r�ֹ�Gf�����hJ�fp?I�ŉe��z��{g�	�X�f�D�	Y+P!��1n��3�����`���~��0A	�w`!���J��.D`2H��"��=�:��T��;3X�jv9I�$oI����)�� ���%eS��v�U�Tq>��D7Z�G؃�^�a�ߤ�b�Uc�
�Y�*�1��f���eX���vWv=��T�z�͚�8t���(��Ʋw0�j�{9f~�\C�����W��YA�n���Y5��=�h+%����+��@�\Ǳ��跞��Pb��(%�VWf�U9+8kI@ �����e	ϩ�u,���"r?:�����RM,��Ƞ9=3�% j�W�d2��"e:��b~lV�@�P��=��2�����k �77��]om\[���/;�7b�Z�=�k�C�B=��?��)�Q�c���x|�e}X���JyT)o�z״lBh0��άQ�>���2�~�F;5��gP���S��|*6KYA1!#4�!d�dzMWP���յ�c@�����E�):h'����ϡ�"��P2�R9vDc��Wa/ �I�3���v�� ���	2R�e#,��bl񈤊07\BeP[$4;0���z̳�1g�С��^���ľ�mA��|=;?����9I6�+W��)�l/�6t�^G=�>̘S�{��gr��	Oj������Q���=��3>�H6U�_[�����{��CD���M#�bZ�ct�(�BX�4\�(�b˞���u�F(t���u����Z�	�9"��%vʸ�����Я7U����?��)+�>������MZDvNM��q��)L6�,�T���T��,
����V�c�s���a�$���n�Ĝ���_3æ��g#XS%��Z�[�d[��>�t�O#��=�`�B*�ѣ���Re�#�G�L�c���s{]����-b�aAχ�'�4�l����=a׸\3���aLMk�7NM�I�_];£�0���o��s�Y�kn�M�!F:n`Qg��"\O�Ҫ���V��-���~*?���7^��~cS~�7�s�v���<Hn����q�������/��˯�L5��_ˇ�����?�\�Y��[���h�ڰh	�u�Ι��z���+]�r�R>w+���M��:V�?��O��ݗ�����̏NhՊ羫�+�1�G�pEn
��B��'�9~����7������D�6��mh�m @�6��mh�����$LG򪾌�;H�o诏�y�P�ŷ՗�(�K�� �`i��9�Xhm�.PX��-�:���F��4eC@w�)�2V�B�n��-�jJf
{���W ����i�%}�&3	�� 9|�8*g	8Dt�&���Z7{�	�^������s��������<�{�A�_�<z��\/����oȢ� |�
�c{i��6����D�߿K��^3�cV��� ���fs�W�)^��B�a��cly�3��
�lL@�h�H X�Y]y�
�w�B��}&��@T3 �y͎d安�w�O � Z���u�a��X��/�kV����S��þ(rVM�m�����)D"ޫ,�X�י�8\�e2�1�`|S�}������S���]f���Yg�q���"G<�ZF���U{��X����ٔ���ԃ9v��0v�!�jC����\Z��F��;��ٓ�TQl�E�s@oV5�\:N%@�����bcY7�:c��v$A��u����F�������8�**\��fz� Ʈ�`�>�s.A�Fd6]���ePE
���jV����g� � 6C>P��+v걈Ұr�mײY�G�Un���1%��Jw��ց�$>h�b ��ݘ�b���]?#�%����9��s 6�~ܸ_��>�|�ħ1��~� �]�s�p��`�M眣�� ��Y��+�] ��W��)��y�K�d�뺄��Z~������wHA�����n�N }E5,n���ruqA *A�\<���핞㎀'+�Ä��[��G��<��s}�h{�����٥��7[�</9N1/a����B��R��.v!�=��o�=X��|n���ʞ]Q�W�r�潯��}�>e�w��1E���\v�y|}u#9���g��r����Z筰B= Qt����5ͦ��F\ 3U��J:>9fϥ����+�$�`7�����w�#-٣�c�9QQ��jX��Y����9>g² ��5���M�En.g<�=b� g�g�/����1_L�)Ob�&�Ϯ0 {���F�N�x��ʬ m-9$,�}�8���ʶ����A�$���l"{�>����9xB��z���ĩ�X���ѫ:���eAO�P��x{Ƞ?G�b-�}���6V_�3�}�I@�m���D�s�BK���}Ael�p�Q�3K@ ��HN8%�1������\�/����h�{�*r<"���ȼ�V\���L!�n�h1���d��T|�p�P�m:S^�]�Z��c���1���Cb��A/�	��^�	��ٓ�{l�<R����{�pHB����0EGIK+�߷��L���Vi}�g���7�Z��YA�y��lM��g9ݵ���-y������3�	��;/���N��k�J6�ڔ�#����:��x��"��y�k3���LHU ըSy������o�.g��_���ȷ�~%K��y$�i�
��-�>���P���ՒW�� sZZ�����X�x���_�S��W�~�yS�]�X��|�?�B��o~\7\_`!v�k���)׬_���<<�C�І6�?�6 C�І6�?H{�艷y֗윀Ӈ~(�W+�}�6���C��*�࠾��E�Bg�����(u���bu=*{!�G���N˩CT�2�6�'��6��_�@6�d6��R��@Di-���@�J��A}q_�h�`�������AH�[T����od��sM�Ʒ�|-_}�)+a`��W��7��^�tN�Ʈ��o�%�.JP3/�����ӧ$ʢa5ݑ�DV�6$�֧Y���L_�}_ L�O��{u��@ �1xZ3���D�W�2�d��$X�X���8���cWU/�G��$�v�n�������ԩlHM;������Ņg��>��]�;���L������'8�kH�β� �@5ڎā��N&��@#@Q��n�5�?Sꋿ�x����uك��_G���3*�́��p������q\ݵ1��*F�=���I���A��ͽz �}�s[6���7 �,[�AN@� ��J�q"E��c���*�D%��� 7��<@�O`��,o�ޗހH��ƿכ%stp=��2�#B`��_ݓ��co��9�OoaC����d�� �
�,�к��م,1�QY�|�燖1����.'�S��|��8��i�td��*Ma0�Hא �J�zt���k��r#� z���߂���������AN wȼ 8�V�\3x���CO���J��bF2*K���MuZ�g_|)G'3�;�n����g46�皤�6NO��z+��O����+��"����l�����{�#����
�E��J����Ւ���r��ϒ�*-`嶍m�'�O�� ��}���������b�O$��6;����o�lƌ��T��on,����͚���3��zsӓ��]���d<�m�`��۝{��&���~�D*=V���iz�Y�5o�JϷ�S���̛��L��5�+���?*�'ٔ��F��9��qO���Ra@=,�c�o�FIBS�6g.GQ�y�����p���<~���ݚZVPՒ����m���?#���1~qy!g����mJ��Z "��VZQ��=b�s�6��]>'i���/�:�{���Uh(��LZ�SY�Y�C���WD�bOb�ö;GĽ�ī�,P��Uy�N
߷�	����ݚ�3I��q������tb�Y]�xX�:�$(���/9���,D���",����/�ԑ���DH�����\�r�[��`��=4a>M�,�:�1��J�ǝ�s�u���v�W:7��M�I�2�s� ��V~r_���kR*��rM"o�2"  :�>��b�@[/�;S&�u�\�ă��x�����Y��3O��N	EUFY�9��:(�A�B��b�L j<���$GU��+]���>�œD�[kͪ��]����+�K�pN��ـ���+�@?���eM{T���d��0��$�ٯnVk���rrv"o�������L�~�׎�A��<k5f=��k�\�ū�����2��]cs�-����i��s��K=�����_��Y,������o~����+�Ԓ��҃�iM�C�c;<W^��al��8�|q&?���G?��ܻw_N��H:#/$�3���o�'�@c����o�=������+/����\��o���I��L�B�,��]�F`4f 삠�x4����hw����l����F��)C�������;4 ޠ��U��/��p��}OY<��mhC��h2��mhC��E[���۫ky��s��3�C^��j/���[5�p�o���mm�L�k��$��ͫ����k�� ���$8�,��Ij{��k/BV�lh:>(C����p�A �����xMƑ�_�J�|�!�
�"���%��Q�f�{؛�<X��g H��EL�� ��n)�{� t��B}�gS�R�����o�Q�����0
EDZ��&T��a�H��`Wi��O��&�1��Ȏ��C&��+N�ЊGH��	Bö��C����?���x���� ȏk*����)"@B
�t��
��Mn1,�p� `��~�Di��R����y#
:�Wစ���SCY	ʊc�X5�諕A6�}��o�;�jP�a^�9>���(����Oy\�% T�0��Uͭ{Ї=
�nR7�cV�6U������o�+M�h,�����`���"�ڍ;T|2�#��̌	T'�J��q���&� �H�����b1�Q�k(#@Du�^Я������u�F�{��Q�l�.w3h|Vf��m��L���hŹ��qkJ��%��~�c.`����kQ�p�1��{k�U��iv��m/�o���J쳍��<�a�G$q,�~���$lC�K*(�i���b�6Ta8��F��7�1�I_9jc��,�,¼����۶qc� q���h��;���5+���~�X20y�j�4|�槼^$oo׼�q|'��������d�Q������_�y;rkݡ����<8�'�%�J��./�p�k����K�E� ��>v��^i;�C*���h7(j��䠷�sc���x�w���ߍf�`].=� �	>R���ϛU� a|Ɔ�WXI�k��ӕĮO�����BnX�c�r�j��k��l�W��9o.Z��y ���d]�E(B��'��Al'~��ޢ� k%Z���HI[{�h��~(� <��
U��$��y��%ߋ����L�.�Xwި����7#�� \@���E�����x��@}	U��(�:C�R��ؑ�{��ڝ�N��^5F�������	��z������ח~��n��P�#ݷ���W��2�|��};-T՗>��\UQ��K����X�e�X#}�m	AȚ�Ŏ߈p�\#�a�� f�`,�+�.�`s�'�����k�EfE�u�����²�����p�7�X"G+J~`6�S�G���=���ZS1̜j!˩[��tB��x<� �=*o�Bs�%��??
�}��A���ƾ�����U�C	��c+��4�xx;pGQ�;���+�����Һޛ�&��,�-RUj���P��=�U�o�=�=�����#�٧?�_����'���P����'r�=�B5��Z>b<`�9�#��C�2�
�v����u��w�x˽�d���c� ��_����G�ӗ���뷒��xױ�~�Rƣ�
�ONNe��3
MZ�������G�|*�?�J>��cw��a���m�k��	B6�]�-�b��#	q��>v{����"��'��_�=g�?���?�p�І6������ �І6�����7on���d�K\�h��8�<�ғ�u^��*d{�:<K���������rx��ߛ�W�o6i�ۖBͶQۄ0��9����t�O������`�@ٰ��	����P�I�Jp���2`nS�%�g���d��c�2B�g�sY����
6�e�~�%rs}�tS�,W4`W�ś7�x:?8�|��$Z�Eq��|�'�)P��0j�
�̓	� 
	X~0u��(Q��b�& `<�������H�Y!$?:��+TAM��/	����$�k�h�'� `���$"5� �U���q�~#^׳�ǥ�B5�gJ_�i��X#!�j~Cୢ���C�P��=	4��-�eB*H��j� <�o�%FT,�Yh"�A� �@���=xb��=dj�e#�o >�x.Q:�qv�.%܄}_3'���;�<��I�b�!�����yx�s.Z%wX�_�r��Ue��>�2*� l���c�j�XI<ľ.�i
�x�c�XŴ�3���Xyi�q֓O�6��_��53��C�ҋ���uO���W�	��L:�|^�.Ivľ?��|L�ᬍ�g�G���	�S �`�n�\qLaxE��EQ�τfDk% a]��­_1U^�s�1�2��%KE�>�UP`���y�V!���-5�״[���x���D}��E�+�O�"��O��oZf��3a{������b�uo��ԭœI��a��p�uź&��q��^˟�?+�*����9�wB�����: �8;���[�������N�^\��q}��nܚ�F^����n!E ��� ��4�x�8�X^�k*����V68~��㩪|�k�� ��� ���"�o1�ǡ�fd�o\���2��g�ٺ���u���Afb�.]_������)RB���N�j��T�T�����% �1�9po[lb�!�����\̹���ɦb,W��?���՞�؞]\��KTe�ִ���[@``����sG���!�ː
Ÿ_�U�4��`7����Cf��s�^]��}KB �AM�j	S_`��.����Jd��ԗf�e����j��p��]��[��޾���c�3���mU=d������K�^OZ�=	����F�b��@?��}��
tO���IT�E� uݓ-о��:�� ����8�s���b�����R.&��ԋi�<��j/�C������	$�x����h��6�!�-[Y0#%�"�e͞iI4dɘ{kM7��+C�@׽����Tu"���Xܑ� ������!P�ϐ*G���D3�H4a59s�B�g�F�_y�P]0�#.7��V4CJ�-��g��ߡ���grۋ;&����[�Ev������j+D��� �aO�}��͓�#����������w��9<�*��Ƞ��r���V�%���u$XbU�Z�a�d��A��BFr�B��
��m�����N������n~��n���}{�|��r-Wo/�39<<v{�=�@1�:�׷7r������_��r��,'8&�g���B�K��$�;��]f�B�2a�OQvT���1ɏA2��mhsm @�6��mh?Z[\_�Ƀ��;�����O>��{gwdp3��Bnoo���� �x2���\��ú����L��؛z?<�}�ձ�����xY$D��4�m�w�2O�yG��O|,;�#�j�E��P]�<�F�f��Z�l�r68
��pIo	��
�.�4f��mr`uqr��W Pa�pI��h��羖���<<�#?E}�#�"d`6��8���PL@�7�P+����cco# ��m5�Z�̿:�݃٬'6�M`�y�*O�o��"��|-�1;�Ҵ�X\�Sp�*���0Q �Yb��Ծ�@!C��A��Jn���Փ
�5�W|��i�@��9�h�d�焁'x<���*_Z}���3 ���(��{H�3=�9dTZ�Lb�^g�MCX�7/q��P�m�DD�ӪDK��hQ�xb����^���Y)��[�%@��x��j��7�g����A�1A<���|謶�F®�EF�﷬J�`�U$49�1������1����g��B�[���?��*��P����oy�*�mS��@?+{�N3U�f�(���Ԥ�{]^]�z��G����`�#*�y;���є�]
*Ҿ���Ȟ��~!9�;�~u�cj,S^{U�$>�D	5(k��,@7��F�S���yǱ�+�@nO��`�K�Ea�{M�5�ENǵ�2��%o	�jT8��:�B�T�,�,n�rw�+����kG�]+1��w�bU(������3����k��˓�#999��;�~�xpz"ǳ����~x_^�?�/^���	��j�s l�v��7��j�2]7��*ƨ@��^�|&x���T��1ۥ� ,-� �"�h�?��H:�}�Y`�dn�u52Rֲ�^��d�`t�b�ִ[�H�dD�	�e� l�~�G��w�;�uT�eV�D�'���R��f�`�U�>͌��"�nh-6u$�������0�B"�)Z! ���VU� ��8����`D�YW�Ϧ��gY!x-��T��	�c�x�6������ʋ�Sba���8h�]���߳y`�A���$���Y�Ҿ��������u	�2��{E�~���/�#wY�&!G	�-�Us:bU_���3�^��8&�l��2FTYa*\Kd�ڸ��{����"���n��2IXU/=��{7�0waEi�%�v\�8#�S��
K��R�`:ƌfx���f���Y�@;:��T6\�44}b\Z(��ܹ�	%;��o�ͬՒ
�nv�'خ���S;=��g�v� ��hŻ��j]�>�A��=�E�,�{2�39�.��n�_0�q���\�6�����H������R�]�rܟ:�@� } +*(�>z�]�짟��`��ߓ��jBo��3�������eo#��^�  f~��d]����P,~�R{£�c9�._|�3���odys�.y��� cpO�q�Xy_���m�cL�=�U���^�g��6�|��v%��7�������t2�},?�-�Ȁ� ��/����|�o�A�6���o��І6���Gi����'Ӊ��ߗ?�P>~"�h���õ<��T��3PY̠�M.k��o�B�C�Q�g���~�X�Wr}�VZTJv�-2,1���= ����<z�.����	PRf�X��ABۏ��$�X	�%���(��8X�xnx��PU^&�����p�]�o6�qY�� AP�${����6'�Gh4Z1W�a�!��� a={�g�Pax,4j���><h�#<���,�VJfI(
 �����0��+?�]�KQ��g|��
@T˔h��bG�;M�~� ����@,'M��� }{������j���SifC��l�X�W��EjVEM_eN�Ju;0��s��eV"��N���h5�M 0H}s�dg��ӉH)Hk+yq��v}N�(�2��G͢�<W$�� %��W'3����9~N�8�Fmڮ�.���.�A ap������1��Td[D)`���k����x���$ϴ
��쏖�ao�E�9{/~���v3�A��u���ƾ̞F��d�����@Q�y��I�6�� �c���� ��f�"��C��cE e��-{��5����	�k�p��H�)q"t��ՒZve=��ɏAG�oѺc0b��e�rڎkW��ǀ{.g��D2�d�`�J�-����ɘJ�mU�$�[_�����J����a S�� �r k-�Jh�ˑIJRb�����sa֋��ܿ����H����H�Rb��9�w$���\]]ɋ����F���d�>oy�`~,T�"��p.�}��C�<l� �B����ź�ZL�3S���F3��}���w��}Pb���n��k�4�5�!�*򲖭��k����{��Ls�j�1�;C�ș�h�s�Z�r��(��J�F�}$����sGU]�57'��Y@Ԍ��8.���fTT����K�8Q��z�����T����^ͥ�\j���k9�#�ܰ�CUi�P �16��s`�^�%�~�)�Z?��a�cm���?2�F���uؾ�vD;4ڂ�ͦ�VRU���U�.�
 ��zݶ��d�|�!�1��u�����=��%�o t�'�Sk��A���]Y�=�"���;�m��;ٵ4�/�m� ���ah�J��"d��#�N��R$T�Kc{uI���>P��$�}He>l�|.�(��j�v"֚�;�qo#��P�E�CzK&X�*
$�,,]?�����Y`��Zi�{�=��E-�:҅�u�^��d8��x�*gD�6�^z�6֡����{������/�omْ����e����a�~����������j�֗zo_'����6�O�<�'O�ȓ���5],�8߰�b��}�/��RWo#�,T��خ{k-�Pv��/�ƽ�'>yG�|�zo{���f�L�{�}�����r�������fqKi���}�Q3�ڃ�39;9��ͭ\]\ȭ[�n�>��槕��[��z{�F^>���[�7������Y�r߽^�Z��ۓ�x���R�X�T�a��mhC����@�mhC��~Ԇ���|�dp n�2l[DR�47 �b'�n
V�.�[�BBtt��a�
 ?� ='�G���sj)���M!,K|�'@�������x:�҄ -��Nj x(ǧ �s�깞@� <���v�d��8^��>�ڤ��5�xΑe;4,;6F�{�ف�Ld;��^���a#�*�Czٷ�� |0���@Sc�+,3�P��Lo�*�o��<�6"I@�l� �\�Q��">��@g��
�VGpת�c_}m6/x�X�V	+�Q9�pY�g �@L���5PM���vI%U!�`�� lV������|�Q�J��@�A�.o��D�p����JЮ���.��  ԒD-׌�b��'}*_]��mI�A�p�'X@��jec4� WT=<(o��V� �Z}��_���Y<�l�!�T �
	��q����c�J|)�0ȰpIt| Xm@���}+�CUX���hEp�Vp�� ���2���Z�͸���g��#���^�y$���M��<��������7QH�U�:7B�QY����޵>��ʣ�0�?
S����
�@:
��<)�E�(��sQ���[�R���\�m�j�u��K�$+�ˌ���:�i%�ЎL�Γ��&�Җf�\�-�\����Jb`ğ��r��A����si�>����J��dFU2�������Vm�a�n.�
�s��me�/e���uz�
��#؆ש"!�����r�xN`�v�"����+y����z��YPV��hF!�U��ݳ #��,��'���]���검� �jw.�m)��F��Tׯ 8����<6��e�H٪�-��A�`l����v�e����WT��&�uψ㙡� ���ٚʹOb�`�F��Tj�*�%~l�\W�\�
�rL�$����%��%�?��~(;�[�d�d����a�U�#�5P�f��ƍq(u`�5�f%��R�����eR��=�z����8o�Y�����B���A�:��T�
�����\�LMB�����K�u	{2�
��넾Ɯ��+UI��?ο�:W�M��"O���-���[n;���1;֞�"u��	����=���&�-������\�KQQ�V�ɔ'na�j֑�qE�iZ+�����4E����`?��kԴ�ohvu�����
�E�m��i'���ېwC�P�B��/*^��P��e��@���+�͹c͜ ��*ň�^c����ޣ���x�K��Tya=m��6yŬ��tF;@+��{���`�+Ͷ���)����O�y$�������$5��AH���`<!����G���D�lV���S-�5�W���|��5~2;`({:�阔�r��b���O� y�������MK���D�!�GG2��5�������x��n��Խ��?��|�������q����,6kw�kw=����	P�=|�T�<�'�ߓQ:����~�w�"����mhC�_��mhCڏ�޾x�P�C��Y���^��}�������}�������=~��������ߗ'O��������@!��`����[������퍂��&t��Ӈ��a�ѣǬ��A /ʹj��VB�BE	X@�SV�L�_�k@�_~�<���Ko%P���㱷�hY5[�?��u:˽�SVQ����<p��ϸ�x�W4 P�!,�m�j���`���b� .��5�(iU�H��W�FTx�ro����쬠4�f�&�|��Gx��@����-�gz����B��#���1������V�U��(l�F���˯�3�"�4"	�<H�U� �QIB�D��.��V;�Yxi�l�}�)� (6&���u�z����& �޻�O�j�`��48����`U=x�Fa;{�4d4^��~$�]����/T���|	6'����^Y��d��4�Y=Q��H���%����I`?Q�HP;�4m����GC�a�D� ���0�*��1+�U�쐊��Y�(H��l0��[�Oɋ-�H�y���ܺs�M{ ����x�X�g�3�|�рm���� �i���Fz�K�Q-����f�h�|��vU��Vή6+g#��#�k���ȓq5� ���T@�
i9C���2�V'�yg�.�P�#2$Z����9��"@/�V�l��	�<�X�ϳ���VvϧsZj.+׿��%q1:w�u�� Ц�߰F��Q@Z	<Z��?ag2e�6��B�y�T�� $�v��ˋ��N̞p�&�09b�����̧�Z�<�?xW.�\�k��]�yK�x���6�:,���@:μr��ik)1��u �A �䌸ޗn��&�r�d������ j2�	��vJ$;�����5]��4lQ��6K^�0�H
��TI�|�Nf�*A�2�
%�x�yD��j}�P����d:���Rm�Ч��@������Y�-� K"��H� NBa,�n�S��M�'��L3���	������BN�OxM��/�^F�
ܟ�,Ğ�?����2���M)Qa{��t��uIeD���-�p��|�uP�_���֩j�V`V��dJ&��a�a��kqFȵ��]n�Cɧj�F��X]�0��:Pడ��<1��Dn,<u���f�����
�=SǠϔ���3˰��r��zA�����3Ȃi��Rj�ʇ�0�HȊ�)e!�*�{Pd��U��] ����Hc�e$ӍĎ��d�{�Qjk��$n���Ũh
�{%hƈD�m�mM��98�(T�J��\�,3���l<���+��X2��N�z5������ʪg��Ծ�JAB	{2��^��@+z��Wo��摔Eӓ5X�AĔ��5�?�+rs�[ǧG��'��|@˪˷!+,gJ�u]n98��h��W>D� �#z�6�777�XXP}��#��`��l~(�#�'�s��.���[��O�C{ۋׯe�^��2Hn����Cyx��G#�"�r�?r�p�$��{�~.eϞ=�?��O�ɗ����#�ԫw�^,����=���(0 ���㰙�����І6���� �І6���(�vyˇλŭ������o�a���~+g�������B�NOI�\^^���V	ϧ3y�~@x���	C,'i��������_��w���K�@�e�?,�� |�C^䞘^B9gR�>ԡ��DE�ੂ����UI�)x<>=�Tm�����lx��0�"T������:$A�P���.��Q�+�Ղ���a�t0��zy'�f��Z������L���ɧ�~&�����۷�R�֔-dC	��}%�6�KPE��T.�U/p�=V�'�U����@M��Z0�A <��x�9������~Ջ	<�Z�z�[3d�9(��^��4'�UҲ�B.����vZ��`YP܀8����l�>�(\N���va�h��W{�T+g���K������_��*jV/��Uϰ�aPt���#�^	����ð:��~	�$�j�b5�Z�u$JhU+!��a>�c/H��v�h�ߎ��M�U�x�&�^kXb���oh EҶ"�G�� Y7jD��� �Ӭ��i�*3;w}�> ��ȝ�f� V�5J��E��3AH1�$X�vc��.@��&_��"���d�w����"]�k�J��nE��7�%JT�w�?3f0`L���!x�<Z5�����&Z�L�t���n���Nu��[p�St��Tl��o}F�l04�DU=f"�}��~*�"���E+��$l�¬U��/ �������5��5 G���7��+؛�ix{{'�[ߦ Ǡ<��ڶ��%\��٘W��煮�  >�V�M'}Q�_�]�m"�נm�!!�ܼ�jٶ+Y�k��}&W�����Ǭ8N�g ��Z3yx&��������Vn���ի7���������}$�;S�y��b��Qۃ�b60��.�ͪp_[ik�'c�2�YZ߭��I8�K�e�^P��D	Aj��u�
3 ׊Z=�"�,��Frx0�|ٶ�,IlN��IPO���=�b�*9�j�έ3
e�������Ӎ�� @V������52&țx���n ;ć��M[o�[��Q���W(hqOG���}�_���r�c)����y?V��>�(%Y�5�ڍ��ÿ�B�M1��Vaou�RɲI
��I�e�?��3���{�f�e�D���@I�P��<1�π�Wj���zG�Y�\Z7w�QFRvm)H�bù5�U��+��	W'V��"7F|��*lw&Q��OO���ԭ��E�\O�S�U�H.(8`�$$��=j��I�z2!V".u�J�M��dX��]���#%|E�*+X���J���ܔ@�W���:�1w�$�f@�^�y�:�P�2��}Ԛ��ܱ8V[�$M|�T�G V�׃���i����BA�n�}��]�wHn"�u3������5����!�.���땜+5�>l������MĎ{!w ӹ<y���o��� �EY��%~�5<�=��*��hH�bߜ�5v��U\'Zى��xO�ɿ�R[>�ǐ�I^(RB�^7s�v�@f���]_��`����n��(���ù;�)��lN�B��8��F6�7�T�@���<7&G�Zs��+kP��Ƚ�M���%��%~K�6��mh�m @�6��mh���/��x �=X�u���J޼z��
�H |\����졄��7��)��x&�N�ߌ>�-,�:�v��������y��wr���lV�� 4:��K�N�gn�޽����{��*b�i�5u�_X�jzJ�2��X �G��{�Z�O�w��Vۧ��x�Z�z�Pk �xo��[ki�9==�����	+�N@�3,��q�p�˔�+9{x">��:��*��?X���t�jM+*(�o��={Fc�J� ����fo4j�B�`^�k������������E M+�������a-}��_�Tm`I�ѶjLҩ�U� "P�*?f�Nxmj)	�MG�Y
0�Q|:�.���dL5@׿mU�0{%He����k�jT�
��鄪
 yh��0�a띲��P)��r�р[�0�u�jb6=���vש�����b�; ᅻ�O�J��XݑhA�>�U��Z�0=I�{����`�C% F����R�Xw� @i�1�Jo���� ,p� w |E�&��A�u�s=Z�cV�G�,����R�J� Є��J�m��9����� pۯ��K�}���@FQ5%30�@pp�u>���AH�I��LF�BXl%���[Vd���F��
���z��P���:!�:d��Z��Y�=h���ji�,�y�&Th�T8A��ٗ�:�@�h�K(�'@g 0@�QJb
KH���8���nEPj2	I�Q�P(A%��B�	�����A<=a`-� �Q��0�a6��tZ���$w�x��?��s�r�YHbƭ�'�G���o���+�;�H�J�Z�f�Lg�L���9ힶ$!K)��+���9r�A̹z��Z�t��9H	;�OS��#�ӻ�y��T>}���}*��O���W���������s}w'�u���Aۘ���b��Ľ'fa��>�=VAp~ ���9P v�R��& ��|ڸ�`3@N�~8�&t׸v}�>�n���gk_���{W7�\`wx8J���~�@�:'y5u������	���M�sN`��\]��k,,q"�3o�X?::�*ܘ�J �UE�����OݘM4D9*Q*7��, 
XW�T�$����Id����� ք�Ɇ�����37�Frss��k�+cGn���.~`���n�mܾ����& ڭI���uт�CƓ�XCԞ�b_b-��%��Wj�g$���[P���NTr\�Pa�>5������ld�ΖY�@{�	��j�4�pp��K2/�D.
�C�Y�;_�@��6�n��)�����o�z�+.A$/P A۩$% r�7J�T���"�{��S��=�Bm���>��ٹ�;��Ֆ�+^3�~�5 4�����?�8��[khc���^��k�" ��uG�EF�\�0S���-�Ztc�s�+ �I.!�{��?���Hz;F�g��|�֍�GC��y$+�֣/5<|*�[��u���@չU�g�P����5l�@��y��7׬ܽ�)q?TQ=Tj!�4���n6\�a���}���k讵�}���{���qTG���{�x
b1�߽�S�䃟0�kE�o���l��q�{-�f�����z�!��ϩ�ƫ'�܍'�Fn̏��Օ/j�t��ͫ���߶��Z�oES���N�Jm3Z����ߑ���C���7nN\���}m���ǽ�tv@��s�m<9��3v������9ב�7����]�N��F�ޯ��s�2�{��]�'������y&C�І6���6 C�І6��YU5��ݝd !�Ch��rs{%K�` �������[V�?~�|��O�W���<y��@ o��V�N..��w_%���/�������{?�@-��3 {)+��r�G�5T�-*(;4�~H�l�;A�6��X��d�i����u�x�w|ޮ�2C"V+�8�#������*aZ%ܿ�z����<x/܃7*�X���r��#y�J�F�rC��Y���?�_�	��A�(5� `KĽ7|���jv�(s0���>���/��G�Ɔu�{(H�	b��V�Z@^gY� �1^�I�Wq�#%|��=��x�*�5C-�v��T,4��
��<uۨ EU%�E㝕�VO4���}����"�[�	�o�b@���Y��}TH"a� ���/hd�k�;����3���zwf�*�����8Q�HHL�»��xH���6�����;��_��������jiC�/R0��%�}�qCe	��S���13 �.�]�>4�&	��	��f��u:���c�>�]�A� M4+Fϻb����R�76p��
.��Y�	���V�c��Ҏ|i�������F3�G��c
�Z������
�~�$(Z��YV�VPj�I~�zy$ !����G�6� �H�ta}��U�>;��$��|IRa��T��R�d����*G'r0;t�(U�.�e��i��ެ�/2���<$���d�5�ƭ�����a¿��cnK����[w�8fw]��*���� ��;�����#9>:d��{�>fp��ׯ�ٟ_�śky��*���!����,��0e�>��Ù�%A���M@[V~p���|�0�ߒ�-��5�r��,�c��,A��cu7*�[�Bڒ����F\ms��T1�~��u.$ lc���ʅy�Z1�E�l6�X��\�k�k�H2�+lj��iF�PɃk�a޹����BK��l9�
��܍U�/�Ky���]�~��䐀2�?�j�l:���}�4ϳ|NM��([CAFٺjvV��ޤ�3�������*�^d
S�XH㳔�>��H�,"��4[��sF0�m]!Ś���$ILZ���&�
ET��	�{����X�u��X�jQϱ�5�?լ����Y���n}�I�ש�#���*A٨�3�(�X{*]ǓQ��#;p�(v�u��b���g��>�<&9��"�׺�h��a�;G� �"���<�{-�w��r��J*���8��>�Q�U�5L�TK�߰�C������{�����E# �3*RF��Ս���p�{1G-�iOJ�=�z���T�� ��f��L���Q�R+��b����O���ܽZHb��0V%�����m��_� �I��s��O+ͳkt�:�\>w���h�|iԎ
E-�:�9�-�9��Dk�ղ�A<8�G�ɫ7��[��B�3q��%��kQXcy:��Ͷ�ro6=�?���UP�-eusǼ����1�p�u�,��~������p��u�v'j��_�����i�����mhC�_��mhCڏ�|GC^{0�`�>x2�7�n�f��ݓ/~�3�O���������h�v�ϟ�Y~��_�?���r��� ���P=H�$����79�;OO�Y9��������ѭA�fq�՛�I��B���
"w�Ń"�,�'�g� ݄����z��$A�>��t?�ăz�P��A.V�gr_�����=�-|6@��,�C�۫+����0i ��>�C)���G��<��F���@K<���.$��*̂XQ�*Ѧ3�!�-� ��H&(#8�Z�3�!F�M����\��wJpW_gU����j����x��=�'
s�H�ڶ� ���Y���8.?,	�����f1���W�F$���S�{��]���	�����eq4{cH���[����z��c/,���Jt��Q�CVԢJ`��0UP�" �>b�~��E<�bA��I�6h~���]ჺA�`i*���aZ�Y�?Ճ]ϱ�!�"����I��g`-A�jUu� ��PNZ�����������$���'<�f�����tj|���� ͻ9 �o��M��~*�}�m@����y{���>�=R= �`��9���["X7Ú��G84�,#�IWE?� ���|X=��c������A���18mؽL��#���=99���� �J?�P�K�*�I��.ܘ�uը��D��9��^����Z��X��U/dz H<rǔӊ���rK��� ���\��?��ʃ�sy��|��G���ҭ�7�/���|�V^�z�������ja�UlVR�����Lß�N-cZ[�5��A�c#YW�$p��%E�F��ժ� �F�}�����
ύ���HNONeSl���U��\*X���u�X3q����,�_�[%q�p��:���˅�v}�� �f��^V � ���tƹ����V� �H$*dhI'KUy1� � ��t�P���vqqMKH�G�I	�JyB��5�{�.�&3O��:��2�}ة�?Ӟ����#G,H��'u߭�F��l�8�O�&��vF�Yl�}�Y��Ϊ���5Jf4�3�q�(,{����3��OC���f�o��"�(�}dd�����t�K�XH�N��
(R�m���6W%���ZBak��Ϧ�߸���F���>����6�e���W/��lj��Xkj����ZX�U��CL�N����+_H����;[R��8��c߯�����j��P3�^3�Ma����#�1�d�K�7��)�e�&��s�[��Q��u޸u�D:�	�l�]q��/b�*�rMݚ?�����ޣ}�k���#*א/��	�T���r{w�cɋJ�w���`���� aa�|�rޡ�V��<���c�7/^�pk�3&PV`�@u��F�xCY��2w�1?<����@^_���o/z�-s^<��YoI�q�qk�z���c��e�gg�r�����BVw+Um7z?�B\`��j�(��>�u��
�� �޾y#C�І6���6 C�І6����R��m}'�d���)�Y�>|�X>��Cy�=<����{�`r�]m ��y-����������UƑf@�&)XAB �'�) ?��o�ƭ�>Q���VK#���=Ќ������ � �ke�۰xB���)-�@h��!�W�PGOu�tv����r��
]C����M8��`*�Ʉ��QY���{(Ge"@Ue��}Ps�=����%l�' z�ۜ �ވ�Er�M�75�{Q�o`͞;ZC��+)X}�)�����Q5ZMn�	l��D�!Zz�{�#ړ��,B��`.��.,}(��l��o�#�xP���V;�c� ��6�wͬ���6�N�4������g��"L�U���~�n�Fў��g�1���l�r����9=ƨ������>��>�f}i$Ư�!Z�e����e\,�@VB&jŴ�� M�	=v�Ÿb��=f�-�	�ꣾo1�^��~���^+��ߝ/���ጾ��[�P`պ��b��8vVҗ9��
�4�0x��1�>�$��x��	�7Մ�a%'"=8��a{�E�"�yj�n$��6>L[	-�Ќ���r>�FUB��Q0��O��0�D���E(9֧0M�Yf	�� b��Ko;��I�.�����ӧT�%�֜�v׵�y�8�(:$�u�js�ǰ��w�7@����48�w*#7�`�t��[�W�D@�< ��Ci1>@�#��]e!˻��}����P5� y��;r������O�y������|+Ϟ�Y�������昇��[Ź��,U��
#|9�|�DmQ��2N��8�M�Ǎ���GR��z��(	ت�����t�{�j�lj�`����'duh�Ԅ��3ˀkb�8T�O#s�����aͥ |C������^����|�$�Ӫ��� @P������|@��qT�[��QU�[2L�#w�W܋B*�Ƭ���ڱ��'�s��<=���n��g�x����B3R���YUٺm�Y�a϶L#>��02�	|OI��_��5�3=��k�ؓ ��p��� ��tT
�H�5=�S｟��kl]Q��*�N��`�nJ9;�c��;H7�%d�yo�6H�@�5�^�����{�*w{G��#H�� �/-��2;�,x�u8рs~n�G.�hlb�)*X%R@b�@�D��j���u̢��Ǆ�?؂a��S�"�'Ђ���M?�Pc�׮�Ru�3[J����y��D`�τ��f��?���}I�UD�E�D��y7^}�� Yߒ q?w��9J�[�q͸�&^qXs�=Q[a 	���Pp.�)�.���Ľ�1���XߠT�����[X�}��'���#�Ob��g=�L^�|�{[c8!��XCǣ���G�Gr|�L�NN��� z��~O�n]�ݚL��t*+��A���{R���FaL[��\w��k�q���<�{���=c`=LGn��/��Gn����駟�І6���o��І6���Gi� 1� �F�W���NOO���ߗ������.����N	v'���o��o��7y����y�B���W�3tO}q�a6���:��x�'�m�j�z�����% Yl��.{ V�, y�uJp@�vv&�ٴ�����'�C$I���T� @�J���+��K� �t�+�Y)=Ҋ��VÑX4�
�� �Dht��'-	r��f�>J����*Z@8l����hiտ�чo�P��-.�5 Ho��m'��p �� ߚnP����Yz�G�T/�ڐ���p@�-�<�^��XT�|��a��W�F��d��K�$ zQ�	b@|H��P�� P��Z���C|����Ij�DN�/(yXY$}�/��+�9����+ W�-��	#P���{����b���f����cL#���%�|����9�-h�p'� m�cf���VA"!Kǒ&���K�ƎJ���
�u|�MEm�h%z��I��v�v����6/��
n�d�U���2�KɆ���U��$��?c=���;-�|5.�( �b�OFTټ�����'Q&���E#@
��Ҁ{(`�
��ú�"x܄%
(�Q�rt⣠��Z�Z�����څ�����ߨK%�"(��)�p�F��N�}�u(U�������͹��8�d,�9��<�9 B�>����۾
>�J9�}�G��F #p����KB�#Ώ:hd2�r,bl �b�N���Re�Y9����QY�.E�����\���v%/^��ÃcZc=~穜?z(�q&?y�<yt.77��o�ٳg�����u���L��:
� ��X[�q#נB��v�~�I|��j�q�
.�~[m�7 �f9	'��t�`}���7it�����vQ[�㚂�-G�cZW���<!8��A�B�k
�Q�f 5�n�\h�@O�v���.x�yK0�R2w����w璦9��ҫ�F-� \�}��j)��%�W/(yQy��g����`��*��ʽu�X��ύQLs�iB[ ��1^B� ��Pq��Q)�V� o8~�w�-��WF��-�>�mk�>�l6W�f�+�l�2[LV�{�^��0�Ś�Q�Ŗ����Fb)���󺣺j�Ɠ/��c}o�oc���,��f�X���^҄;e����B�n}�w��00�m������'�/�Be3�͘;�WA��&�q1��~2GC������5C<�l1,X#Ȃ�����j����N6�g#�YJ�p��
QU�D!�A��m�H+�J�S�r))T���������{"����e�2T=�������'�RU�e���0M�
��iI;X��L�Ӑ�Nu<��P�d�su��8Ӏw\\\����/��|2���u��ݗw��	�y:ކ���1H��[��Mwr|_�١tnm<t�g�s�v�e_��:-AQ�0M�n-H,3�íKP2s� 1ֆJD�k���@�T�r����5zXOp�"����Э�K�P�rY	��TA��%�xB&G''�$��//ehC�І���dhC�І���ʃ�h D���ز��s<�����������?s/��</��X��������'Y.�Y��]�je�{p�dLowd'lWYoK��h����VG ��@���Z)IVX������ �����Q�)h�*:TjWu�{��!q�\,@�,� !d��A�'��Be�f�>� QaUz��(Hno$ґz4�^�U�Pw0$>^6?$1b�<�$*� g�"�*sD �m'݄{�^ۊ�F� ���7I�t�k Տ�N9
�NI�f��hV�i�
N��@:V=���4��Z���ϲ�q��F�D{�G�;BZ�Q�^�qH��*z�PP ��|�9a0y�Y
�ZO �u@ ���$��(kI�ع�1���66�A2 �'V�6֍t���i �Pq�����aˠfZ�y��@~(����~�L�so����J������Nu��y��D�`�y�� �J�<�b���UMÞy�k�e�|ۿ���� @)�:Ж�N��� ��s��S~w]hjH��1>D|�2��nִ�H�	_�z[k�מ0亂�V#[^W�M�+���(	��g�d��ד@�c-�8��QU ``���t"{ݮ��+Q��������c<�����$)2 ��K�S%=�Zmi��2C6$˵���j���MQh��O���L�+��������f]�"�G�s��H��j��\ke0�_���E}'u��1���ٔǾv�qws#ח7�ݷ��W_}%�����ޕ��9>>����}��<}|.��rus+_}�s��.Ɯ�ۋ�����^s�>�d0��tV��:��âI�[*.z�X2N7ٖ��B���V��n�j#wM��Uv����P>$
ꂰ ��@o��Y�� %
�>���VK:&k.�x=�ƅ;O�q�s�����@+Щ�q��ք�FcΟ�:oQ�m +�D���Io�W�,�>��|+�O�D�5G��݂{��+n@��~M�=J� ��� �Z(�n�)~o?�P��Cv��4Mz�����v>��2������#l�P=���`�ٓ�%W��3�gv�k���,�D��я�f�γ�Wjݯ�f���t/h��o�3�l5^AD���[�A���F&ǜ{������ͷ4���CX����`��{�T��.�܇�&?I��l;�bX�pu0��5�a���
� LmF�kN��v�%�'�����]3@^��p$��O��c��0�c-��:��5��!��Y�zkP�ӵ�%g��ci�I}%��#��ܺ΢�>��fҪ՘^���n.��s �[_��q��c�灺f5Б��\�C����ڭ�E��RՁ!�`��g�qOр1Ů�y1���&�Pk�
ϟ�f��KXgv�� w��"\�MŊ������~ׄ�Oŵ��>�b�ؽ���o����2?<��>���&E��7skg�{<IV�V����*y�� ±�������g�?�Q~����j!����,_~�%�ޡmhC�_��mhCڏ�X�[W^����{rrv&��/�+��g?�¢���V�a�Ͽ���?�������Jf�a�|��p�~��� �O+���T�{(���b I��� 8�*ux9k����q��TI$!U�V� ���`%ح�]/WZ��䈠�Z�0k��6���]��2;P��e�>�v	�c���G�/�Fc����?�& �z�'>`�g92Vz��:hxz.U�3� �@���d��O��"�ؼ��{��=��?�n��Z?"��*_�Gh6À���HF��G�C�Y���TJ�)Z�1-@�b�� �q�$J���.}V��ծ"�7���].J��L����~u��s\SUh���*}t��x���ư���aaV*��՘�+@X񞺀�}��6+�7�_�N6�]��΢J�'T��8����� b���k�� ��ƹ1ļ���-��I{5����r�*������;��X�V�)��k���弪˶�9��v
F�x겿� �F8�\�jh/� Auu�>&���&o8NR�
�Ŧ
���&���
'%(�P�a}b�����|����l9w����X��#(=��w�k����=��| ���w���~� ��c��i��s+,A�*����ĭ���8=<��Λ���p�&�s:����ި� B���b��R�P5C��F=(,�Re1c58@���CQwxx�1�_S�w �6��@����̛��n�6{�u������\]]���@=d:17��H����d"�b���o���B^�vsj-�^�$a�0�΀�F 2#�k�# ��/�;��C�8�9�����~��uAB���!-"�j�Av�\�����̔	4C�v�7�^�صjJ�.�~`��+8}Q'K�7�MY���(�t���_B�c��k�8��'���~3� {� �)d�In�}�s�W�������v�Q���� ~��X�(
�����?G;O�y䚄u(�~a�����l^�a���ƘQU\�3%v�5#M��#�?���<���4˫�6r/憎���ȾJ���p2�ۥ�Wn�5$V|:�S��� Q��;W%�2�nYtk8���ⱄ��a.oA~�2��2��
x_�B����9��_������^��F���~�p�5K�`wm�O;O�yUd�hD�Z6�bo�J��sȆPr�g���$��2	�0�N�~uOn��=́�B� �bʿx��Y0��7��� c$��(��k��B��c��21/:�{��8_�.�]V�/ܧ�6��ƜdP�bo�}���tT�P kg�	H���<yJ�O>���X-I(*�*<*�����ƭ�~J�����\���f���a����p{�ԭ��Gsy�½7�1�
��a7Xy�Ʉ�D��ݿpl�~�/�p������T���Uyo�B� 二��Ʈ��՟_�?����k7>�2?��І6���o��І6���Gip;��Cςթi"������G�������#.d���y�Ju�h�z��uYz$��\A��+�CT����2A܃*�[Zf�|�l� �VCjU�&��s<4�U�PE��5֊̺R��{=��$x8Z
��F���6R㊭���l�I^��е��[�vq'G'�}��fI4�S&  �=Ȃ� ���4NU� ���j>�W��)��jTE�	��:x��q�	{/T�"K��;#���'���6�h��f#hp��MV� �|��~�[�������<@7��
�,S�H��[HE Q�-�S	4�{�Hij%?���c����5 �e������������\h�}�z�������X���H��P1�|�i���@4�0&$�ϰ
e#<Ь�خ%�tl*�##�N������< �ؑ�Hz����CT���V�-�pn��2��PO���G�^��?'�0���{�1���!/dGr0�VJ'�u��%����9�}��|Ƹ�k����~F��s&�9������Z�RY�q�[����QBժ�8wm�m�o[����݆w �ņ�2u�?a	�O��^5��^�}�Y�;���_��!+����U� 3Ԇ( ���
����#9:>�`�\�<�𡅚��PU}�x��k�w �Q�8�H �*�a�{"7�֫-^��F�r_P����V�٭��t�3���z{�Sα��`S�O����B�s�t�v3c�@�e����Ņl�#y���-8'��ى�?Fr|vO><��O�'���ݳ��o_}#W���"Z��s����
	��I\T;״*,H.G�[�o�1��-����f���s	kt���m��@���8p�u
�s��)�~I4"�1���tO0c-B�5�O�Q�uNQ4A�c��$�øZY�
�ϧ���.�1o �Ls��y�z�}����|,�F-!1��-�E%��Q�$��6��
*�6oi#g���Vh|�+(�Uz;��P��T��]����Sb�n��i;O��NBú��2I�sH��j�,�~`�gk�)�>����In�������!��5e�,��2�,�i?g��m���ح9�u6�U/�שR�M�
9F塚���sI��Y-9�ݲ���1��E�VI7@�J�%�`��u"ȷ���ؔ����hVN��r�C╧ /CU��ǣ�V%_EFN���ԼW�ώ�2��J�O0�����VL#��J	��H�N�zp�0�4�v� \q}@��b�s�p#C5��3w�� G����� iŌ��1�H�YTW���z�o���:qkr=�>`L�o<�x}mo֡�L��w���ݍ\\]R���)��{��(��4��dR��)�����߃�&�x���fn\@�S�������� ���y��>� pޭ��GP��s���a��k���Xj7N��������ȗ�������T����!��І6���m�� �І6����7�E�����{'����_�O�3y��	� �4����4�{6�<��?��>�P�����d�)�����'�YM��ߺ�N�o��Ϥe�&��ՏK����_X��(mM�^s �G�v��r6c�4��׹{�ۺ�[�7&�����F�9m�����_�?����#��� fGcn� �ooe:C�y��PZ�hΫ��e��t�F������9�yA�5)�œ>��-�d *���v�pZUV��Y+��Yȏ�Q��H���a�lъ?U��Z���!�"����
8���RU�*�' ���.��A6��f �B�o_Ӳ�z�%
��;�hgW�z���g��;+p�σ�z�TĻ/��{�BL�|+�?w<��j*Zr������Ѭ��ˢ��2p����%�Rh�)��Jk|���y������V�?����R	�������z���K+Nw��]Oh��3���B�Quo@K�+V���:�8�h����l S�쪔�0��S��`�*#��&'��y�������V6e혳����0W{�Z��$�Q_��!�悈��P�)|�g�qM�k�y@���t�Ji�#AifP�Ŋ} y+(@XX�6�[٨���U�y��*
����Kc*�0�`)d�d �0'�٘����J)U�����~��mR�s׽`21�;u��o�n�����\I
*�ǖK�PB@�DC��<��1��i5�����z
���#�6�oX��Jb�: �6��`�%
��g�j�r�X�z/g�N�� �WW���!T���ƍ�;�� �0.�+�v������ ��D8���H��q���˻������x�\���+�1�b:f�x�E.۪a_�"��0YU_Ri��$���6�v���)�殺�5Q��6�Y��%�d<!���ล���	���vfww7��5�J#�u��zj��r���� ��hnS��&䵾��$�R�� ��:�a�*��c� �⎠e������`~?~�� ���;_7�E��]U�}	D_�V	|1ä�S�ykB�[X���Rת������J0�,�d-5r۔�w�z����S��Q������Wp������� >;��>������U}�6��g��8Ao{�����ֆ�5�����d� 9B鍰������$X~S2J���S����?�$�b�;�>�f���5�[�N֭�˝�Z	���I�Tf�����8��P�%�B�m A�#GÍG��?��Y��ڝ#��rd��k�T�����6ފ"��$ͽ� s��9K�A?���E���n�Nz��B0��,)�ޔL/Y�S�9Y�µ�U�g��T�oI%.>c��i�T���m��ʍ1���'��G��Z��utc����T?�%$�眗 $p�	b��ՒcY+㩻O�Vr���m�U} S��u�k���4+v���ʩ�bĀ��}9�u\�K*��笋��P~0�)�O�7���&r��>�o�;��F����5g������n�c�����ɟ�=�*�������wD�}��І6����І6���Gi	�o� y�������a�D����RR��������G��Г?���������9:8$�����{HBX#>��m� L HFe,d �+�Y��@2xh-�9�1&��1?:�E�rYI^l���V�6��{��x|v� �s�h��K�,���*����[Q����ّiTU�������ԞG�8(�Q�P�5D@����9E�:�o�����,l5�@ +=���V���`M�Ef��#!�p��!A�'��|�/�C x�Ө�mS��a��
��?x���0,4�����>l��{@n>�z;��Q�"j/A0.聨]En�=�����#�� �x"`���4�:�,��j��Ƚ�a� �̏�l�z�����# I����C��'ULYb��H�є?SP0�ǧs�l� ������������[��{\�Rq�� c ��1&�Q Q�pk��~Ҹk�Je���$���kT�x��X�8�後�h��nE��b�Y�yf߆c��X}N�=�U�Sy{:����i?���qO[%$@��_��eD�
V
sh�n΄���D���S�c�k�@ږ5� �����Bm����b�'2?t<��#U�
��6����\PD�s8FS�x��dX>�t@U4TB5C�ׇ��܇"S��N�DUr$i�_����P�Զ�>� w*P�2�wvx$�+���l�k��nε����V^l^��͊�E�Md~x(g����L�>~��5H_���77r�Z�X�r���łc"O���t�x��kyV��V��� ��$#�sUr�d��n]KG�}�QNEE�`�*�mgj˦W5��K~>麤�;��A�;s\�Р���L���k~���Y��`N�"lߖJU:n���x�Zǿ-��g"��'n^���v�����=�=I��'PIu�>���")����#���t�����uJ���"��n����FrX�X����=������W��z�{tw��~�)���
?#Э?�ĲA��߻t���
~�eNY�J1|&�����<64����I��|�ֲ���7i�%��Į�1����P ��� ����C���V�A?D�vZ��M��2�5A 
U�5�zC�c��s���,��zŒ��Y/32���op?�s�O�~���F��nc�5j�٪�%�X�=I������}B��D��h�u��3�b4�e`yl�}�E"m����kc�}���(�t=���L���������n@湵(���RJ#�@xl�`�-�Fl
Aރ��Ȥ�{O����R�E��c�E�'�z��?\\_�ԡ�W�S����
��.�m/
#r�����d�1�<Ǟ_�*#?T��̓B���!�<�-�n��!	�c������w�Z����R��4֟��5\�Z�N�g����䔁�i�l�|�G����R��5EAU�1D^�:�|���U�~�]y��cy���n+�^����޻a]�Hs(��[��ַ�}c[O���o}�[��� ��R������ز:�TMIOc<����)+ԏOO��_Ǵ�x�o�!���?�	���7��$<8��� �@Jx�">�j��� B:Сn��� Cd���n���c<�T���J6�exp\�!�״���a����1}��� +�C�K���_�֤��`H�~V�'R�ͷ��sY���W(�cV���P����:`�{�eaP%j"Ҫm�GЪ�)�����1ϕ��"����a��.�
����ch�� �0�JV�AL���������4��y�>��w'R�Ѐ'��` ��T�ʁ�AK쫖}8:��#��Gk�à���>��U�����Y�<���j+@V��}w2��6�-��@�/�� |݁�Nq`��Y�9(�Uʘkb�U�5�_*/24�CǷ��Z�@� �1`�D����'�� $�Z 5�|�|��@=��q�*�@��`t���03�P	AVৱ嶠�XA6�W Gd��f�2���
{���TYq�s�^�� Q��$��>��	�y ���<�d:&�Ɵ�j!�66���Dq�9�c��-8K�L�$2p(&��$��:h���3��o��Sďfܠr�DaTJ���@���e��ߩ���H�X�L�j���g �g�RnP1�ʚ��i^[P¸�u���Z������r�,4�!l���c��ܥS����d˷��xHv�����rk#>7�� a�Gj��f�E09�pl`Yȱ�a��kp����Z�*"��W�م��]plM�>�'o<�w���<~�P�~�Z&�cz}y-7wsYm����F.^_)iu[�vP�~B��x4�),�8^��5�e����n��Z�W�X*rJE��amF��X'�3��p_�r}�	{��h������&q��b_C�;��������zc�l��g'�1���{ޡ�N���sź��!^;��JXX=�7+��~c��Y�F]f�dts�Usx�V��l���2?��c��P �g8����eu{�����:�`.���)��p"��]'�5�'���ߣ����;'�����<�	�Nk�6b���*S%Ə���~���$��X{�4��s�'/8#p��H��nʹ<)�!��K�#٨�8P��Zr���`N�&s�A�$�+#������W9	�v�X%���� �mQ���JA���2��+�X7q*�p�� ��W�[���9�k�j?=��D��5�{�l���ZHۿ�2l��aM�c�uXf�a����D���Ϭ�^�(��(�aX3�wč*�TN�lҢ��R"�`��n���( AߐL
}U&����m)+*?v�2���%hQ�����{�X�F��ڏs'غ���&]H{�.3�,�>�}`��f�Z����_����������|q+���/���/�a��~�{I��{Vk�2̝���V���G����'?��|����쏟K��ַ���__�	����o}�����\v��lFPd��+y���o�a�ϱ�R�������Ex=*I�pU�`X��E׋�Z�l���Z/7$-� ln�%�1�BU� ��y_���� �� aUh��U NL;�p.xx=;=p��ަ�^E�R{H�D��v�a�m�����d0�i3*7��'*���=�� @��0���m-GJ�h	�2�d(�3@��J�>�2��h x0�^�r�_Y-״j�@5<�{%s>2Ul� ���*(�_od��`�W�3d8v�?�*E9�P��C=ɕ��_�����6��P��g�쉎�%�(�4�!q|��8|��+��GT_@R����H���z��g��*�0���#��KWM8�� ���g��;��/�wWr����@G���P���Z���k�.�[T���7������Y6�ꗯ�S��� W�*��j�����u�t�u��{ ��u������5���/[$mi`OU��0�l�(y���{��Z�l����{T�Lc>*�%𢭂�
6FW���=fwB7f�PEF�[ ��n�vTd hĜ\oִ�J�N�Q��`�A+�5�#@�:\�X4�7��_lvvJ�2���F@�����
x�]��Ts��� �}�>O��"Q�!y�1�o5_�f1�XȌ�±��%K�*���~.���j�`�C+y�r"3��;�2�dL�|����13��``YNұ��,is����þ���V^_\ȗϾ���������U���y:��������{�+��n)��Wrw��=zU���_��UG���K`/Xֲ���vV6oIjg1	X������Gµrm��꜒n��hu�Y�D<�H+��3Pi�7����SdY�s��ئ��y���5||�0c��T�h�r�@8�
��&��Œǃs:��tI�{�^qw������ I�D��P	T%�j2�:����Ʀʭ��ՠ�{Wéҡ�2�|��5ɭ���/	^W��՟+�p�n���^{�h�JA.Y����!�e��/e�����:�?S�\��m�)�x����`��=	svv�)|0��^��'��ϸ�(��v�Ii~��**rU��8���K�\[à �K����0^��Y1��TXQuck3B2�Ѭ�(#�+Ɋ���2�W)�ݽ�JV�}	�{��P�f{x���ꕈ$ ��.�qi����t�mp��k�b���PP�]o)=w3,���ڃ�+�D������cW��k$JDڧ.��˗ry�Z?}�JC�r����ܭM��$F����\eW� �YC�h��-Ȧ؈���O���/'�Z�7@ģ����'�W��o~������R�\�A��S��^/A@����p�<����������_��������ZU�?z���{��^���È�E/ �[��ַ�'@�ַ���o_k�ŹF�4~�����?�*�At��#j�̀o�ó��v>��|��T [OfSٮ���{�$Ϟ=��z���U�U��bUPW����A���Nl���7���q �P݌�`��	L�3>�MEk�a>2�ѹ<�G�L7�v2��<���3���E������� �! �Fa}X���D�����8# �1t�Ԅ�eMSI��U|��V�u�`޲�Vfc f�}�oaD-�!��PV|;(-]52@���h1�+��4b!N4%����O_�V	"�!6+���6<�XPU@Ӹ�v���,������ h7뉊a��g<�m;��П�����PѮ*��N��VF9�U��=�����f{啝_%d��� �pH��wu��'ҍg|�s)�^���.ש%��*)?����z��N���Ɇ�S��}�ܳ�:$u��ۃsƸ��Wb���������`-�\7�/P���L	�봖K4�%�r�Y�nTa�j�;,S�(�j��S�D���T"����8�8n ���B�y%�Jf��WkQ���c[����_AFT��Ɖ׆
8߻��,_ V+SG%N�6;�%�B�4�3*d֙u��x��h�u醼�Md��G����6幡*� !�8̉])[ �FN�AD!�ʨZ�c+m#Uc��v5�W@ί��������X�CKe�6����m�fD^1'������Z�0uX7q�@|�DF�P��[�s̑@��
(�l6�a5a5=�c�)v+�|���c�=��w�Mk,z�� H�'o����p܋�V��̘�/rsuK/{Wg'3>��Ws����Oy�����&T\�k�%��b�VK &�an�K��@����-D.Ta��1	���㪪C?!#���T߰�=�)��i�V|�2�P`�pBs�<fAT
|��ƞ��DK����@�a��ڀ�ă�{���̀B���A�*!�[*��O��_��t�D�1Ys�:�k������ۇ*<���?\��������䄓3NPh0������PD	�#'�A����Tq�E�w��$�1_A�m7F �t����Q�B���!��e*M��	�̭��a��j+(�@d)	2�0�i_ƾ�
 �T�:~�P�u}�HHD��� 0�W�j&��#ɓ4�̯0�b-��@�5Z�����&�	!𺉫N	DҖY<s����5i�v$S���C��(UEǻ�I��E��V�%Dp~�Y�L�P��+�)P"�{-�`�`���5쑼��R'�x<�RD�M��],Q8�b�d�S�U0[f.'��2B^\x+��fvM�v��_m'�k���X�Ix���sB.��jކ�d6�'�T�����p=�}E[�:�� "kWbȞ ���Ev�rM�z ���h�>Xs`�{4;a���D��o���,V9=l$܀ǀ�M8��;����ٙ�����'OH�@����cPOr��u��	"�����w�ַ���o}���� �[��ַ�}���ZV��Gg������[�lw|�5� >�&S�C777T���<��~�]9��ឫ�Zi ���@�t2�m�mx_�Lأ�UzT��
����7U����f��F��p<��G|�B�  t�R�I�Mg�E5���<<x]�����>�D^����Ϯ̒#<�3D����*VT�<�r}s�*v���;p����;��h�p�` pq|v.��W�zC�jT������ 7IaӰ��`	:��U����:!�0D�'�s� ��:�-���k�WX�
p�vc�=S���Vs��p�z��� U��v���h̶��R����[<>��Q�k[$Bh�P|�?�tw�?�wv-��ȭ��Q�m_Q����" IWa�!�e
�Y9ɜ�p�ſ����#U������(PKEȈ�18���Ed�w�>�&�,����� E��[�&�Tt��+��\j��}sM�ЁE^�ؔV�0�¼���F��݆�k�A�UѬ�ř$�2���w���w��DJs/*�5T���-IL�j��3PFan��A���ύ�klCĲk@����� �Ԇ1�T���;�~@�@�d(�fK��J����J9X\��on���+�;{�G���%U��u�W�T
k��O$ׅ��<^䒠��\�>K8Ǳ� �2M�YL�6j��d@/���P <��6V�A���,�V��U��,k� �[*Jp>->M}}�ؠ2)!� ��8��n-��Jn�sZ��A��˲�u���Ɍ޶��>q�@V���(�>�S���N��~��?��9��x�
ƪ������k)����nN�2�i#����+�λd8�W>�.dbwT�@�|��Թ��vQ�i�Ϣ�-�{����Ah�UL��(��,�7$�EɅX�dXU��T��Ni��mؿ=�	�/(������Y'@~�-�:�Y,{���MW����W�����S�����������s'�}���nړ >��u����u��-�hɖ����j�C2��`�|��j׽�[ ��!���[G�>|W <�T�N8�F�ަ?��żK�	��0����FJ��b�R�^S�f�{E�����%�7��-��&�z���A���R@��9��E��������M��9�o;�IV���;E�:������'�;�j2���h]j֓8d� ��/U�i��h�q�k% �\����(5��KBuv�,����*���Z���Nj��W�����^�1����W���u��D���X#\�pLUXC����$_�2���螊��ڴZޅ���U����ۼ��Z��eb��b.�Z�D����$Uy����=�+��f_	�/�>�����y�V��?������pϴ���1Od4{S��~4����:�,�{��gѣ��ۗ_ 	7����r�[��ַ�}�[O���o}�[߾�Ƈ9_a"Ex�L�+����<z�H��p���+y��s>P\;>:�o����@N���I%Ex���ᡲ�O?�X.^<cE�x���Q��ܰH@�8�@Q=z�o����FZ���P=�G��o���b%rR�k��t�*3��^���1�G���Y���J>����g�ɋW_�k~8���%=Lو�ixxC���B����-׬tcैU׆��p.@���64ZᇇOTe\-��G�1�t��L-��@Q�YZp(P�L
�C�#QK�.W�DHݕS*	B���nM4�9'
��`��
V�N"q�	!A��T+�+�Pю�DX/�� ��NoX�C���l�k=��>9��E��!�k(3*��xԁG���DI�&V�7�t�ڄ���E
A�,5k�MG�F�K�+��ȏC��6�~�Ċ��!"{Ыi#;��^U��� � TP ��o_�� ^+8�]��!�0��&�8��q�}�65z�}�u�{cD-�F�f� �aȪf� �٬7����B�c��D�$jU�VNYNb1!$-`��i��(���t���W�Ve�X7`�,5��n�� h2���V�Z��LLPz0�y��:S�q�S�� `�!ޘ*y�Y�%���	Dr�2r�=�I� q ��@3>
Z�liu��D� TY�0�'���H�x���D�#Y1UQڹ��x#�Ϩ��8.Џz=� qk6I���:�Vf�2Y9�����5�zJ�y�x7��\�
���65��.5x^�f��p�ӳ�9��waϘϯ���\Nϖ� �x��>����d�-���/��D	e�y�\� �<:��;O�j~X���%c�W�����';1�?��' �0&��`�*6��+#U��p�i��2�72n��^mOBUe�=̝H��S[DO Ym cښ�N���K+���04�˓�����
�G2;>!YCk.���o���VN�tk��	P�l��d<" ��
R2�	X���N���6B=�֢�u?����!`�u�lk��x�ZN���|�v[.�#'�ݦ�U%�gґ�f}��&j+���-�������a��a�t d�����~Ɖ�7���22�s�zFs@4��c(�%ӱ���0���Q� 9��1�q��b�f�} �a� �t���^�O8Qq=R���D�&��n ���������
C�?U�a��fO�B�L6UY������觧�}�n�ם��5i�6�6O0��F�iJ�y���>��L������h����O��;y��5��`4��o*�"X\t���k��1���1�*��e�c_��0t�1As���$������Y%���+U����0�ѧx=�Q�|H��;wR)5�����A���J9��P�f�C�$��a�k[� �j��:�|��Ny�����ȹ?���؛Ӂ^?Q�Eu	��Hϧ���2#~�{�����ƿ����s�[��ַ�}c[O���o}�[߾���kTD��a������H>y"g��O~���w�+M��_����׿��l�+y��������7�7���V=���JOT�><=���g��~����x_�s�=1@t��pH���{B��A��O���0���r|<~.�Q�P���ޫ�F���������駟P}rt25/��6�D ���F <`H��G��3�d3H5_�nL� �����W�&�@�����t����t�߹�	
-�e��LTE��;R���((��jV��=,�������A4��-Uj�Ăҧ����B1�Ƶ�(�]
�%S���`� ����,����cZ���L�a�y]���*�g&je8\��@����׃ zj�����۞mg	Fh����ڢ����\�#�0_z�[�<��Vَ��n憸�W}�H��;��6�s�=���$��R�%!��@#�N�8i1����z��}	����M�����2ū���j�܉Q��Ħ�qⶳ>8�j.ڟ ��l�a/Cنk<_�	�n�msf�1�2R������N3�ʁ��I�|V�ZK]k.	,����ݵ�dݵ�i{��G��ZIU�����B��H��5U �W|��UvN��f�,���`�s��:�����f�Ϊ�ygV�+��@p-��Wţ?��H�a�C5GC�!�ڰ'T��uX_Q]\� ����;���+_�\����P�2�t�N�1�J�H��^ T�>EXnYusC��ֆ�f;��Jm���"���ռ��Ȩi�&T���j�� ���I�kc����qss'g�k����B.��y<�>��8@NH��|��G ��vH�)��w������v�e�9ɧZ��h2
cnH�ƕ���(k�SC;���^���$a4Df��ǙeM�>PrS��k[S�fm�= ��wr } �@p��U�P��T�IOJ2c��9Iu����l�� ��������� �rg,,�K���5�J�aD0��~mL:���h�c��6��gp���';����߾���ó0<�st�j	��~}sh�U�%Rk��[��X���	��}�5���]�K�RU�=��3H�@-T~���hyU�$n�k����㺉I{�;
%�V�����@D�vc8��s�pu�{� A���[�k�Ԋu_�L������Iܰb�M�mw��Y\�p�ҎE(�Χ����J��Ŕ��h��M-KkS�T�>EX�K$Gj㧤J�k
�6��rTE;��:֡�G��V�ix�6��P'��l~a�n9���b�pn#d�h�:�������v$Ot��8W�T��$mI �$ln+ل���/�u�q�CQ��q����_��:�������f�����������y��i��<<?��~S��VB�A���j
�l����r�V��[�<^'�@@�׫ڭ�loiVB��{��P��gT�:����/�4KB��fGι�{��� T�42��2���Q��e��o6��v���L�>�e�m }�[��ַot�	����o}����bG�C�ÃLʾ��w�g��o��wߕǏI�`Ȗ��{�72��O���ȏ~�c9=}�@i����8==����� w&�v������<;Pu�*���-}�AP��xE���ɱ�x`
� \ʏ� ;�X�%�Iۭ�N�?~�y��σ����n-��\T���G�SUn�D^�6�C����T���;���}^>Up�sq����;<g˛o����Xw�pl+�H�
s������4���M�@\ ��!臊9<��H��� l�pl��q�#����]N��(����p�����Z����# 9��������w�[�-�|c�*A��P�}��T��6�� \NȨ��`M&ғ����7*�ILe�{i�RC�����1�sę��uc��,/���*c��xSTM�����@��Sd0��
КG:>2�E0��9��l�ZaP4�Z;��|�J�k �h��*x[�ݪ�6��4�0�P
jnl}0�㸔ރ��,AjX���"vPy�.T�NA(�# ��䨫&�{��ہ/Z��
����Zc1.qM��K3�m]��п \��;�[l��Ø�	Ҕ ��k)�����p�]	�š�睅AY���20*|��ʭ�9��*��,ح�|��`L�`(*z�ő����[�e%A#�M�X $
@�J�X�8���0zwU"�8��QYo���	�@� ă-
�犆_+)�`�o̪��(����׋��.iI3	��T8�5�f����&�?�7(= �`\��</� �܋q�
kRm�:���I�&V�[�D�|���9�A�j�]����[�ޞ�q��jk(' �V��Q ���a^n��e�Ƭ$fvI�Ne�)��ֽ��S-m�/�Ӷ�R�?{�ղ?�!��Z>��S������H&��~Xl7˅4����}�p��З�y�-��?�3�����C%�U���a�����@�4��s>̏q8�I��8Y��B�2��dV�'��z������L�G'T� ��r���r�Jk�ͭ�C�߄cF�aoD�&a��Y֡�d�5`.��Z�ۆ��)��no8��=�^	����qus)ߓ{Fp7�^W�9\���I���w4*�B�< X�k��Q�lc����c'n�� f�z0z����=[*\KW@�|�/��?��A�o��Y%{�]HR��߭i���Z�� ��:�qO�6Oa̅��5�2�y�]4��*���nI2VS��������I�o�sU��\��ݦ����(�ͶO���d@A�!lG�˃�Eb�j�ᾨjTW�!�(�a6�⍙G�A�"O�B�MU�
��Ycփ7TIL�)�������m�{���GD��j�v_�g!@��*l�rfl`u��UB+���+��)�OcjZUA��N��S�Gp<�t�
�X�A�����t<�ޅ�v+����bۃq����I���|H[�8���U��7o��[�����7�����"�+���j�9�͕,�}�$�+�� ����r�� ��U�밗,`�wq)��x�P	��M)�QA�A�uw{�}`
�֙�F���Z����Y��?�Gߔ�o�)�lD�&��������z���Wr������J$��0aBi�����a��R�q}}���ʦT���"���9'�RI:�6�e9���!8�MU��DrQ�m�Gj[���
�@^s�p�+񷸷߮�Q����gó7��m3�2�q����o}���~��[��ַ�}m~���>,^N��o�ɯ��3z�úcv|��R��MX� �l+>�|�i ��R��H�<yD2U��/���- ���p���r)/_��o}��fQY�V�j�{�g��zKd��C�" 	�?���)Y����Z�������r�1�|Q����*	d!�<�ov%��+�h۰U��Zm�����_o"����E嫆@�=a >�6R��4��V�0(���k��Hc$��g�| ���A_�H�`[3�V3^"Z+�|�0�:�{4m��� ��B�F��29"�g�- x����ɔJ`�Z"�k�u�%B�/c��h�&� t����4��4ǮګFY�޲e��R<�f�/�U��x���|�;�x&�6R^y����U����y6Ws�z~�gp��5�W��R��j�}�x�yn��?��fӒXPU�Dq�x����%���N(R0��:^�v��v���c?T� @kl� ���眤�P=Pja-	�v$ ��a����-�g�� Q|&(��S��®����h�!����Y��̖0�3��5� ����C�P�����(4�[�wAv�ِ�z��0�i���G���F��짩���f������*�5c˟A�1Od�ށWa�mD�-U{�k�ui�ز29'�Yk3T��N �c���bS���I.�dP0D$F#�ױ�i7n1n�hh��#$j���5��Z?��u
��U��Y@<�]VQCu�UӪ0������C1�j%']h��3���X��(�|��e4�"�;O�[o��5r��d~{'�'am�y[(b�ABf"��{���h*o>},�?�R���' ܀�=���VC�cX:��96�F� �%�(���v��n�.$g��0X8>Pm���A�(տ_�+��Tk8~F�VDe��j�E��_�G�Z:��뫛nl"�VC�'�WT�*7�7����b����+�|L�1V�#:���Ux�x����Jv�}A��1������u�m��\O���q���\W��2N�8��Ҕy��R�V�g��9�=@VM7�>��u�$lxMM�GE^�o�'�y@5�ja����o��{k�ap;{��$�笐l�	ye�T��ȾĲM�ZT��-�](j1o�T�x�o���:��-�����KT�����j���{�����Z�Ge��O�{�Zm��h��,�ڮs���v��-�z)�T #S���J(����=�zi���p�櫅�-��Frtt�u����|3W
ꖸ�wE��8�Ə�Qo�V��Iǂ��P�T[U�VP�6T��=��L��6�L@���}u�f��~���m���pl�T`ll6+������((���LNٗ�~�	הo�����#^�u�����syy�BV�m�@�c��9(�����w��d6=>� ����0�^���۰6���l6@�g ����܅����8���ziJ쿪L��Z�D/R:����kdE�$�Aֆ= �,F^R�w�x�B������f)g'3�[��ַ���i=ҷ���o}�Z[�])� ���S9=;��ь��
 �F��n��꒕jx�Beh6��tX ̺��";D rxp�⅜���IxX}��76{yqI��f�$p+�����a_��:��y����t�a就�ϗr4;" ���ۛ܉�B8����Ε��}��!m4T@9��jy�|	���X훲��=�2_�����lK��c�|ă�x6���s��FZ�G�Kxpfq~�U�V*�_��@��iO�j6 A ><��%�Ӂ�A)%QjfS @BXe�	�)��b\ �i5o�����p'N�.��6���@b-�\���[� ��ңIj�,��gҁ�[e�{�0�kB5n�P��k|H�YN"�--�"�D��l[��a�L=V�%��RA�d
.�$!�p����n|1��v6W�O{_#��b�H���o�wn�����n��VN:@�d���,y��I8N�x��SB�"���R�������*�4� 7�y��wD��
��)���Z�WR"i�Q01��J� Xōz���;F\�-��S#2K��G�5_�*�hs�(���O1c^;�U��`� �X��k�ʄ" NH ��Rsw�����m4� �E$�<�$NY���r!��0rHɽ"��n�rt4"����<��l�k��be�\s�ej����`�ʀ��D��Px �wp��B��"��$���ZIǡt�-��ްE�pV-8��t�*}�"�M\�ʦT{2Qu
��%�d�2����>b�U���
�b��Z��9�i��P�1��Ϲ���S�PT�.��7T�]\\�O�hn������؃����Vl�5,v�k�L�	�.}svr&?��ȗ/^�o������&���k%��1����P�rI��*jZ�`|@A�P����ۢ��,A� L�>P$"!�\*_��V�љ�o��i�������(� �qmisEa��ym��A+Ì�2�]���ɔ�ȡq�+��ҕ��t��O�+J=Gi�c�:�N��%�.)�1�B�uT{摯YN�z��f�s���55�,��R����ß�M!��Z���A,�1�d��a�ScDOed�[������R��qH��ܕX�%eg������~����1H�Yñ��JUfA�%Q����E���N-cb��vǘ$�gpq,⚂,a~�`-Ś����Q8F�TE��`l��{��������f�X�N�X�JK�B-����QUbtW�06Qˡ�F5�p�k?"��6�:���0?b(���0~&�1�P+(`Lq�B	��EV2�dGV�&P�2W#���mX�O��{��f{\^�
s�ۼ��؋)8V�a�b���_�{��BU�o���~��\��{����J��c������-mOǓ�Z���q���R���������&#�����X��������+m����}���<��{uܥA�<�������.��?��_qLz� �8G��8O��a����I�_?}���J�������y���䍷�w}�v�o}�[����k=ҷ���o}�oE.} $�ѸL�-��HvMEX�����������ٳϺ�5����Z��?������rws+��a	h�����#=�<���_�Cjx�ݡ�;yyyɇ��T��^9���D��	 ��nXt�Ӆ?1@�T+r�?o�������ǐ$c�c ��n~��bAPҫS�BZAx���݆�%�n@P�`��gfU�J�2�h	�z���P��*I-��7@iU�E�.�d@y(RP���F�+�$Y��F�`Al�W-}�3=7C�%��1���������t;��PMq�E�����BH@����|�����'8������>D�J:�$ja�a�8g������q3! �/D��b7�@R�ڇ��m ��'��I�CBk�����C��!��K��:�	�]��y!N�xճ�~bk�^����A�h�
�jJ����N�.�-�CnG��� c�DK�`���WG�d�'ga~5�s��(&Y�Ъ��h�e��M��Wl���O;��hvY~��f�b���u�⿑#��󔚄�>�(C�A\n
���i��-�E��7.�ݚٴл�`<�����lC߮!�`LT �U�3m]����$r�T1��|��o�Oo~�}(�ʪ�e
 �v�����r�*}��YP����]r�܎]A�~���^:TP[����!�]����Z� yű�X�,+bƵ ���h�\㠄A�/��*��U�_ʥ��a��������V�#��B�|�XUN��V�P��<�=2�rz<�i�/^]�9>$Q^4����ZU:`�0OB�z�fZ)~�����G�dc�|�ͫ�rP0��p�Aŷ�O���T�AR�RY�S�㳱�$
B�=Q���d��e����@W���\\ � .]	�JK\���{'�g,��m�<���Zrwc�1{,ϝ����6~�믏/_W�ؙEb:��J='K���~��`l0\ݬ,]5�[��uҳGt.W�T}\w��d��I�><�-q����̔�~^��Z�W�#T����	��=Ţ+��I֛y1R��C�k��[���Ƚ���V���舓���^�﫚$v���
3�����������w:�;zܡ�q��#�u-�بl����s�@��'��+p����Mµ%�M��YqQi�
F*O��K�*�$�ǖ��8nCN��/kU�U*<!G�eW��o�!'a��~@�>������j�����U!����9���S��npI�4̙���>J�ET-��L�J�0%�\���w{9�Wb����U�����jkX��EV�&��5�n�|���S���Kd5��~V�����������@R}��r֖ן#��M�^P�da����˼�z��ة�{�{�0ڗ'O�u�ʲn����o}�[߾ѭ'@�ַ���o_K�¿J\^ ��i��E�|�_�z!�����?�/�?�7�>���1Gِ6��}���OTq<y�����?�1ɏ�d,��5�MY-�*�A�ψ�@?<��|�B���<|���),
Xq�Ҋk�t3�`(g�2`�t~�`�0X�� L��D��x>������T��@6;>�q�a��bA�)��}����<�<�H��z��]�TBr�[u��ח2Y�� It��hH:�?K��F��!�"�ڡ`e,*�+S$䴀P0�fE�7���bD �%�o�h;�#4pw�B���S���[c�%��<d�O[N	*_C��������=��g1?c� ���P�������i~ȏ܇�Y���U@��<c�8 ɏ)ڈ�����Q��pҀ��`�{�g�8@�`���W�` ��=)�B�ESZ��޾
��VD��a�z�{Eǰa�af}�t��}������U���շ
�an�T	�̐� a�V��
�y���cN$a\�����#-�P�߶;�N�q(��^�К  &5 ��-\�jS��'y��*J�<�Ow�C��Xl,�g�7�qJoi۝�	S��E�ٖs��J�DI9T2w�:eM��%�E¬Z��4�'n��k`��h���0<�$�b���x(�:2!�`|�ZB�qX�" �0�}���*�k�{8o�j���M�)?�6��Ъ��)[P� ��m���X˼��bE� =�)s4lN$������������8���J�}��i<�{���E^�#� h*D�z�oK������> �h�o��b(�7׬R~������y������o��Ɍ�4�h���hk��"JI�a]}pv"�~�%m_b������h�T
c����j�L+�[U�1/��t� �h����+�H�s�&>	��S�oȆ[fU���,�4d^��
�a���L'
���;�A˳�CёD���e\B��zg�gE���I77E�P[�&-��cX��0`����i\{]�-�@40� �U�G�5�WN83_f�J:X��r��~��:\�;�!��/7�>*񹞗U��N�8���j��[�)�by��70_�S$���/%!�u��ye�[��7|���"���c�����$?"%�v�{��
����|�1(V����� �uQ	�%��-+���Z�&�d��J��d<�<�x��[l:�2�{h��X��8w0�/X����qԑ[ ��]%��,J�����$�S���b%wCU�p��d��H�lq/iF�ψ��$):b������3թfY�Mkj�!�ev4�T�{<�7�=��38gXӆo�%�{�����gr||��a�-g�~��������X4���_)�T�.:+�00=�_� )����׍D�p½�Fi����s���)_j��~)�^��l;O�������ۍ���b�x��K����/n���gϞ��?x_�|�B.^^ꞏ�#z��1�{���#�	{%��K(�
��Ř$Y�}�H��W_,��]������\�ַ���o��� }�[��ַ���xP!�[w����������ߗ��o�V���>h�> $��W���RTx���yx z%�����o<�w���<z�D��<��ё��C�S�LH�z ��^�'"O��*(�t���`h�.� yswÇ/�q���$�v[�w�* �g�T��a������J�����U��|��
��\.���a�+�?�M�Ö��Ņ�CNg3�c Y+X��?���W<� �/=X`���0	�vK��tյ�������5́�C�6E�@��%�r#j%E<�v�����,W�E���8@R k1`v�[���p��8�j]ɏ�PR��P��Q��a���ӫh�zׁT��9���]�r�f  ��EG~�%�gg�������B�BɌ�`��g�*:O���
�U�{�Jk������W����~4�.*���-�\�`r�U^�5��jJ~����l9�夐�/�k�]�|N6�_[�6J���@3�-��V%+�����^�T�
�
���x�כU�[Z�A��q�;7 ��c5q�66�{oӡ�ت��B2���J�mXw��'��{ ���2�ck�6��p��@�/���ۘ���6�Ih�u"�kh����M��q$j��=����i�S"d�N�0� ��s?�dI�l��6n�ʁ�
=���$�o*��f��c�|{{cc��i;��d(�ɱ�1�߶R����аt��,��+I�XsZ`��\��2/ d���T�M'�\q�F�����YQ�дb��L)�#Sn�TN܆�e�Le��3,~��qts�Z>��dv4	{ő<zt.o����fJX6�6����'��ť\�1� Wt�F�mI���Z��[�Pd`/��R�
�$j�G�8���T�l��P������*%P��q�߁\�l7�Ǵv�k�z~�-��U�cOT�d��)礫���[��=� (p 9���v���+&�nmDcV�����j_�Vg��F�;��\u��� _��>�[����vX���=7�J�Ҵ[S�0����Y�:E	ֿ�Ʋ���7��K]v�#$���j�Ղ�ց��g�Q�6Wi��Ģ�_�S�_yڑ>���ߍ����`�BK;�Ȟ�I��D	�ϙ+dD��PP�C��pv�Z��Q
��
$}f+s�Z�K"�Ì_J�@m�LMBcG����΍JAw�s�G6Vk������kE��BJ��K~��:M�քy�T��"Q�(�A8��p����F���@���`���:�����Mk^�E��m�䵭�D�}��k�óc9
�ס�Rv۵#����ꦵq��+�����~����O�m�cǞH�%�(+~�U�.\��FƉf-��-晞������ɔpγ�XN�fry�J>�����r�D��؛A�*1	�[�u��/�}���s���O�6��~���Po�Z��oI�a4�С�0��0�,����T����

��m�o~�*������w C�o}�[����o=ҷ���o}�o9r&b�ޮ�.�>�'�a�.���~훭��d8%PD���ɗ�~.�/^I �TkI���*y���G��+�_�b�$��X���C�g_|.ǿ;%p��o@5[�lX��խZ�y��S0&W��%�V�\ ��M��$n��׀s���Ŋ���c�d����x8�����纺�����s�܈����٢���y8�8�<�Q�� ����+��ǌ���ه�Ղ�ä|�ժZ���Y���z,s0�%Ƭ#� Q;�N$�R=���򁕡��<�`T���-x Z����$jX- ���l!�[%<V'Z�F�|�i:�l�,B!a]��T����T��9��yPe<�q7۵�UQB�)Y��AiQ+QP��- ���
\���.6]%���A''�	o�hN�b���� P�k��&��H��]��Ս�-��頯:�"Q��̤1^"D�4%� ��~ǚ�_��3c�Pp��` �nU��1f���{�Y��}��p���"T	x����o4��Z΁�w� wn�0ז�'~B�����F\=rA+�����e�Wh	��,� ���,K��)�ƿ3��D�s���j� �Y'2i{�JIk�T�v� =���6B��1 ���A*:Ǯp��ݭS�Ū��9��1���N�hXnv̵hw�����Y�ͪi�6aj��e�s 11�*U~(p�PI��i�b��È-U�Ԭ�w�kx�oUmÈ�ؾ�>Bf�@���"�$�3��r�>C�	:��a�e�x�n4�ޭ� ����|ns� ��쭍��Ȥ�2b`_5��Q�6������gH����$�m6�5�i~K�����l:�{H�6�B��ʓ'O���X�Ɓ�iX�10##l*A�|�pa닻�4P;��L�?����ܯK������2E,+ ~�X�R*��{=�%���Zlň�����&\��^1`�'#�������=�_!��#$p=�8 �>̔� �\p��X�'3�F
�z���u��#����H��	Uuj.�(�����+ʐ�k��E��K���U`i�����T�{�X�AlW��f�E��'�A��:����׍$�}]�����#m�*K��!�Ҷ���}c([���U�N )Y�3b8ʥ�"''��2d9<��%�$�k�)�4��%{Y��k�B�$�-�ɳP"�2�\[�q��J����
��\�P���vk��𥊛%� �N�S�������܀�h��t:�<�q*��?/���
��]�žm�j��=���l��e9N��ce����z�
p�w�n�h�
Bjd��\^q\����;�?ٗZ��BQ�(��utzB�#�Z+
��ýI�<���Ӊ�v������dz��%����ևa�1�Ջ����|��GT{%YL�+���PpW��)�>��cy�2ܳ�������<����'V"L]�h��������ժ�&�Q�B������~���g?���/�����o}�[����l=ҷ���o}�o��ʫח�~���d�a�k���	�P�eh�o���D^����>�H.^_�Ul-�r_��*���n6������9+MQ8��
� Ղ����1��l<�y+)c��D ��T���,"��T=ć1��g���Y��7���v����L	Z����˻{�T�wW@~  ���h���������m��
��������	���Q����9��Lہ�꩞3�עlv����7�U �:<|��5�1��*��P�E�g����AN�(HX�H�
�C�]XgC�<�]�����1�Ms��p����R@؊�d���C�5���h؁�U�Y����6���^IK��*p��. �!�a,�z]Wk@x�Z2�Ĳ�h�!*�=�՘��y,�Y�-�7be;��6\�eGT$��2�|���_��|�ߢj=O	��=��n'��#�2J ��r��f�������c�@�A�K+�傿�]�x�� 	8�����1�1��mg5k8�@ `@\�uJ@�,�p���J�&�m�{?�-ㄕ�v��e�XP���	B� ��簪kU��� � � ?�U��7�p2����>P8��i�mC���R:"��pq4Tbó���4��Vwy}u-����ո�5xI��k*�5����b�p��6�Ҩ��m�8���+��scVx�cf��Gj]Ӣ(�gz@iF#�5`!�ɝ���+��X���k5�tJ�;�y��yX��u��!yv�a,a���P��סu�-	|�Ӱ�cG5x�Q�)���Ǔ�����r�R��"^��zC�m2�r��q��Y!�Z0͕E( �7�̸�p�B�b��N�b�;J�b��sم5�s�c�!T"��?rPjR;$��d�`D�`���Z��$��؋>z�{�����*h8P;K���nE�#� i8�u���Z%�]�6�� s�,5����L�����fk����� ~����^�k�yg3h�'��6	�BC�S������2��w_3�?����\��,�U�=�^���*��r�)������Nz��Ͷ��)V�YH���D=�Ȣj;B�svgUԁ�i��V���7����=��5���9���),���9̯��uI��_Of�`��*
���?'pIVq��1l%˩�����mdB�xP2����� krk�Xoc��srySl�]��⭰�]��?ӵ��� ����{���?���F�'Ȅ����g$D��E���w|=x�嶖�|%w�s��m�Z���3%a�ZI��6�I���*@m�c��N�ِ�i(�˶��L�N.�D��º�{ݰ��-�
{�@a�@��G�@>��ð6�i_��}#�[`W6Rb2\޷� ��������$r����!���,y${E�@ Tr�E-
'r#lPT�
�R����f���������K��ַ����z�o}�[����4T����͜��`�ml���g�O�8 Ѐ����[�}x����ǟʯ��r}�Z�CT�����j�ŋr|v�j`��jҌ��z�� R�rˇ7�#�������/���F"l�:X����C&�i����q���W#��O��trD@��#Z��۟�´����A5�����MY��Z����c��?��R��@�����ꔙ��L��Z%���ڬ�#@_j�nF)��XA�'��6_���T`ʵ�@% �d��R�b�A5�9hK����-AK�WW��� $K�����@�*��� �O�B �6�p�X��໊<�����w��
]��ǃxYi0.��Cb���I �@*Z�r�;�������D�rAe��P�4iü���¸ ����>�Hi�*o�J�3��
������a��S_n��ǲ4`ǣ����[\�����@Eu�V?nE������ު��D�/䭪}X���^b%��@}7� S���@�p�Z0���s�_� ���*��{�wd]��f(�'�]�
k��ی��6ˍ����faF���(�����:���2=<K�w�OF�� @f4�+��:y�G���
��YԮ7kZR�΋�~1���VU�����0��a���o�p�Y�����z�5HZ"�� 䍕���Ι�0�k	�H˱����:�L��F���l*7���j�&�H7� ��%�F���n�c���Y1�ev\���<
��hpmnd� W2��2��ɴ�I
��"x���VG�#	י*���,"��"���
{
2��'觝�3` ,p ���� �����E����#��:�K8�P��B`���<�}�0>���on	�a� �*aU{م�ú��t��R��%�/����>��'�[U@���W#k6s�	�f��-�XIQ7j���8~]ro��,�+���'ƦF���"+Ɇ��4�'O�f�k�\uA�T�X��`;�� ��� ��w*U��ǂ���1R5$r�]w@����A���-�\"{�lz���%Z��Q	E�#a|�2�T}��͖�!%L}���h�td����Hm��~��h��g愽}�����������	'b`Y�Jz�+A6��|�7�YP�>�L��x&ӣ3��d����Hb�Y���G�~i&��屼�7I�-[T��*�m�@�$X/8���-3�j�7�XU`�Uw`��P�`��r���%J��=���%I�|�!؋�ךq�1��5�}�%*Im�W:��e��a��{�����J��� w�,���_}��v�Vj0Xv]^^�k���]\s^N��p����i��<�*/�o���6��OH@��?{!o}�[aΏ��DI�M��1$����x�/z�1�18�8F����ө�L�`��ׇ�#'0�L�}$G�������\�����b���لsu��T�;��LIr �)μȡ����(�� �Hp�=s_v%�k�"fI��|4VE1�r�M���m0^"��L�����_�/}�[��ַo~�	����o}�����ώh�����k׬�ժ�V����CV��on�ً�	1w��|��Y�	�Ǧ��I����$�rrvL ���vG�m�^��mB��Nn�
�� �z��
$�������U���yc6Z��F�(8���y���J�ix����i �����rqq)��?�o�����;@E"A��*ᤥrݪG6�!#�jdu/���	���*�t��u!��6E5�����3�Ԏi8�^�`uDP=%p��K���l�v;r�Ҫb��;`��B4Rܲ@T���ʂ�}Edqv���EPv��_����:bd�?2&�?�Ic�U!'|�vr@�Kn�$Ҟ0���+@@��TC<­J�������L��l�ԏ��l�0�5���N!�|���0F��#�\�1�d���E3W�X�:�V ��9��y[��!{�Yq�|���b��"�Y�$]�W6�:� s�0��;���߃�Q{%Z8w7��z�\�X�[#��K�,�0��*�s��{cv�B�rXsz�85~�(;���� �@`������Z�s��p��W�S�:�c���Q��'���]�TmͺL�Z�!kH��ؓ�j�B6Pe�q�Ж+VS��s�Y��� ސ��>iA�T���2Xx-ɩ�����Mh/S!��� Z�^���X���~+#d @MW��5G��qT� ts�s�1�hf�B��q��<�f;A%F�ֈ�^c>Q�U��X*�zP�!#ȇpo�a%=��b;�x�Ђ
�)���z)h]��V��,wk�̈�����=`7jGT!������xż'�Ky>ұ`j"d�pL��?1��O@;�� ����$�~{ƈ`_�u؃�ѿ$_M���2��#�z�sq]�$�H�x�΀g�)�;UR��FJ���Z7J��A,O���fU���U����$�>P�*��������"B	�}h�~^�e�fS��ڬ�lM�r�<��P����Ao'y٧[��Acl8�� 9�e[�ܶ���n��:�t��{�`�a865�s���ć�����*sEܦk�4��&�����p�ð>L��8���|e�� t������}�rrr.���}���R�����s����4��e�pmk��%U�_5I�R��XT��yR��P�4l��d��&��R��:�1TM��n���玈�r��r���u�$�!�Q[!E��.�����Y˩$Q�:�ט]V��KmA#�mG32��#r'����r7>b�γg�hߚ��),-�`þ�j������A����:I�)
 @P�.0�)(J@$�Ę�/J�Ϛr�Jm�~����g_~NZ4�u�W��}_l�׹&2[��Fb}
�D�fW�g�3��w(O�>�JX�v*W�U7���oZ.��C& �Z��c���JP�!8�h�#W�	 }�[������H��ַ���_���8ڃ�c��j	 9x�{������������x�J^\�������"<�g��ӳGTm���?���~�m��F�r�kT�%����X�[U0�LxHk���P CmD"�P�]�_uw 8,Y]$� ����G	,\]]IuW��o��&�� @����1,`����Քx`}��[�Yn���_���o�n~)�PC�i�P��❴�� �N�� �Z��:A iK�*c��ǚ���m:±Zݠv�MX�> D0�$ 
d_��|&��*�*��!�VAV@��;竦�8N~ �SDC�#�
��U�eZ8ӓ:���6W%���0����|�`8�Gf0��*xZ�Eȩ��``�Mj"�}�wh�V�:"�n�zo�e@�ۧ9�r� �!p��s�;�=���Ċb�ɎC��Z�YJrY�p�UR%߳�aM(,T��	Nw �A@0� � �A�Kӑe,�]��@
��N�rE�J`rl�i��Xmkv�����pj(_�:n�u+�1|I`�8���� E@�V�k���� ��D4�ch�(H�ƀ[�DeH��3x0�� ��װܲZ��x׫��h�+��n	�I����\�fO�Rx2���J�(�4��j	�j~SmDV-QevB�_�s�H k�-�{���������*�ql�ꆿS�s�Pх�,Pw�&���Z��X����knjk>�
}R��������c��W�3��̵f%�Y8�®���9��y���gJ�ЮI�eYl�TJ�VR�#�v�`�y��Om�z�ﰕY"+h����L�̭@�>Y�������	��բ)Rc����u�q�:�ʂ����%ρd,��D%T���� �c���	�c�iӁ���
ǆ��+�u2�7*;�ܩl]HԎ��ς�+̽��ھ�4S'%���;��/�CLu�k2�vjOE�3(+��&�`Ө���5�u�ϥ���7�.��.��#^��`l2�ڔ{�)�4�d�����T�:� �V-�#�l�/W����s6�e^�y%n宅q���+]��|�}���s�}���`x'h���c���#�1�=lvR��9ޜ�qUt� �]�b1�qbN����ӧ����V^_\�j����	{� i���P�����>��lG�J%A��5D�7�J�b
Vfa�c�N��K[��]$�Ŋbo='� r������Db8Q�������[��{��3��f�{U���ڌ{+X#��j��6��&�U�A���z-;�+Y��$��Ǐ���q�!�J-Wc���Kؗ������=+�5������,Wk�w���O39�Üd�n�����w����)���_��͵����v�"fy��:X�A��Z!��7Ԏ��L�C{���ٟ����g�����2g�ޭe5_q�r�:�77W�w�w��{����W�.I&��Fi� ���*�[��ַ���j=ҷ���o}����A>`�@�mxhB�����2;?��G?"�5ȧ�}&w�g�R��|�Z��`��e�����?���z��gU�+��B��{_�z̀L����F�,�cJ�}y���>���o|�������/6|�����ʜ�y>�.�Z��Zu��-���ʯ$c�.��P�6e�����E!@�?	��Gf\_����	�?fX�@��2H>�g-�x���{�.K��:���ΙYYU���H�mS��^�˫ZV������~���Zn[MI$E	aL5d�t�������ŽY )�EX��Y�yo��9g�o��,m `1�U��u��r�4��p���H��ʬ@ "O��*�Ճ9���o]�z��HE��N+�Y��h ��րJ Kj�D�?�=�!
Zk� ��$��A�|iR��GC�>�Kx �	#J�Z�8��r�a�,��׍Y��:}��?"�e�?+����������A�jpU�[������v��0����dU�]4|�������Qy��*�=��B��im��;��Y#���O̺*�� ����T%��?V�خ�T*{pqf�$�:'U�*��
&|Fh
b�ϭ�A��ǩ�e�9�B@��)ǥ�+a���F.��-9Tx�S�����lo��P�jY�QĿ�{c�J�8�I��vj��؉�c:�HռԠ��%5u\���w	��,�I�ܟ{��9H�B�T'���
XW�]�JJ�3��9�֔[�$'�N�0�i^ȍ�߉�έ��2�� X��a?ރ�a��"jGeVvކ�%Nhk�}�$u������)�V�܄��z���ʹ�q��SY6#��8��Җ��sھ��������`.�~���͆s*TvT���,�����VC�¼���܆���	�b����^�μ_���e�/�=~�)�����{F�u�`�õ�l���;�p��.#�1�*�Ցy����\��{�>��:;�T�p:�Џyߋ�MU�0��d�U��uJ�*��p�(�%�gȃHu�>נ�Hc�� ���:�/�#��A|��z''»ZS�8��_#NGw�p}5c�����CN��E� �w�ߎ�,�������Ɍ#���fsr��Ӊ�>:�Q<6�O�!����p���Q�+U�x.4|ysˬ�m{��9; ��+�s���3Q�0�"�����ִn�������ѣGQ�>��ҋ�'�s>��y㓏�*�&�;< �P� 砨ZSx�'�c���~p��!A��gx���I�9R�uD�l����)��C�욻�!i[�'pT>��PK�Z��Z��YX��si�Y��Ă�D	��w&���
��ۛV��"��a�M&T�m�;Z+����j�Z�g�4ُ֧��d��뼯FF�3�*̭��B&�p.�����%ej�~{su%�z������k���0�����3��8�'�2�]�T�����e�H\�7^S���ߓ�}�����M9p��s�x�����*%�o׏�?d�K0��}���8㣇����X�mlc����Fdlc�����4��2��"09�M��8GU�d�q��Z.�y~����ߐ����}�uY�洌*�b���ɒX���ÂV�=��>���'���'����g$X  ��]�V�w\� �[�",=zLo���N^x�e%����	>[��v5$|��ɺ�(��Z.OOW�b�Qc5�b�d�:uY�"x�������W����(?y�Y_�����5�C�W���c@�����d l,ܢK�K����Vg���\�(�C���xl#�y�0����4�k��}fm$Aˠ�d�rV��;rV�i��2@�E~A9�̊^��̄�-b�w�	�8 �! #R��SP��ѾK����vՇm����Qr/���z�q9���"\��Q�6&x�N��  ^|U�Jꢖ������}��(�?�T�3&)+��d�=��V�٤0�A���3�EkBG _����r�w4��b���D5sC૥��r{��Q`Pmr�����@��	d�W�qE�����̱u�n��[��Ƥ��f3�|�c�7jR�*V���j
���ң6�3 [�3�0xS45�?���� ���N�a����N�C��@&�Z�>�X�;��a��,t:��EC_AHb ����<a�c&�W�dYKUDg��m��$Y:!!�1�}j,��-�@��:���±�z��@�$4b����p�a���ӌ%�����~��h+�~��"#�؏#7�L���j���g%aF> �s���Ϫ@�( �.%A���/��1kQw���Q��/���5WA�RvQ��)�V��'���&�@���b0β��*J��x&��Tf�%mf�^\p,��	ʸH�/d\^=#ؘf��O=����z+X��[��L��^G}ԩ��*�f(2�Jʹ�=�Z�6d	l�D�R�Y�jɶc���zdv3�5E�����:2���A1(-Z~v΅,�FPv������[Y�h�8�.��G�h;̈́"�����V��P�0�}�m,/g�|&�Ȑ;�,�|��2���^P���	�L�7�� �0�ʡf Y��� NH�,W�}�w�@X ��̦�-RqgV~� r���Ε/N(:qrl����W��&,0�����02�D�A��}�]���=82�fx}Ե�g�K-_�yoq��l�Y@xN	�  ֩��RV�#�ɓKf�P������\�#��<%Y҆�K���umc��7U�"'\�c�3�>�����j�1��j�5&�"��ڂd��C#��THίa������M��*"�@��I��3},T,��$�<����D�C��7�a��D��8���c��.FI�����9$Ϯ*�OC7}��F��n�&<3�/|��_��/ܗ9,��6e^���-��s3-��k���VD�j�\ܮQU�� �}a�zz�D>��7��˟�����~��)��>K�  ʒڟu��ރ��3I�N�N�{�����������jl� yB��:'��E�Kj���_!3�ZP������$���Z:~��7��_�R�6���ml_�6 c���6�/��f��f1�踽���g����>,0A��(/����PcX��{s D��r����Je�������.?���#�I+��(**��0����P�K@>�1���������"�v1_țq��8��" /��Q�i����F�f���A�����fjEo��Y@�w�޻��O~�c������?��<��qX��#Xz���
�w�g�,� P!�OԦb ��PU � vJ4Rj;��	ۉ-ؒ��@l���9H�	Щ:�1{��|��߭J�FG@>�Mi��)�DX�?����g,��<Q�&b�	�W#*!ܾ	��T"��E�V���ߵR�� A�2WAÜ�c0�[C����&��(��Q�|o�����@?E��[�8��6)%Q� �9 �Ϣ���5�:}Mf�a�fօ^8�K�����<f#��'�hJ2 jX���ɨ�wP��;~��xn�=^��CTm�W�����X�j��*?����sے�Y-HI��[�"�b�ñ��*����W�y�����
�:�	�1�in)���+Q � @�J�XI�v o�������n��ծ���J�}��<�[�O�X��ֱ�$��n�^�O�*�/(Q�6��}M�3a��i�{�V��Aޠ��V8�'�KV���B	3,��6 ��V]?X������SGeFx�p�t�ov~�8�خ�}��U����TF�6�;�G_)+�Pu��n^n����M�S+�{dE��
�P���1�<f��$nTE��@.�uY
�g{������SZ�lv;9!�͘���}��d)����O��Rg3X&�����S|���$�'���1��r'�O��$<����ӌD�Į���8�ISy�j���$(�C�-(�8�Qѧ���+�,�d����Ϙ��Y��J|���L\��k�����$�����1�n��ԉ |G����J�k�x�oT�sӱį4�GB5:d\��U48�y��'���j�c"���*ݓ8l�hs�͟�J=�N�@�����Nv�?/���`�q�L>V2O�a���J�+��c��.���4�C��l��a�;�|�HR�Ԫ��8W���gO���G$V���������Z泳�����7ސ��Z./�B_.�G�*J�*�c ��#1�\�IA�)��L��sp��ӎ�/<;��p��u�ۮch8���s����(��t�S��EVXw���9!�*k5���|����O��R�QА ;�b��ZT��w{�٫ben��}v���/��<����^��٩L���e�e1a�~OVrO�(n ���
�wf��3-r�6;���O������[�������hH*(��خW���d8��[����ԃ-�o�!��η��7�B���r�j�f�	��sUbCu�簈�a/���((X��xᢪPb6ᰱ�mlc���3���6����KmX�.���-�~��x&���]�!���-!2�0X�r�c{P�n������h������O�S��~��oXa�w��?/)�g��L��x
.�2�����5��>!0zvZ����0�m�GZu���L�_I�U�(��ԓpZXa[���I h���o�����/�G?�{yz���0�m�&��
Ǣ;����e��$�/]��WcZ���������H��U{%MZ�jm3e%=+&��BJ;�Ԙ
�s�V��ss%���@��F1�T�ö4�7V?~Z����V�r ��h��Ƭ[@�h�gbU�F����}A`ib��ee81t�q *r[/kkW�{8�6b�TIP��{�d$���EK�q$<��7mڰ�7� ��Ԁ���^���-ѵ2*z�b�I���p�d�*=j����F!��dV5�� @��rՊ��Z]��l�^�v_Wo�҂~�UZ��WU��y���
�{�[z��	��7�) +13�����C�6�zfO�r� �b��q}�j�:��UШ�E~�6��ꨭ[]T��,��/Qy�J��fT�q����~'˙**`���o���,���@TF���a�1������)qR^{T_�v�l�Jn�{��4����@�hn��C�l�,�����"?g��b˰M���z��T�=B�1�6%�s��Ek<�u��ծd�5�y�׃B,%�b!�Pe�&�Oz����U�C��ްB�Y��#O�˘T��#�>��%H���\o7n-�'�&f9c�6����v��L����{��fC0�6y�lR�[؟^	�j�p����T�:7_�^K+`]�{�����ݾ�'���a����
����y�1'���J ��W����><A J��Di�\*m�l�$����td�g/9́���o?�'�h��$ �p>6�h��h�|�|����B])h��Y��m���0s�/��Ԕŝ@j';2�s����D�J%�-�_�S��I4��X}� TZL��͠�����B�r 3��yc㹋�Sc1�$��`^��ا�\�v�]���fΉC'���{����2�B�Gqhx�齀�Wb�&ef���Y� �������9$�,橎�>�PA��T۠H���r�a8�wT PM�7T�r���32�"�s	�ʶW;�F�D��V�o$�����v��.����M�y����Pm����:ӿ=�~ �$H�q&Ukj����B�"wl7THb�Y����c	�@p��d�O�Mg���R(6�0�y8ƽ�#ux�X�;����Z�./����&_�-Y���8G�����������޳�DU��Qv��j��e�=}z)�����]��Ï��ޕ��m A@P~Ԫ�Cn������z�@���*L1�1@x������_���l���&P�Oi��q{P%E�!�'��ַ��G����gO�r�S{V��8������U����mlc�W�����6����Kk9Vvaq<�-d��Ű�z�م�zW�o�!��PY��X�,â+�/�sA&?�d���owa᭕̰)���¢�	L���T��,� V��z�7]:x`��?�M��j+�a�X ������������A��Nd���p�1*� �f�LY�2,��/��_�/?����/���/���������'�rp�/�Q}�P-�	�P��W����I��%U�$�2@�3bSJ���p�1	�D v ���ؗ������ Џ�ֺ�Eh6� h �Ѵ�*J�����Ge z�j�` _�ꅝ���*Tc����R[�9�3�����a�5�.,O�]���ctA�+�a���%�f� (SKZ���x�`�gx8� `Ž�ՎJ�n�W��Df�, �J��Z�6��
����̪�{�+�Ơ�M
�3���֩��U����=�+@n� ��t8�{����}E%ͧ����ny^h��������`�=��=�k�,�7~��Y$n �)�h��}b�~̌�� L(	`���'����T%���-�R�9�jjV���A�}l`/�<��8�*Y�ڥ�9}��H쬔$Q��� 2�ﶦ��YS� �Jj���f�N9�򎟁]�i�U��ļ���ڬ���dl�!(�V$Ӣ��`�_��s EbU�4)u�<�΢��E�X�4����S��eɌ�J%x%{��H&�DGE?�}�d(@Yd�H�Uѵ�TAA��[����\A�ߓn2sN�A�P5
����5�@�5�-�w<wM���x1I�ܬ�=g��8㡐=C�aÅ9F��5��U5;=W۽ܮל0����xJK�/�S��[m�f�&�?I��	�"��܃��,��GH��ឈ1r}�`�>���a���1�▄��+�2�	\z�}>�1�W*6�g\������@�➄�HU��˸��k �]�I!��ڸ�<;�4��N>_�.
8�.	j)�{Vy[v�~f�9�d�Tg�T�Ċ���[�N%J1�U$�\�A�e�%���Z��,��Fߓ�=�Dݽv��؇E���#��Q��(����HY��U&�M��Y$`����\6�К���!�ˁ�����`�n��s/3��xuk.'C�DƱ��4�
��VR1 ���!(��(9(HH�ۮv F`��� i,�6�0�v�,%?��\h}����r���F��z�ȣ'_�q�uu�jT��a�m���P�C�*���ÝGm6��D-���6����F|$ff.�  ��IDAT��u>��nTfm��!"?�f9�� �v�͵�'��sz�/��3�C��H�� ��?N��m��1=�|���T�wf����FNQ��ۮ�������/�C���;��e�# ќ��]U�B��|�{@�b�gm
���{���D~�߄��:\ό�RR��8��ꃲ�9%m��c<<ܟ�.q��Vsy����3�zsC���YK2��
�_��:[̕���1LW��öA�����_���x�D�0O�^ڢ@"�elc����?N	���mlc�?{�5�t�@5W���v�_���{����_�Z&S��G��كsY.θ��E ^x��r5��ח�aᷡ2���v7���)ACT��� G�R�$hb � �a����GX���=B<�=m�zu�:|�:|櫯���Z���Z��Qy[�����aQ� F,^7;�������Z�{��򳟽�?�w�<z� �b�"(���,|nX��{��߅�g�Vd૏X�,�k�5jI-�3� & ��b��>|��Mp��A��E5!Z� �%�؇ŧ��P�C��yM񠑚��^�	'�Y��B	U��;��?Z:�ϬF���A��4��\Ct���%!A���I��B?��@�� A������-q�L�r%�VH��>�v�Bo�1,-�70]�R#9TB�ڸV���Y?E���L[�adIi�Sn6SB �@�K�O=��Z�"V� ,��f��PB���UG�k���T��Vnnn�jaT�S5�E�N���,�I�`U�p�=T�3G@d�VPPwl�~L2��`��X��2NP����^K�h�J
V�G��%)��ٔ��Tx��%�4xXsNP}�J�u[J(�p��`9����b��׼�̳9+�Z_\\��y�L�4�xXLRD{~@(�/ ����k���f�fh�T&�̐�įe�XcfyvN��m�@(�-�v�=9��^�C?KY���	۾7�E������#�ӰtVO���g��[���g����������{͒�5���c�")�VlVo"9A��2z:{�Jz�s�f��]�6_p��� ���*��Fs��/۰_7��eVNx�~�g�0�v_�'1���"�,�y�9z:�q��rZ6��/0D:R�BO��*���ER8'.72*>�s t�o�����Ç�GO/�/u���U�I��[���Ϟ���!O�̨p���p_�K�kC̔�
��������$�o�"�'Ϩ�XY�x�r�Ӿ��v�������vס_�H��-�g�ߧR�����e�j��L�c�7�3TA$�Q�Ed��-�J���6�ia>�R{�r��\[{�
�^�l�;R��
�U�L���j =��Z�؊]A%�<���S���f�38�d�{UksgA1̳NJ���ܮ�1�8��y{����;KĘ�Uݡ�4Um�Q��s|��$R#�.h��iU�����U�J7#*��;�n�C�|��˪	�i&'��`a���%�nD'mp�Jf%9�;�S��ej�	"g����X�&�{���nͨA��G9��P���n0 ��g���H�g	�ˋk�o�𷳳{$��x���zQ���2��QT$�1W�x^ ���CҖ��<��F�u�}��"|�Z��|g���M�\s�:%m�8W�0���}ɕD1�Ix�r
��#��Xu4t�װ�9(LA0{kʲ;b�V��Hh�yd%yg�ϑ1N��/�؟��h�PuH�WKǰ��u�{�"<]�7�ʳ��0�>��^xQ^z�ey�[>gdF�MXܣ
��@����{���|���w�y�E;O..�5c.܋1'E���ܭpMzL���/*��W��Qq�PB&�j��fQԡ�C^|�%>�w�0O�X�����~���_zU��/�E�	�Q �;�]�玖����
�)�?���o��wޑ%�|¸����_���"���mlc�ؾ�m$@�6���ml_j��b�D��^�a�E��nM�ջC3+�~�'�$	����N������g���D+x��9^���.ˆ X>U�|k�Ȫ[m�I�z'Z�U�z�d�+,L�b������J�k��'�=
��9�/X��V��԰��9�� ��8���<��
�ɧ�ӟ�#?}�g��oh����� �P�l����\<筰3�h�9@�ln*�NN��i��$�-V��"��� 0������ ����Ð�ʐ���Y�b�=�h�k�5T'T�X�0��h��*�^-�P{�k�wM5���Y��DC��I1G䨊�uI��ęh��I��^��0�a 4x���M�Cx���ܪ�� ���z4T�LEf�L}��J��X}ܝ�  �*�X+��>Z~X���m�ݘ�ϧCe3^G�,S9`���9#�G����?'Ehi�i��sB�I���V-�~p�/,s"f���q�j�fTO�!�����s����xU4��
@&�m�$e���ulc�ۭ��ef�5�t�w+�X(�k5�m�'��t��_�MfJ�E��2���ֶ��Ns1�ʈ,������L2B�L-ٰC�$'�_�-ABT���KV k��nM�N�N��J���[�i�[\�V��w��=��g�1_U YkH��)�ɬ��")�!P����:c�h�vo����LԡM+�c#[9F`}Sy��V�c��(a^M�2)`��k�(����[_�vi/�^J�!㹀Z�D�XXv]3�$��]g�XB�T�P"�~�A�gĩ���X���8�$��r�|Q]No�E����A��{�d$ S��j w�`�,�wf.��y;�����4��0w#�	D�z�W�y�.2" H��[�,��+�øù��m�7�\��m6���u���~���%����>�Co���P��V3�� z���FUO��cx1ԑF�b�e�Y�F˨��d�g����w��r�3�G��va�O�u��Cޒ�Q��q�e�4� �\ �m�g�
HG����*Њ��ɳ8T)7��~l��9DT��񐡡�g�9Ym�Nf����;W�p.:�6q��z�5��~�HҰr��Z/1�&1<z>�Q��
�ː��RTVyd�iԪ���p}k��Ѡ2DN��9̒tP1�=��/r_X��:H��	�d��D�iQ�z��<��>/������W_����?
�/Z\�g4�[Q$���*6��H{-�,�m�c�BV��_ ߙj��C���´R�#H��:BĬs�J�xx�P�����B��ֶGT����O�L��έ=��#%k�*�i�/��Ch�ıa�i����P�]��p�����'O.d�ZRŋbĸ�%�mɩdU�So�3�Z..�����O�>�k�3$�95���J�s�R�$�L�;\
����5a�fڅ�5�5
C>��#����K��~�_R%�⫯��b)����=)H��ް<{#�O>����ɏ����O�b�mlc�ؾ�m$@�6���ml_B�*��@�6$�z�w��D�bd�(��*��.,����nЋ�X{��T�(#��A�;V��+��HnhCҷ�,�#z�Ǭ�D0���wJ�x@2�a_`=C�9 � �o7�v�>����#�*:`CV۫�p��>����*�R�"�*jQ��j�'��I�<8���Oa%A��Ff��t�]>��L63[%�?�)i �s�JD�X���JD�1�;i�V�*F+� *(q@ �v� Г(HA*u�Zmq��������۔�U
VǑ�U8f; �"/�!`QҺ'���OՎ�ճU!U����>bq�/��Sp���݅+;Z��e�
~�*M�~H��@7�Y|D� e�x7c�q���S�"���d�`%Ϊ:qln}ճr�7[���� �t���I>�y �3�8CS̽3m��J(�P�Ǵ�`��w,X��\ ��TRKJ�y��Z���}
������m�V���<��z� >@��9d��#ˉ0{Q@s*���cOT3�/����g$1	����y�U^�v�诜':<�n2zBK�;Pz���v)�Mit��y��b\T���P�A���ǌ
w�k�E�7�;]�{�y�p�i��v u�~��u_D�b�yΨ~+��(�#����"�*�p�X�M�R��{�m�5
��Q���T��>�!��O����b���Lf�ê
�d��*9N1�1��u{D�P�*��3��B�=�O�uB����6�obN}��a�2�u�2��3�A��UQ��A�`9g�$����[�����@�6�'�Z�����;�CEB8��tAEC ^��Ne��ю
��|��6���r*���7��at��U-� �7a�� c З�M�g�gϠv1��^��b'�<��܎��}"5�+|T�ݚْh^H��,��b�l���bI�q���8����xȃ�"� 7�LYE�jO���V��!�۩��!��EY�"��!�\�g��P3�8��d�x= [���`��L�����0�Ώ�x��v�n;埽a.������`��ܶʕ  x��s���,�!��`cs�b����=�l�b����|��_��>�1��1���w2�?����$UrU���-���z̧;>�dzo��5���!q����T^~�E޸���9h�[s�PY:O�����l�T}�p�������ԏ�s�Y�3*�:���*�����N�>�A�JC��ӊ �/�ڪU�Q�#�]䈖/K����a����s9!�=��8���%�P^%*��9g]��6g�Ǟ^<c�3>�5����w¹縧�Ws���=��Ԯ�ex^�<ԐX�9&m!��A���7��E{��vdM��(���FUE
�]����ǩ���������g�|"���������W�L�f�3@��?S�^�_y�ZbM�vh����!��6���ml_�6 c���6�/�*Da]�E�r�$i �����EFX���	·7W�=
�Ҋ',�_}�V�>��S�������'����t�,,
�v5���1U ���be�[+E��K _cѦ����9 �oo��� gevXȭ�"���'a1Zp�H��\���B�}��	��˧O���X��6:ն��s�k�p��a�
�,����pVT}ƞ���\�3�D+i+���6�A�����/McU�,U�
��63��Kf@���YԺ����m�sTrIk2��[�3��Ił�� �]��jႦ�jk��	U �?D>�*�p_z1@����c��f#�\����O��� ;�7$���JM���^��+�� �1��ᝨj@&�&&�k����l��T@:��[U��RS;'bP����N0 �F�@`����_���1o�z�l8v��D��a|�o|Q	  �����v�\��ʓC��
�+��ˏ� ����ߎ^Ū�ZC��)s�9�n�k���lAr�AG��a(�qRWJ" ����������u�}
�4��0VP���c,ࣨ�D����;3�7��ѫ�����)>�? F�RJ�k@�$�� _0�pD�-�Eā�p�Joc�p�`QX����v��w�A�bA�h�.	���gj����X��y���~�>�J�pl;�3�� ~�9l� tW���h�g� f��:1��ï�B�w;f	5��8��h�������VS�C8�j��1��v{���������x��)�e�k>,����\�~[�$	}cu������'	���^\�P)؀iFxL��yJ�i����-T:���A�X�A�Sk='F��$xzS��}�t�}���(�Q5�����$7��>���M)���-��ܯ�^skx�E�t~�Y�@[ػa�t�@f8���<U0&v��A�crWŹ��gt�-ֱ��Ƌ�M�YL���c�1pL��繢�$���ߎiWiL���C��ɓ��2˄��qrP��� �q�0WETM6T@�:g���M{�\�>�٠���<v.(��4��	%<��Ӹ�ꬮ�=!���ə����\�\�PŃk���3�����L1��W_	��4<���S��E�N����iU3��GjQ@su!/F�-���ܩS*]qD ٘Q��<���(������Nڡ�E?����������~��Z\)!���Ҁs��h��J\%C���=�B'�=��ǋ�A���V��\�6��C!��`��x/L��7�/lc2Y�{�����r��ؔ$��me��5�c��#lw�J���C0g�n�� �@�Cŉ��bn��cU��t�q���ˠz�ic�{��ٙ���[������������O��\�?�����6�����Fdlc�������b&��H�[���a�����8X3��|���YX�Z�M�s��bᎨ�`yy}-7�grzzO�u'��R<X�b�,�+z���!� �������¢xb��O����߮�sQ�<Y2���2��ۛ=��E+;������#���������sy��W��s�l�)��.B��"���Ry��~8���"@��jU�b�jc \�Y9��7:.m�5;!�� �xEk7���U�� ],��&Lp�۴���H�s��J�W
��'����i�0��s��Ix��e�f���꥞e��z�m�8Ե	׮k�T��#9*�<
͏���=���oK�0O�.�R���,'�� ��b�-��ZV�O=<V��(��:Vݣ�1|��W�z2TB���#z�2(�a{��~��f��A����@� J�VzO�	�n #j�"@�W���AR����W�������ڞ`�+��we�W#{Ŵo�mb���GZ�3%+Z_����8���ȩ@W��Z�x�k�~崮I\ӯ�$J��p��N[�����0&�	�	�:�߶ù�U����}�s2g�����e�*��p��g��YZ��<N8� �a���p�t+)=wJ �Jf��~�Z!#��`���� �/�v_ʤ��A�����U�T�@��~�t�����2u�ʏ�*�Įm�[ӆ���_=��7w����8�H���67S7�JUi�%)#����
�7��	$\�F��AE/���*��+����H�RE�=��彀6o���l��F+��7 ��⎄CD?����9@������y9Qh��蜼�������^���G^����=��>R+�Xqce���p�,Al��T����8Ƙ9��jE���<}~�6b�ֆ�����L�h �C�wc�}
������	6W2`����Oa_Af--��8���/�u8g$%��3g(�r���C3�z��m�j����B�R��Ox.`��WN��U���뛁d���]Ć��86W0��q���7'�]��j*��K�:G*)�$;ޫ����Ξ>���s^4��T&Ef�f����[a��D$TI��5�[O��7ryP�EZW٥u�1
��9�[[��3�ȕٵ��1�� ��YGO��y��Cy�W����,��'O�p<��|���-�H�#׬Ѣ�A�6�j��F�f|����.�t����b���B��mU a��~����C��X�����x����*u�[�����'J��7a鉩Ȑ��c��_fj<�P�6|S%�f#�����H	���pg��FBD?��n��؇�񂓌�M�x��*uk�AG�Gt$�G}�+��R���Z��7!qܵ� ��꽳3y󭯳����H���X桯<~��|��5��^{M^z��п&���o˟�����϶EN^��HB�6���ml_�6 c���6���e-��m���Z���dBpվ���K�v��o������YE���H+�w��"���ۥ�����1�� 4#\��Hß�\����L����Dc�Z�A��*9G�+L��6��5���<�\�
Q����3ӰX���/���|�U� ɺ]$-VeaNNO咡��`�@l:�3��������k�-��
T������Gꕺ�Yyu?�9���nn�Y�bYă��P�w6p5Kբ�Ag�W��w�r�G�|&�e��}m��A_	�j��"�mP���Pl{Yf6Q��fsp�05����
(
�;���<%��^������f 0����A��BȪ�c�Gw� ����[k�gn�䠛W/�m�@��yޗ$F��+6�� ���gnăC�F���t��I'/�v���G�#v�q���[ɦٝ�6��ڤU+ 4 �<��υWj��?�G�U���.�Ԫ�+��jy���i���z��a��L��<�]�v*2t_��ߛ"����+!�V�ĉ ���y?�Ʉ*��X�M�:C�������X,�<�P���;څ(�Y`gp}����r�����K��ʊ��B��홿��.����X� �� �Ϥ\�����dp��
�0aK�s.�}H�Ʀ*��%P��|���H�|g��7p\�)g Z-f�4N�@}P�J�I����+1m��~U�ٴ*�w[=��hg�r��$�,���9g�h����6����y�����H�>�m��ٙ���+h�擿c�l�v�k�Ef�u�u�~�+�`��#6eL�J}�ǐ�Q��kX7FT���b\2{�R2�0� fU�����M������f�YcUV9�����^	�=��a�=�w��<��vAi-6����@�?B9/!`���]��U�qku��܃LBH=�l�P�7?(ƚ���b�m(Yp�ON�)I՘Ed|d�wP������Kn+�
8��jk>��n��ھ�(�	ϡ���{؈�k�� �)~�d�׹����x�ݗ]��}������h�S�X�i��d��4��8��-����E���mY�W�$�f�]!;msKPzu�ܻw�>��֊sy�j���2���bj	K6�Ǥe���Z�5�nl~����a�ɵ+�q7�J%�ļ�v�)e����bn�|��������w�q�����w埸R��$��*ǵ��H��?7��V�>����%V;(�Tn/mB"s#�d�;��HF�Y6%!�0�jX�{�s{xI`;h�<ib�h�p����L1�f,d��o�Ϫ��,WN���e���̈DU�qL�y���K/�w���0_�m9p���r�חW�����ٟ�;��ò���}����$?�ӟ��H?�,��2���mlc�궑 ���6��}��'��̆Lr�'X�{�4�m�7%�wT_��V�.Oθ �����r[&�ݛEG��������ȗ����~#p)2��G�'���	�T j�P��r������FֻR��C,�/i�X+�Q/�P��
`T�=|(�_|�חa1���MZ0�}���`�f�Ż�H�D+�QE�Ʋ@ r����*��Ia[7DDM-�	��%�|j�p%L~�qh��g5vX��&�d�Mp�:��=�u�R%V�Cz9�h o�hŝ8��j���ؼ�3���ݫrEAV%�&�|&�c �g����%�f{������ҭ��2w���o�5�z^"SY��H'��#����c�LU���20�o�����@�nO+�Uɢ ��n5W��� ���p�T�Jr�n"c�C�)���؈��(�C�Jx}��
�E4@��T@@����X��,�=Az��Q�� Ɇ�qf�m�oZ�
�BCv1���*�8��_�]���y�vt��
ә�t�B߂}����?W�>�TYtEe>��xj���2b��P�����*V��5�>'���#7q���=3Hjf�T�P��8go�k:#h�5D�l��P,��T����߻w�k��=e�5,����&|��7��yW�;1�@�e�1X�W3�����y�����*/�O�_^՞�U���H < �����[:*�V[��H�*z�cX�0���,�A�s@���ǫ�kBZ���Mf,U�� `�v��Ǒ 1�欰��v"qJ��[��EOP�p�#����w~F0{B��Ϻ�P��^\\H��WTB��X�K)[��� t7�~�M�<��^"�[�9!�ù�;#qj��ٚ�����
�������4�x���
J���p�JAJc<'Cf��(Z#�@m* J�o�҉Eqdd�υ���k��ݐ�D��?�]2����p��l��t����� sr�	�ifA�N��vv-�ĈW�����IW~`�T��J��@��=�A����p�qTL��	-�9�_�GtJ��$#��d
�V	;9�(�L�Vo��-����M��O/�Y����c��6�6�sЧ�܆
U�p %:��.H���+Y��! �NW9	�<�
�s{s�����"�k�Ϙ�Y�;�/�kLT��iG5�No��é�VP�y�]�6�(����V�E�Nr$<����]�&6T��p;��L�w�o�[b�d�m5lK��B��kx���1�i�>4�~�|�M�i��`-XU�Bћ[�
'�����x? Ɂ�if�U�Ο�[�R��y�)9�dF"
�\���ʎƪ�ʇ"�4����J���~�c�6�O�ٮN�����Ձ�`ML�����Z>���z������o~SN�{V�'�yPo���|@�l�����\�6���ml_�6 c���6����pY�T@�p��Z�NW�E����佁j��Yoh�ȣG���씋7����CZ"�jρ����3�7ro�;��T��U�퐊�� �O?��`� m����W�pUw,���b�^���5�~�u'�U"�.��r�b_���,hʶV�ܖ� o/;Z�DU2 0�B�f�[��@�
�!ˁ����G�bd`X��k�j3l ��b6�g��p�������$�}?T�G p��^%��J�'+K���v�O߭U�Q�Z��JU�%�o�N�j��� ��=-fh����U{ �r����me�^q�� �(k��Qp�18u�:��M��kAՆ٢�Ok�4 �l�%�;>o�EVU�U�����s.�o��������Pq�]�]���$�qV[�w����yOz��� ��;�L��<��+�]!�us*�@��G�<�����oQr|�t�v<������|��X䩕��{	�"/��tV,�������Jִ��v��[G��HxTf%8� k@�Ԫ$@�4�y����I�ץ�^;�h�l���p�ED����@�ie9�9����u���J�w:%>a�ԥ��l	n�6�4̟����d�w,�9
z23d���t�,�F �Q����]3�XN���L��j�`�}/>�n�AU�kS�ߣ0��Y��"m�pu��MC}��6�]8�iù���<4ɇ�|W5P� ��2�p� �wf��Y�3N��Z=�/�����0��9>�#��?�Z߫�.�(���31�sUր.�L6�J��< ��d)7덑����q��>��j�q�٧�h��[P{����c� ���X	`��#{j2�YQ��`�@�i�N/��r�j�0n�F�4+'��c�ʥp�W���;�X�����w�O��l�K5�4o!+q_(�xh؇���.���n>~�=�#�[~N>MLœs��A��5U?���jD޷�w�-�}te���N���Jxu�~κԈ�)��V6#8Oz_̆��o��;�^����=��$|E�s��̕u~���A�A���+9��98v����}��އ�<l�"%+���"3���n/a�<��+��{�ɰD��
N�%�>?W�L�[Q��n��w}s�L���W8�1^��?g�ʧ�}"����$�>��YP��
�C����絾�8Fa��q�F఻��)�V�M�������U��h������v���?�G�|(g������9>&W������H�k��>�P�WD�,�Ӆ$a���^��>�d\�QQ�H���s��$�������
'��$A��h>�ڽ���1�$�( i��VVKͻ��A�X@��F�<o �`��{>�-xf�m��Nh���>fE�_x�'�|"Ϟ]����򗿔?x�$�Q�/�r�Փ����2�ew���?��W����?���mlc�W�����6����KhX��b~���?����=� �ez�5�w:� �����D>��S�! ��Gb������_��<���T+//���l����4�@r�
� ���ܨ����>6�Ǳ��xrs�u��Y�UɨZ<�D����PQ	`>,
b �|+Z	�67�< ��9�H�bu��� ����8�w��[�����+Y�-���{������R�UI���f�M�iD���l��)}u{����k��>M��t �&��`��#��o�C@=�*���@"�Za͍zҳ*߉�o�b���9ǁ�Աt�������svV58���`	"��q��e�&]"�H�;=���N���%Pª�\m#����W0��cע䛂*��F��Œ��ԥ���z�+0��*#���I�M����GE��k��� 
8`\W�=�����@�z 	����Z�Qנ�| �����|�ߩH�g!x�}e�����86'Kp\$'��L�CA�ְ����WU~��� �%�c�4ЮUR��Cz�ϔ Z��
���,����Ŕ �0�fa����#0U�1s�4o�
��*�q��"��bɟ�g�.�He�iM�\�f�U��c.����Ӱ_-���L0]�Y�3-�v%7�:���
�"�c�8g'�p~-ϨW2 �#CpS:��s����[9Ap!������@�<���R�0��$�V��g���a���J ڰm�mJ�[FP�yL���ga9�+��G:�Q�c㆙A �C?` 3�4&��~u���k8��<��-������9�����`#��2��(���Y�
8K.���牤;�+��� �u؞��ԃ�"n�9�+ų�S�u�;�8�h7V�q�ĝ���z�VJX��ϊ����[ߐǏ��o?���>����*+����[}�{�Ӣ��r�P��"'y*�ɚڼ�:sa�8� ��[�32W	��68��f�9�:��¸Ƶ��n��.r���O}�o@*�"��۽e�T̫��5�+�':'�MŁs���i��{Y�*�}�9����y��.s�	��,�;����n뇟��K�r�X��p%�����٠Hq�Ǜe�)FS�5��s���u����8KHTL&�j�N���qӪ�Tj1Ǟ�}��O���,�*�-G*U�9C>�Vu�oy����Uwɠz��V��7�W��@���n�\_��_�瀤�5�>�4����0�U����/ȃ�O��+>ەe#�Wײ�T|���1�ҥm�y ��x�k�n�yQ�CtV��S�@����Nm6���U8Oin�~Z��ՔgyTr �_;��`c�9
68����\��vWN�S.�q�n��ka�<~�A�O{�r���ztb���o�&�g����;����+�����3�t\ ���U�B�/�|6f����4�Yo��GFo*��p
�jx&���M�w����䣏���7h��MA���m���<��{�<�������;��T~�?�|�q��ȯ~�����K��믠X*I>���� �p���z��o���mlc�ؾ�m$@�6���ml_J�Xh�X�O���1�nP+E���+�
i����]�~�SfuLuAU�C�3�,�Pq`����y���Z*����KUX|3{�|�,���-fe1Bӕh�c��8�4U+��;���wB���±�}��aqZ�wh]��zn yu,�a!�\)�Z�E)*��$��J���>�O��j�$|F�n
��%�И�wt�ο��kp�Y�S˫E8�q�61����$s**��r�'b�����*�>?j�Uזq�pq�Em$�'��Y�PW�wְ��L����L��@�A��6OLw��Btd�4����Py|P[xf�^�vr��US�Q�8��Y���v�݁\W�W��A:W��� 2i�����!Ʒ��ͭI`<�X����C��qu��Rj��y$�ۖsB�Cs� ��w%X(v.�Oj�C*y��@C���H��;1�u�*�\��#M���JT�p�J�_|7�?��������#<;��,����ZU� �hC��xX���<�M��� 5��Q+ �}�UI¿eI�*�'V-��2�� �* 4������Lj� �KX����|��k;S",7���s�f��5�>�cc�v>���T����x��o�j����A�4�M��s�^�X�3���Noý��u<a_'Fyؼ�ϫ��� ?Ti�$Qe�tj�p �҈�F>XaU�������\D�%�}�D��e�����$v�L�U� ��>�I4� jai5�AX����Z�pb'�^42��G��U髽�:�S�ե�$���s0� �d��"mF���mQ��ca�ǣ��~L��!��N�	�gʹ׭�|�R�rp1��3���u��ܿfa�8�O�j�yl�?����1�{(����4C��^%��@L�þ��gd�|��!S��)��|:���SꎃMd?d*�2=ˆ��G��yx:����T����;�r|]}�,��sNTs�<�m�w���1��=�Y@PJ�Z.�Ł��]������م3���x��0� #����?H�i�,�����JϘ�K	՞���Rז����J�+�c\,N�Wtl�Q��gT�v$g*	3�DP6�������8ff��j�[����4 ���T��-�H�C����ck���xA�i�#�{ Y�W��\�Z>�&�����>�t!Z�a��+~W��a�$���������s��3�.|l����"�ʉ��~��,/��>�fj�k,�?���k��z���\]_���S���������"ܟ�p���Z/�c
%a}����Ï~,?���嗿�� >as�����}�wz��Ky��s٭7q6aK2��{3��|�����6��x	���mlc�?{�n*VoT~@M�
�	룎J����Ch{,�Â;*j*  �V)	��J�c�[X���c�vz~B ���+��.���v#��	N��P��ѫL��� C?�W��	����+��EdlK֔��	��7��pD
��鄋�V��ke��S@��Ζ+���n��b�q ;�l`�W 0�I>#�AK��0FU��ZHq�@��?���ތs��:�VF�e����Fl�	�5;���R�"��A	�D���eܯ��M;n�s*{�>әJ�J�<��X�VV����u��o�ѫ<��!��jh�߾�9]M�DO�� �t�w��U[�pN������z�-�7T%
�����o�5Lh��)��Z����,�Z�'�/W��w߁4'_\��D�)E\/��2�� BW���b;�V��Ȁ@|/�s�8�؁S�[J� ���\��i>>[I�/�!���j�b�K�"��v۰Ā?z�'����^c�xS'$t��_a���Eq�6X�܏�C�f��l���׎���7��NXo�ڀP���/�����Wa���G��T�A�*D�	�!�=�X-U�� �x�G�x>�P���/3��kЏwi��������/W��R�q��a�o�m���J��C��4}Փ�P�Aŕ�]j0��5�$渤��+B�LH Aeù%�H4e��v���E���.��	�����A�E��.I���g����-�j�{U�(	L`��qL�3*���6���XW��k�*�0�"�c���ɦJ�UP�\���v�{�����o�̻A��f�+���=�Ad�$���q"UxO�Ls7 I:65�'4ǧQ�C�s����ʆ,l7�tÜ@�?'�q0g� �*�	�/�`C�O��Q=s��H���߻v�	�9��sps�I.���ȼ�0N+��d�H�4�[�A���qHx6���`��vV�4���N�ɨ��| ����9:���z#|�9&�]��j>:�c9��_{L�`�:i��g{�� ��Z�P-vP�6�����ޏk%63���\yHygjז!ױ��~~�>�
>��Z:���q azvr*���r�#�|��G$m�HI�?8o8��;"x\��>\�ͮ�*
%�+�z��
3|��K�H�R��6R��ò$�<a&�q{�g���3�ڞ��p6\'��'�zC���	b)N����H���T_�Z��LԎP9��
U�~���11�Š�������6�\�`I*�q������
��I�g��ޞ7PH�[!B���w�E�q��J�r�<�\=��!���$���͞x�Tת���?z,���ߗ��[y뭯�k��&�_x(�0�u�^Y̏O�=����w��D.�<b�������_��S�v[��x&�����$<J�c��J��N>�،mlc�ؾRm$@�6���ml_j�������V!�"�UD��,͋��R@DmV"�P���rG :�,T���.��ood��5�֬(�r�����s�,��ELt��Y���G
v��. υ�lQ�5u+�ɔVPH�f�ѲJzb��z�k ��G.^[E�/^�P *1���w �v�ښ h����wT�z�%-�x���fJC��,nR����p)� K�LW,�#�PdF��62(E@o����h*zz;h�
�!L!ɉK�$6���$���I��x�;X�|�"O���Yۭ����a�����*�$2����ؙ�hM���e�c����?�1a� ���VYC �U	�gc���r ��Ӑ`��A�$�W�"��0���C�X�}A<+�-/�*�#���1��Pe�Ta �þ���-H�A�f��� 4*�r W$��(&�TCŶ�sTg��Y�:�¹ Q�g��}O���n�� B��'��u�<�䜫���j5=�+�B.,'�T=�h��LY����j ?h�d��q��G��EW0��3�,a�zA�4M"����n��=�v�eQ��ߕ2�'�sa9SA�q
�]���d��Z���V��(��D�/I�d(��.F|�x�S�6���p~zx���B?��x�:#4+���r!i��:��!�m.C��MS��}S���<'�J�)Q�ϭ��Ƶ��Zv �2ݫ%,]�����w~.'�+��UYp�D���O�N������Vn�7ry���8�4�����7عdru}+W�m�Va� \ ��!��׾XߘMsZ_Aeu�!�T����ݠ����EC�U�ZǍ���'$�1ǁI���s�q�+�� ���Bŭ�,��d��m�{�|�����������NN9;�ᄩ�՘4�~?(��g�������u���2���pe�N������סʴf ���Su�׫��@{ �ϣ����-
�{4���[�9.5b;�ͪSK�$�+�R����;��XŜG�����ԩ,l>���j�@�%e�L���"�-�a�j\}��ÇxIb=����vP�4j��,��TS�nSb{�-���+�xF����_|(/��I��	�Hx�-�	�Ԟ����;{��,�����*���m�~�w�ND��[���ȏI�$�����-5�9��)5���s��8Qh�P�*�%9�� ��4�|��Wz�%o���ůï<~z���f-�p�~��\7��x��>3�K0KԾ��V����
��Ǹ���É��.a�����~ �������~W���o�{�C�S5e#�}�X~���g��T~���d��̞��2���\<����k���N�K�D����w0���EQtx���6��}%�H��mlc�ؾ�rb5;�7��\`��vk#TOp��n��g���xƿ*诶J�{ �G��-��~�N���d���ꄡ�X�#,!ƴ��T��~m��	�O ��β1�aۺ�B�k2����f�'�u[�Ȋ��E�m���i:+-�~��@�,*G��f����ڡ(h�򓄤Ad�
v2l;Ve3< ����XV\�{���tB�j��5K#US��]��� 2D��AK+T��^��!t���/V�
�� ��KϵLY<�4J��t�ܳ�a��g��(�t��x�?�2�����ݱ�_���`�!p�����
�u>��M	�fx�C3��^"�6�[ձ�h^I�a����l�\9��@��mX��s��Ub��[�	���@���^� Ў��� T�΁>R�|��5wC�|F�VWC��V/ MUr�dP�>� Ŕ�h	���"$�U+��X	�X-g:S*��_��ھ�c��X�OD�t\3k#PRS*�b����dƪi��&��;2�Z}�&�b�-�ZD&�@`��覼�ӓS�w�$H������sȘ2�?tڶjt�c��jd%8�Z1x�>7�ݎk��waXV� ��rjX�0sb?�h`@;���&�0A��5Jn����,LW�x.�����t�LXG�����} ��/�y��P�0�B��0�g̪�Y��j�B����m ���dJ�&zL8ޮV�j:���[�5���6���&�V�e��1g1�U���d�Ԝ��񄾶XΨD\��������ES��(�"QA�8����v��pM�O�V�d$�+0��%^��ꔡ��ju���N��	�3��aĸ����`�'N$��qn[S���Wl�C!�;D$˕�l:��~7 �~������|��L����g��L#����e��o�6��Oy����;8�9���T��+9����w�h��1��G�5ձ�]�D-�\%W�(5�t'`���I�4C���D;V����ʂ�}�*ծ="{�B�y_�\ά�V��O��8�s�*ji�ұ!�}��I��w8���oԺ�W=��$q0_�1���H� c.�����j�J!��U�Ĺ�,�jfIM�+���6�Cx�1	�c�W_"I���ޒ�����=�Ǐ䣏w$�����,����������O�̨���rB��W��|�營�Ge�>$8��
��J@,�����!Ԝ6Ww͟o�4Q+ޏc�=+� J�t�g"�}J��}e��?�~��/S��l����F�;�ϖ�J��)�	�L��Y�ۘ�w��E�P ?U>3j���-�)`ㇱP�;f��n��?�W_}�*�bWʯ�{_���{�٣O�,ߴ�9r�\��!Uv�[���ʧ�qU�w���qw��(�wm��e9c���6��D	���mlcۗ��Vn��2���n���eUY��c��O�<a�[���	�ŋN�p�����X��#$A�����Jva�M�C��H�F�y	x >��W`OU�^������w���w�S[�2ޫ�4��c�"N�4�@��T �"=)e8[.���J%��@-���ͩ�@0}�Cñjٝ�6�|������D���� q>BS����i�,�u�s���o� 0I�"@[�(

�"��ϰ��>��������!Ph ���7ݱƜ}��{g�{h���4.�{�ު�᜝�k�V.�i1�s�;z��n
}��|Am���,���ŪVB��|����u�W ����s�*`����n�v >��9;^�S���bP���V�H�m3p@?�%��)ի�f��f�<bע�{f��G?t�»���n.�̮\8��z��X������8~�w��x�� Q�V�D�@Y�S9�����n]�]��in�tx�h:��ý��8�'n����j�r+T ������ ��Ad��� g�5׷�OÚ������L�� 9��V�X������0��C��C)�E�ł滰�����%R��+>�m�l��p���`o�w^&r��鳗$_4p9�jƞ�| <����bI; ;�YN,���j�Vb�H-���j�QB�| U �'�K�4�9�J��m{� q̥0���8��<fHz]+�����3£!�����Tq���X;��R�D/U��4�V��g��VAq�O�N֤���*��]��Nx=hXw��R�,�xsb22�:��N����L$j��uEs�S��i6�a�#c��8�mK��a��7F|��6e�.iq������~��
 =���H"�j/d�9����-��\/�p�<G�8���������N6U�z��?	k��rȉ����udjԦ����1X��,Oyno���lX�êGxݪ��?�����0:S��^���ܠ� ɇz�a��@l:Y�?�k������*R%S�!�ɏc5G��C&a���5��ͦ�k�"s����u����[_�ݞ����;V����X�ՂZg&�5�氟�`��qJ��-`C:S�y�ֶ��1��oe�Wȕ�a�
�?/���u���{�<W�P��r��g���>� в\�`O�@�Y�~L�`mםj������D�s����rv~ivK��׷z�*�K��fc���3`�o3����K�Wu"v��J�C�1q���er��ȭ�YIb�*�֯��)x�Ĕ%���������(xߌ�%���R�x���\G
�_3~�{!�uNW$�^�^�N��,��,H��1���A�:i��ظc2��r�'���(�V�;�O?���������%UmM�˳�W���K�>�\#,U5�{Z(5�MXë��`� ��*|݆�Y�q^�8�1�q��z��8�1�q������Td����Z<U�؃Ob
�� �͹�����l��P�(���^4sWk��2/��vt�hk]����A}*2ZI��blw| ��L�)��f/->���f������QB���(֎ӮQ�����k�� s#��	qi�^��(��\N����f�ٰ�	�������"�Ǥ�[�AU��S����B7�z`�d����Ȍ`gإ$�v���R��vIǴ���:���B1m,:�"(�B�K����>�����^��ͅ`��#���Y"��DI{��h,���'��V���_���e! �����@�D�"*h���K#|����[���.V;	�#qb �v� ��[t�z�~���YN�f���5�4�E
 +W�hy�s{L����s| �4��ZTU��þ�6U�Y����
��@�����ă�Vg��~�NS�����h�P�� v*|��DJئ�f�gmH�T�z*��]��ĺZ��˘�Pe��ӎY��%q !i�%���z/���Ȱ� vD�A�_���0�+���9(5� �_�f[�V,���r�5����n\S���҂W�z���a��A�<^��2�DA��k����C�L{�N�咠��<�q"����qn� �V��$��v�u@����eW@�b�i#��-ն�$`�1�ҿ��B�ދY!�zL�y��E
��ĀjS�)�&$�j�js�2W�6f�����+��B�Q�����o�:Oo�ny]�C @*�q�^Jj+�푅�Z�"��b��C�)����&� _���9�5��\� <�j�MY�<+�[%�z���u�p-S"0����׏A�F�8wR��3^q.P#u���ZuM�| B	�Kg$E�s_�}�<?!�CR7\��Pz���W鄊�C��!_����U�-�^^�\Q�x����4�g:XP����k����Td��W�9�뤏��z�����T ��C�8��h����Z$#���N4i(9���ש&��8>��#S����p�0_P�Tu�k���g2����i`�Nl�Mj���z�摽*�z��P���ɧ��nS���\���P�Ta��yLQ�W�i&��,�R���}�ry'�Z3b[q��D�; �y�d�Oy�� �?�nK\W�W̲��T�:��� ��hT����~��pU�P��7���L@~O���0�_��H,�<1�*��<ߦ����O�B�Gű)��D�=v�?�p�A��8l���Z^�>��Ex-�ڮ�Fµ&����5U���{��M�����Մ�
d��XH�����/���2��`�5�>[�FG]���P�&	�/�`\z���o�6�0�����������?~*��8�1���1 ��8�1�/f�;y�ʿ��u��YxX�	���O`L���;�o����<�L;6Z7�!�]��"#G�hK�d�.tY��$<�o�nLN�N�B��V5��4�� �Tx�j�R���^v��z�3� ��բg�^�9[�6$��3P6�ޤ��~*�qw'�]x�\
I���zև�|�܀!�N�SZ����$!غ���V-D�����Z��gG?m����C�%<L h�gTG���� �ƙD�aEo�6�ө����Z���BP�sn'���۱��Q��i<tFx�����
���:|�����Nʿ�s��?����Z8�[� ^?=Q�K��+�B>ĬY���E /��)�"vM�U�gx��q��Q��y�1���c��"���na�,�n]t	�|�� ��͘��_�.��L �:��[�EG��N;�x�^��^�"b��#�vm��i�]��^���#��ԁ��w�����@��Wb�d��
ۇ��z�tJ��rzq�5�`ꫛ�FP=4�j`��oI��v9}��0��;�,N,��3�HÀ=�h��Y1%Ѓ�:�4�a}��2���^A}����HB'\��ن�YW+��;�Z�:�Z@g��b�� Y���AF��H������n�n��ꥴ��ᜮ�p�\R5��W��<����Q�� �g�� b.Q����AZVS˹��c����S�P�Q�AH��
�GkU4���V�b��5�f��vE $	�9Ԇ���c̡�n��� �	C��u� 
��>֍v�G)��pLo��f��8�$(�Q7u]��-幧��iY?I��9,��F�w�rw�RRj�^H�7{��XC �D`Z	���*/8v�A��v��� Z�9ANR�T��a�a> ��}(@%��f�����e�h�D�:
��n̴G]�|!��)	���^����
��9&Y���xL��4��_��	뽩v��P\���	�CH���pB��j�L��{Mu��k��]���4��*��}�,��	a*q�dPs���]'�<+��d7rR��!����?7&�\�3��  "��ϊ����EUD��\M%���H�,��A��dRQ��XΤ� }d����a���������7�ɛ��y8�Qw/��5��}�f����,�k�K�ض':�q��k�?q}}j���T���A��$�y�P[y帧�E�Xx�7��ϲc�GG`�zX(٧��OX7N�$���E�ƕ����X7a;c�@��V�ג&���tJv�����
��T������8W[��׶{���x>O��E���;������h��4	u�
�L�˴̲��v�Q�+����S��U��ِ��!d�b^��b�����Tv��s��>�����lPl�Zg9�������AZ}�O����f���8�1�߁1 ��8�1�����s���P�j����B��&�A'��2?=�o�O��7ߑ�t��:<T�v��������䳧O�l:��fY���� ���F..0HvWmd��h/�n#j�@��V�w�2�y1�r�'q�O��Х�t���;Ic��j0��T�ݝ�CJ�iB�l>�I�Ӹ�&��B'>��6�%P����� �������F����q� G���ԀҰ]��$?�]ɇMv��J��[��N2Z"E��B�iw ��hʐϐ�
̬�V[�rrrJ@V@[ �Ui�a�c�]�
$�}^JiG#����p�`��aJ�4�&E��(!���'�Cv�SE�� �Q� �����a�L���6p��S ������ř��#0�2 �"�C9sT�C7t�׌�И�~g��(���En�*j�lo�f���*sM���D�]� � �����T����Ϧ�>��$i,@���c���K޷�g��ϐ�P֜��y�>�}�; )�y ���dT_dܷ��O���%?�����3G��4R[-��W��7K[� Y����A��g)�Q�5�.�=���2[Li�rq����f��|��"U��4H��-��� A������	���uk��x7��=A)�� ���J�՞k�9�e��m�z������`��X`���&�O�f 5�1���/����y�^�;�#��ȇ��}�]��,�e%���/��u��8��*�S�JΖs�آ�B� ��br��:�F �jR�P��*dnDB� d��d)��\6a�m¶���ԡ#� �y�_��'�6O�>�P5���^^��)�h�n�e����I"t#���K��Y%8�e��L�A@��+��p���O�RӘ9?��**v�gT}���u��1+����k=ԃ�*��yj�|z"�p|W��?������~���:����� ��Y�Zj��˽��0���3k��J��8�	�a_��c�Rbk?:X��c��N�"�DL`��R�~��p��^7[L�#�������y��^��Vc~��"�&�(<��3(� �@2�� t�#P9����*̋\-mZd'M�C��q�4����PW�a?]E�u�P�0�w��iQ+q�d?^K�LX�fÁC]�.\��[�o��n�D�;S�� p�M��J,�UekX�z������f�V�%BW<���p�r�k9�m�=j)&o�d�C�jt�Nt��뇺�,5��^#ܾ`&Y�Mh;V��V����i�L!�ɝ���F�Ƿ�-�p=��Ts-��*��'���G�H�LBm��?�/��&?�ɇa��9˺��N`ND�҉���:%�H�w�Z���d=���}D"�����4r���;����\=���J��'���l��v�#����ʱp��D�ް�I�v$"�?������Tù�=����ߺp��P��(�j���c��K6�����@*���p}��:*��(�Tn����2����{�_g�5�|�q���g���Y��`545D��O2�A�ϰF5�,�}���B�\���ek�N(8An�XO�s�Q��K��ܛ���F��y���s�qa�+�kkV��Inm������4������wG\�������8�1��l�H��c��8��\!��eD��- �$��˅���w叾�����������`��C�ݜM)'g����W������Ch�t)ә�{%���=���;V��$��d���3ڻ����Ƥ����ݗ�)�Zk��8�ʁ��w:v������,�-@8/r��jy��:��i$��f��v-��W���g6W����"�l�Ү:�7�BZ���O����wJ�@UC�.W:1�2�2("	��-�h�eky'���^oؑ �Ć�T����#��%$�<�X8he�C��ں���'��0�F�y|SZy����g�v>���UT1B�Q���x�� t����v�k�td�����ڬX (��1�^�dG����	�N&C�9�< ��� �ݳ��`~�<Uc�B��
U����%TN�j�*(/�s�7��vx_�z�}y��Exd���٠�pu�ް- 3���ok+Qе� ��4+��ܯ[�p�X@�qN�f����<W�~�,�0N��j��T��m����\NOr{[��@�}S{7����+��yOK,�[�٫�
�"������Ay�� ���?�~�:QN��jK�	 lѡ:5V���B2��"������z�L�a>���@m��&�ۦ��غ�8��+�Ւ���p�?�#S��<��ݑ��$����BO�j@8�F�v�o��B��y p���M� W��j'S����C�<��,�bſ�vPD����!��A-�Z�qZЄ���z���� �'Zs�6]�PD������Rs$`᧙:8�k��+���r�_�w�>��	h�S����:��5c>��˥U��m�y�v��ean�y݁�j�17|"����6�����o#%[�D���K�=�^@p|�s�^�cS� �oD&�@S�u�Zc:�����T=\�������#�=jh�g����q�k�K�Z�0�"�)�`�{�4a=��EX+���֎}��:����A�)����p�B=)x�`��H���y�!���uN3���!�h{H������{f��<	k���Vk����"*��]�s*A��,���v_�,}F���x_D�I��Y�b�����lZ���Yf��P�;����"ϔ�nX����;MN$5f��:�����Qe6\`%&�$��:b
U����&F�o��@�us{'W/o��x�����F����p��\�Jm�v$h&��T9��@M,�v�=�ޛ�5U��[o�-��Ux����@/q��54Ռ-֜��
 �<�*|�Hx,%#��>�UI3�~��:�{�`��F�,��]C�%�V��a�׈������Xx]�g�I%�<��������������H��ɜ����y�ד���#��j����[��z_ڙE�撩���GNRI�C؏Ĳ}x_TuFht��u�Q�(���फ~���f����D�P�Y�Z�����KU���A�5�Ab�mU�Q���c��8~�H��c��8���l�>:<v4{t�����B��� ����;oY��-���􄊏�ә�������!{t8]�
̩#�M�cWsk��Μ����1-`�2���k�3m�r��٫�� �� ����VUYZP���P�r�=��~,���\�0Lݯ�
Y�,5lz�a ����ro 
�k<n��?U�9 $�t���B�c|��{� �� ��į6)J��j��=��b�<��K���՛��z��yQdb,)��x�D"iЕ��ve8g�z��sV0�����,ҽ!h���VE�/V����}��_:tb����1i��c�`)���X�	 B�fH5�^8pO���7�� ��Ɖ6,�m��7$�t.䯐T�H�._�����)����{NJlVXJovƀ��X��\9 �nӂ��A%�d2Xt��ʱ��^�7X3uamkη8ҜfH��<��$= �)hW�qE
s���6��O�lrO$O�#]3��{�'K�Q%rwwG��h�����wr}s�]��{��PU;��T��2б��8��nEd ����-AFa��	FǍ�r���@��n+���-�͏y��ܯ�e�V�%���qT�,'��P�FC �Ѕ�*`���{��*���aϺj���)ä{#�@�F����!�;l;l�v�5�����$��T=Q�DT1�,�5�L��{�����S�(P� nc˖I$���|*�f)y�d+�)H��EP�jr�lc����	ǡܖ�Z��1I���4\*~.����g
l�O=B�P�M\k4���э��z���T����uIm�2�Q���`W��d�j,t�#S��E��� 0T� �pܙ#bK;�A&����bޗ{�I{�q"�咯Y��ẵ%���ח���c�'�Z	l(RrZl���$��I  ��9��x-(�L�F��ם�����&�����Q�%��]��B�1V��	�x%�J�0��
_'a-�R%W�굈`&ɈĈ����et\C�'�2�|�f����0A'�pN�g��@�N�ˉj �,�;�=����[9�[.��c{v�,rn��p��*��6�Ϭ"bf¾�{NBmlh��󱞨eꇒ��`�km/��zOÚ=[��5=\k�F�z��pM����h��ᵭ�������}�}j�vSɋ�/䓏>�G��I�y;���}������v�Z�{�&-�<A��(�GDɂ�X�zZ���1����=k������95�M92l"Z����᚞O�&k���|	Y^)��*D�}��Ƭ���C�!�4���NՐ��B���V�e��ύZg�2���cN? T%�V�U{$��B�޲�����,g�o-Ą*����V$3Ӹ~�_Z�N���fFU���K<�}��ą�����+����D��W�p�đ�.�.��SNC������^�E���DZXS���62���	�wF��nǜ67$z?\"c&��$����������2�q�c���#2�q�c���� �+�&ry�P�����[Oސ�|�U)���H ��D�}��r�<�'����ߓ���l�k�E|�F�ٳ�!	��F��@ұ{wO�IQ�p��O��'��l��������etց^Q��� �����{����`�K��=���C��5�cd���� �ѕ����&�U��;��QB�W;�#�,����M��:�ԫ�#@����n#$��UP�n>T���&��y>3��J��v)�>e�P��X�k�Fv��_wy�u��y�,>��]t�C�n��2 �%�)⡃U�fW��`�*b��v+����P.�
�v_w1o=�#+?z�s�,�<�>777�I��{�����{NDw6��p�����`�>���{��>��޽����� ��U�+��U��<�u���^�I�$YN`U%	�93����i��w.;!�$ !\%�����ö3���k +֗�E�Ֆ�|�YSu$<�ކ� �=�nF��>��A�%v뜤FX�unD�=���{zz��ȮҜ�q��{���I�B����+in]�z��꣒x��iz��q�&��Q/ O�jG1��|B���-��\����CmB2�UP� �����`i��CY �hP��H]$�PG�2_�yF�6�����`m i�V��<�9��$('*%�޳�F �揀�s���a��)��$5�I̬
 ʡ���d*��ګZ��C-���1�7�VL%ۮ�n�w�S�O���Gr2���/4P�0a�~��ModY�I�u�� |۞�Uyx]i��!�~�M���_�`i��VPKA�����5�"|o:��p��8� �uMuH8&���+���j�;�5�_��fu�z����assM{��fE�*MDݾ׊n���M�Q���PXiM2u:]�8c�!({�W뮆�v�=TI��$�(�g	�C�g�P����+�2�c���5O��Q>��F���Z	E���Y�I: ��o��Mz�M$���!�E5_�D�%�'御�T����"x�ae�)\����駟�6���Mr��ɐ�M����	���=k9���ۡ]��#*��5_��ؓ'o�u��g��_o���N>�8�!���n�v�RD�G\�@:6�rw�����#y���8�-�ř���;T�~����oI(zK�*�_��ϲ̈����/=��v���>�$�Ή�_>���dy&����^>{���%�X\[�6R{2��x�F)�c���y�9�"U�mV���K�ɣ��a�UJ"z��0,�-%<�Wޏ�%�[�u�4���pj��6�JxCY�u��0�y�;",~�h?�˿����s���#�E��ESK��x�	H��4`T�o�{�AP��N3�@��N�[̈WL�NL���L�*~�P�%����dPQ[V�����	ȽQ�1�q�c�[c$@�1�q�c�����?�����w��x8�}H���K>�;ZD�V!*��| ����|���{�M�o�����Wx =]��|Vȅ��������V�� ��>V�D-��a�m����7��4��W�@q} DڡI�%�k�S<U��3�}G ����څ[��f�.Cd����B`
<�c�a��I�=<h8;^�o�v���!�i�i����F�7(u_�x ?�a�%;`3�`w,�`6��.�h%��c�. b�w7
*���"�yD9ИK�̎	�E��* �t� ����)B�	���Q0@S>a*�[¾! \m��
������O����v�Z"�WG��? U�MC���6�A� ��Z	���\;I`Ms-H�$V��+*������EU�J
�`=����yײXH=@��ΣvI��
ۼCG�����W�`�'�۳���9,P��`�~�UU����2�a^��'����s`�Gg9*X�ئ�Rb$��g�|�*Ü(w{���/�y��!����(c�h�S�%�0��"�����Y��FB"�� ���v �� 	4�"a���s�f�Qo�� lv�no�k�	��~F����خ� �Nz�_"�E�����kB�vɊ����4�G���v]Uq.^_��(Yi� �Z7u�2dx��N�KQ���X���J�a8�Ɗ�?�Z���Xb���������
:�a�c�8��$|J!!��BVX�v{U��]���@a�!+ !�Q*��� �@
䙒m ��2�M���,��Av�棔-�St�Ecf�^ȼ麭�ެ�ٳ��	���^��'k%-MB{~�4��6�n�E��y�{�X�nbFXw�^��AV�S��j���{�A$'
�h�z��&Ϡ���^o2C�0T�ԭ���2c�N��q��%��C���jc�����od��?ýcfO�*���]�*���0�8�:k6IJF�1Z����/gSA;��iG<�s��F:��d��3X�a>b��_Ku�醁��`G�k2v}�+�xl�N����I�V�_]�S�Y�1"�X�v�^�H��߁`�X~�w�Km
�8�B^��մ��0G�0�(5�d� 0jh�}H����5R�l*8;=�7�~S��[,���ɓǏY���x*/^�;�ʣ7�E��GY7v�p�r��(7k��ӗ����g}VU�j�$s��ʋ�k�=(dlv�L���y�g�aP�0_�p�_��5r�6%I������˄��<l'��P�k�h[��<)���W+Q�k�
S�����*�Sd�c9�Q5�hy-��5��Y���9jjvA�h�MJ�N�=j1���vP~֘%ÜA�N���Q���ȏA5"2d�@IT�k��H��jJ;�_A��H��6]�P4?ԝZm�L��gn����Al!���E�H�Ø�n�Ҏ�텢�i�}OY���V-�H���<��1��m�vc�9��a쑝m.�c� 9��_�'��8�1���1 ��8�1�/|$3�Ve��[_����Ů>������?���ǲ�'gg�,���7d9�����L���o� ������_���׿�uWE�2���}y��~�`��z��sY*/�C�ryb`Nt���^�Oz���$<���5�н��%�Ӳ$��":�ڥ�f��=Ʌ�Y���v�67�A��A���s���S0�W[�֟��|�HЍ�Ax %�SY�jL�  �q"��uѮB���e���^)���v�B�]|MX ��ncؐ�Jt�V%�'U�$@L�G��1m"RZ��$3�7��@�; 6�����E��Ah!�A�]w��F�3~��6�ek+�W9ڑ��6I�v��`雎�V ��P����ӯ�.�z�xFGx��4yn�39A����e��� �<g�ؚʻ�}_�m���n�uL�h�q;���%�x��<鼳zr8�����n���8l��[Rr�̍ R��+J`)�W����v;���O�d8b�AS�PI �'>�9����� +�s1͕��]�w��$�kF��2_jť�4�j�+jF]��y.��*3�`�ņa� �z�c'~��O}��*l;�����{'�4��"��-�-I�����`���A��d�x�*d�p]GT���
� ��G��ݽ�"G)�U�;���Tah�¢+��~>/��>�a� $�a!am��C�W)��ToC��(��p�� vT0��,��{X'w���v�,OYc6���8'L��
9 �:�I�C�0�Faq7�y
�Y��}�����w\�v��� �'��YOY��ݞU���F����ڟL�Xo�J�����u@�y/8.a��v��7n�n���a�(���L�\��'����sv�㸔%r]&�n��o�Kn��1������̕��-WK�*���6���}ބ9|\o����TUH<x��JλW�#''�$�,��Ky����	X&�P�Tm��dP��2�5"���T9V��d�&<�r���� a�rPyԴ����|�u�����S����9���mR�R;�>��t��BE��H����k�[m��~%~�s��{�����'2+�r��\<x Iن��c3�!��$I�/(Dc���TV$ѐ}v'�¢�k�6�U�@�}�]f�<��~���pϔ��`�+�+�,*�3ԔEX-���|��3�ܢyVg�,��m�e����&��� ��p����3C�e�dnۄkS(��zǟGa]=y��>�Ռ�7��Z�Ɏ�X��2��w���9)�At2@�z�z���2����ز��T`pP������ߋ��bi�c婾_lu\�Ӆ�5��U�Uel��O-`�$8����آ���pu�!�a~���ڍ�:�W��'mQ'P�0�nc6^T�FF�RVmķ��-mNS�$y��}�:s��k-m��}QC@����>X(&����l�H�僴$_C�C'Z�^e�8�1�q��u��8�1�q������#����ExH>]��W��u��W�&>����g��?��|�{��ҿ�{_���b!�wAD$�>|$���?�g/�3tq�^ɟ|�O����������~.��g����Cr�6��2�,X�B.�1����	!D7<��Si���Ɔ5Z-��d)弢5τv.�y�Gt��Rv����V�1 ������g�tq"���:Wv�  C!�Q���P���|�䍞!�`3vt����hj5j{���<����Mx�\;]|��c� ���i��F�s��J�)d<�L�VAE��sS�?��k�=|������N�x� ���9�����������	k����K��14�E�ɪ�17x��0K'6��y6If���>�-@�lho�����ا�U)y���ǁ�m{P�hHkg�2�{T>;`�#
�)���n����l%�큥mL`?Ѩ@\d����{m-�j 
ic���~~̎ia&�Z����lĆ.g$3"��i�����J��F,enF7|��ɩf�t�����u�Zΰa^��&;�q����ig�|v/qW��I:(c֫�@x�ɪ�bÍV�e��[�s��5�-n��s�|��U���T��d�uO�����̓"�Hv;�훰�2�O� �>/��܇y�gS��(�A��R� �m�\��� �8�}�m��q��ܐhO̰k��6�t>��Z�5�k���nk��B�L�Nq���,(� &N&'����3��I�g�Ij %
�͸�D�(��GR'�'����$"R�z$��ME����d1���+3EL����9��a.l�gT;"���J���v����a]�\�+�����ULy�/)��Ѫ+|~#��qM�����v�Zs�Q�Z���T �`Q�N z1��@� ˬ�`�k�4�=�E�fKP3.�n����U`5O�6�?�=�Y���R��M��N�pa �Q��H�%l�&��R���O�1@�;��Q�6d�� F��U$ <߃�w�vY���~
5�B�Vؿ����۳	�ۆc����3�T����n[���sS��7H'�3f�DѤZ̄�Y�ߑܻ�����^��/�?���Sy��K�z���2y㭹\�?�0۹��v֏	�E4n�;��t��O�nn?'Q�k�<��\IO�Pbyt� �W=����r)󰦻0/aS���L5[���ٮ��I��bJ҄s��O��.���G��/�q�W�<���S֐�T9���������V��䘇$lkf�V��D)r����I<<zp)�����^]��Gr5$!;S*�3M�fa�j���������wJ	�	�^��#>@*� j$¢�r�*������5lT�ƹ"�`o(f�����̭6�z�p��Ц���6����޴�9B2̭*W��7�>8�δ�^��@�8�qQo�v\�� 6���0b���"KH̶��Yz���� 9T�Ŗ�zi# �)�O�	+��rkK�o�n��r��#w3��%���`����������?�8�1�q��{��8�1�q���������¿��_xK�z�]v5P�]��G�|,|��gEA�x���$�Ǐ�{���\���o�k�������Cy�𱜝��/^�ЎOXZ��3M����J�j� ���}Jx�)�4X7�W�ļ�]� #��/����c(�:]�+z��o���_S/+�����W�r/����P��M�]n�A���	�[�缘�A�\��4a�n�IL�k��N�`��hL	���ګ�`M<�k t��^��6�Rf�Djc��Nf�P�������S)���: R���{됄�&Qp���p�:T b�F�Y���&" �#p�Y���H�Ulܲ	��\��W�C6�JF���'�B�mL���^�w��%��5e��F��m@�����>����m �ܯ�㡺�8��+�>q�~' n�N�@-�čw3����T2 �.~��7��^��<X��uGko�)����r�K�-�0�����`?�^��(� 0v���1�݆���T �a��Ǔ
	S��Od@Io�5H?����	`O�xׯo�v��a�@�`����q-p�X݈�F1r5Mx���7�*v���k�����Jm���|ա,�U�����~�4	ǩ��za���}Rhw5~��\���ڑ��[>��"��ĉ�$Rc=߫�U�!
H� ���@��˘j�x��d��'k�P˹�]�d��{4����ql`�D�kr��� �D�
�D�"2��n����a���g��C@s9B�J�<`��XP��sɪ��.I�N���6���C������M$K\#�N ����q�����5푠�)���5��v���ܘ�s��w �܆����?X��j�D�8?��ֈ8�C�=��7�7$���J����k�i�I@�4��s;�Rؿe$�J?3[��Kk�Lx:�l7��v��F�k�-�M�,g���
�}ڏͧJ�º�j�x�٘M3��{�q��fr��h���6��J����˭�z��p��|is����J5X\iM��@�v���z<F$�*%A��o��{��\U��rw��Ϟ?����#������n��Vӧ2�.�z;'����$�ׄCC���JT�f�[�o�9<z�5�l�p�p>�x�y��!k��0��S]�u�4%�Ь�u����YV��\��Kxǻ�{��^Pi��-�$� +��Vb�~v-�T�`�u�9����׬�H�W2n���gO��_�җ�=�cY,fj��)��?	ks͹�vU7]�{���w��(OY<l�n ����"�=h���.�gQuPEeDCՆ���b�FB��U�$[�j[5hQ��U~���}_�Gs���ɯ���u�ab����Jɋ��k*�;�HϚ��؃k�z�ӷ	���<��E��hR�E[u����X�n��b���j��j�:�U���X!�#2�����T�p}C�T�i���Y�������(���yl��C�k3m�� �q�c��]#2�q�c���F^2�L�I1�˓7��Be����������L�\v������/�	d���9��?d��f�a�w��'r�^�����V����� ��[@z.��Z���i<�P_�q�ix�۩Ն��틎E�@x C�n����~����nv\,ih]�g7|���<x���~�!������^ؽ @E���d�ngX؜_�I�-���.Ήv>�Ax��1����Lg3ZH�S�jC�?�b?�F���49�{@�L��^��`t�Z>j� N@�R�\��a?�?���*�@O$7���2 �@�j��S[�� Hm�n���֦e�d߇�Ui���Z���y���+C��:9t;���:x�8� ����0ݞ
�P����d�lT�'��|�$��9e 3ڃu��d�]��]yf���'N�8iA�@5w��e':� ���������y'�u*g�Z� Йʓ>�@�NW#�Dt�ڃ��Y@if������Bxo��r�Ǒ�����c�?�4*���3�������������}�� �o��|H��Ё���>z��Z�vH
��@kl�}����Ǿ!'�A	�1�̑YS`����Zm`��@��>�٩���!���H��A��Y���`�vˎ��}�s�[�㽶�VN���H�@��X:�
ͺ�oo��6��K�E��O>�H�P.�� ]Lg2+�TlPw9��-;�c�:�Ib`nNB]^�8/�p��C]yu~r�@y�P�V#�$����C�x�bS� O!�i�2j��,��dXjU�|��p�,X �@�n@]�s	�f�9Px���v`Nt�`�J�c��󬙄k�D�tX6�1��`?�j-��>���_��.�$������:̕,lK��u[*��\��Y�z��v�	�*��R�W��MR��
��aN����/�,"�!�|�� 3Q�%��7���n+[�i�Җȳc@~�$�`%�,�drȐ�
�!|���D����ݯ���	G9�y1@��$0_.X�=S�A�a/'�m�������n����0�W$J����ڛZ�cTrtcVs���8ܘ£��LL�ג|�C]���ێףfa{�R�����,�ñ�����ˮ��
p�+�d��K�u�n�Z�����H���a� ���c���FA|�����������G7���v�0���z�c@I5�����l�H���:^ΣpO��m�|� Բ�h0 j��~y���"��i�<�����r%uJS������zUJ郜���� 9U�a;@ܿ��#6H�ȯ0�d��I�2��h����=��6�)�ݫ��)�l�yyss#�?�s�����B���
�}�/(����vA1��͵����D���[��g���'��`��
?�������8'�cz�NB��=`�k�[b��F2TG�8-ɽ�1�+3Yb�*���d����^e7>G�Aj	*�$��*8������\�����Gh��򹜄zZ1K�L��������r�'k^���s�pq���L#��Y��iȽ����/�H��a		�2	��h�$�uekY'E^���9RkK\kk���|vR��,4�$3^����տ�o�?�čc��8��#2�q�c����bq"��`<���*�z�W�pZ�:e�����IxЁr�x�E������� ���		���A�T|8�	n��މ?x����%���.V;}���]��0l{����N�Z�|���5��6� ��'o�3�X����	�۾��/^���b�s �MG�t�C���q��д��κ[��0�%��-��ᾳ�5�X���s�u�k3����o����:�ɓ �m`�;�ZD��#@����������M8����Qlj#H,��0�E�6�u:Z����5���K�#���x�����@&��G)�nEE�-�_�m	8<�%;�CX�[� �⠼h^��p�sȻ�=��p�CѵC��8W�8���sU��v ��R ��2�M������A6U^4���a=�cxݦQ�����ӏ����Y���$�2-�<� xv��)}�c�x��L��<�"����9LE�ڼs�D�)�"UpЂM-P�NPI����p�.f��^j�����5�4G
�=6j�3�#gօ��<K@;��6Ww���-s�$��9͖�b �]�:�� X�N�a���=۾�2�a໽\����f!���u&w�7\�X�~�ɮ5�<b&���k05��{=�L{����-|��4�Ly� ;�t�W���}8�������Vu���6{�ރҝ֗�<�5�]H>cN�^ꨉw��v���O�a���E-�|�.�g��x����Fp��(Ȣ�l��n#/�n�&�yu}G�,��\I���� �<	�wQ��d3,�,W��.�|�rߙ��w$^\݇���`�T-e�9M�J��H�\�q�׎(�mw</T6M&<�X�  x�0�`�G��9>=S+D Z}��)����P�
>ی`v~6�^ےJ_דi�u��)�9kjO� ��d=�� �%�m��p�*%r��y�EÄ�9�UE�*�6$�&l^������>��M#�W��=�r��1HQ���,�Y��{�U6�~��g�����_I�B�'����u�{�պ�Y�@BQ�Ʋu`نkTC�9�q�8��9[�F�ú�������ǵfK`n��İ]�Ӂ��&���u��&�.j��8A{�  �p��ן��q>4l Q[D%lT�Mn��.�,�h��M��u�z�W�k�3�����[W/^��͚j�b��cY�9��'�Ia]w�p��1�@�%�AJ�d�^�5�k�X�/�xW1�mNk�W�A)��;����ޭ�^%� �Y;bSÒ�	%!�Z�yWy��^Cs�q܈K�p�4����սs�iY�<�����%�ͱ&���)!;���W��"�v4�h
�����[>�*���T	�3�^jU�)��>�Twi�j-��Z
�'���q�uV�tW��M���d��8��3Fd��8��t���L����X�Q���	՞�]��;�^����毩���������w�����ݦ�֠���'�@��|�����	��}I� �fU�:�(a����>���t�@ی	 4l��]+�nÎ��>VYt�6� (�vky��)��7?� ξ�} �7x�^����ʎTB��˭iإ�e�|��Qk&<�� �����I}�l;�x�|v�)�i 4@�Y�lЅ������f������?؅�y	��6R��*�����>O�V)j­I�ݐ�X�R�� �Bgg`�+��u'�;6Kh���U�nȿo6X�W��ډ�Y���&�4N �A������k�>�t��a���w%�5�[V��/���� OC�DX��~�`���In����Ҟ��`�1���Y��1� )�W;͟�G w	'����j�]L_:^� R�(a��+|_A�H	�L{�r��v�15_ڍ@%�|�'���y��7��?�2���a���"�j��x�'(%4���{�'fes{0?�Z�@��D��xQ�5�<�=rv � ���p �
5���^��%F�.-A9��<-l�G�f�M�~��-��w��ݵU� \���C�â��z�I>?;a��~�fm�"���LNB�m "�wC@<ױ/~����'�����I��a�2ݿ|���M]�����nq����zs�ըC Xq�,����� ���i����2ppn��ú�Qo��:�H� lG�'㪆 2�a�N	U���A|�ܣ.fE&�I��lj�K���?�b(�N�?���;����zSs�hIȠr]�n�$.@�:�%�þ���c�)�J=��$�J!sr�>�x,pN�x�K�ŔjNt��y!�$	��d�����J/�y��8 @Xw��I��#�H�6�~�@-��b���4��'?_�Bd�v�@�ܔ�"����I�0g��5��&���@��e��4�H�Q	��>:짴6To���Z��zl��@�z������"?��8{/|>�k��!���v����x~�	��yG��"U3��۰�=})��s�釿�gW�pl��&�6|�l�I���Փ�k	Hy�f	�Q�?4Ulq��?E��d�
�=��C�`�V�T6a?��i�a� IM���0b���,�L����%��vC�y=�;??������*���i݃ng�i����	��&X�e��,���>\󫔤���A�w�~��l*e?P�8'�߹�B6�펇�c�?�_h�����ڍSk�9�)��J����둅w'�ݯ$�rdh6����:l��{ؖZ@:����Ѷ�u�����{�?T٪k �9*��*�:��h��1o���>���&��Y��Аa~�<�$&�6C�T�Z���d7�Z	�PSbu���_�Fg�	�{B��^��P�4礘�$�`�J��L-`ŉ��7vO����}�`�rk�
s�_����8�1�q��wg��8�1�q���r#7W/��򜝝� ��ݤ (>x$o��X~����fK��\���������s����?��?�o���X�Pcv�#'�]�t�b�6#1B Z-y �s۝��ϕ��ѧA� !�
���QhtqDV��փ���
�*�*�ر�����<<X¢�  ������˧O�ˋ�i�``<�,�ݳ;h�k6�.{����2A�X�@	̲�uF0)6(���Cyd5Ģ�m������}#�C�R���+	�>�x�u�� M��z .�X3R�g�#�Z���ǿ�����I{"�m��
�'�C<1��P��Fr��_I�q�$ �X��mo�]���8����"q�C9�{��� ̭��\q"�Xi�
|`&ȳ�d=� �"�WH�OrE��acU���៩�N�`��~��{�k=����D=��<���N8�z�7�7?UTM�%�D�k�YN�8�xlv|<0=���8b��6�4�~ }�� �
�J��Mr c^� ��	s@���kIC��� ��>ȭۘ�cdRe�_���PcS0U�.|�W N�Y�d�3>m]��v8 o��0���6
��@�:2�v�� #6-����{IV
l�����.��.ԸP#�t�%JX���+�����P������E�}��ɾp��D@s��p')
ɇ�:ũb�* ��X����cL�b�
�҆�VO�<�<�^��<4�}#Zi�)�ݛI�]פ�Z������9�Z+�T	E����2��0���)���J�>��s]�>�����7�ܭvRbn���"�m�̅� ��	b
��S��=�ޚ�q����`W\'8_J�o�G
�o�[@�8�A[�q���bɟ�Q�:�}G�~Y7jm�������ބ�p-����ś�Į+
��Xc�;#z1ܞ�sB4�E�X��"�'1�kc2���TMNn�k�4����m?��Jpt6��t֬��PC���"Ïϱ�dʬ��JN��rNI�ֶ)�w�oF�(Y���T��(0U�$vm$y[��V�xy-�������}��{��ȓa� 2-��>�#"ǙLP Q�ـQ�#jbө��J�޲���+�r�4�4T6C���s�l�êr��jYE�������F4���(�\@���u8H[��1Ud�E���$���z�v��a��6��$�z��)� �������Nܿz�2l,5���Q��kתƃ�x��ه�ו �u���m�������ěT�ڮ$�^��V�c 9ڎJ�^�5Oծ�^G[Ǝ�I��7T���܂�`��;@{Q%�jƔ����38����ڊ*P`饹T�7E.�,�8������kv��4��Rs|j��y�H�����&�:(�p]�u0���
�0e�
	V�Ϊ�--�y�*8��ߩj	g�7��9hʘ��U���_��Z)��@�����jѿ��w#ܖ|������3���c��o�	�q�c��>��o���F>��/�w�$o���}+������]^|�
�w�A�)e� di%
���v��ʭ�6$_���eyv.Qݘ�BCi���"�!�"��
���LU�Rl+���
1ex�fX��FϠ���F p��uٗ�,�C$��d���F@���	��g�����G���}y����vzI���'��p�3SIc��rvN	~��}Ϯ�~�}]k��oP��dj^�ؕ�@lt����q��D��.��h�W�Jf��H-<�L�=�%����s��Fe	��{;�Vm�[� ��8@zq�<�W~9�ÿw�;���k5X�bF����lY �� ���X� �m��c�a ȼ[~8���u�6VN9�Ȍ�����1	�`ݱ��xnե����iwr9��g�8(�k8�1C�p&�y[��Ȋ���5C�xkQRH\�DAx���[�����\�zI�އ}@�k�ر����Y��-���rp<~��=�N����߽ZIa����>b}�#E1#yA��5R"b�Af�u�bq��~�.�YX�����.�L4(.j��S�p4i���4�rV��Z�T���%���'
|a!���;?�dV>w:ےV\Uc��N�E�=.g�/3W�GG�z%w��� �
I͚*��/���m�͗<&����o��TK�ؤ��˷�ºf�:�� �8�UI `?��~�����5���yb�W��CiwvS�҄ .���-{`�a�2���vS�z�7�]gJ΢#�0�6�Q�w����v0N���!�p�@�_߭XZ@�� ��[n3�	�A��꭬�~�a;*v.7��j,��g'F
���>�h��ٚN��rL���Sju�Y�+En	H?6L�J�5��U���u���o~�����-��e�\���6r#
��P�D�W�ᣇrrz�mD�	4#U��$�
�$�"\O�� �co�4�B�����,���HH6y-þ���1f
�����w���yJ�W�vs�(�t���t�l:W���%�Z�&j��^C��=)�|r5X^�r �1���ڬI����K�*�h`�����V��6`���2̓pOs��k�N�.l�O Y�N�5���I�r��������1u��j��nMU@h�� cI��<�5 Sv�p{��Q���`�I��p��\C�v�{�G� E�uu�]�{*���RNNR|�+2	��Y����O~�u��UzO`��okyܺ�qF��c�*�yo�./rL��9Q8f�ԕ�Ϋ�X�έ�Zq0]>�`���0���Tե�v�p��M�V��V����R���y�\%h�
Z�sb������yAj!��=�q�`�U�}9�Y\0�j9���%�U
�u��e[��Sb�j|�)�N'ạ���ٜk~�-�`�:����Ҭ"����P���$԰��i�'��b��i�oR(	�>���8�1�q�֍� �8�1�q|a㽿��z���z��|�ӟ��Ǐi��X��2|}�����ݝ���������U���E���?���Ӊ�����}����3�N
�$�,���n��=DuZ�i�6��ωy5�'@Xq���3�gue8�ac�]�v�O��Rv�	;�V�Zr�J�A3I���X��ϋ)-
БƇֽ�x{��4]���o<!�s��;���C@�D�;�D�6�������BО�Y�J�,��� 4�'�8XA]��M��<�h�X��[��CGl�9@���p*P�����^�ǎvB�OI��Y)��	���	(؉��� ��D����]�t{c�N�|.1���* ��`��xP)x.�S:<"�f@q'����~���2/ �8��$ɱ���8_����^��瀣�x�<;8�?A����g�(X������� �z�,�M���2/��$&��s�'���S���K;��A��j�v�Ӊ'^T��L�W, �x�E-F�A�
�2�!���})�g�$Y?{��k�z�/G� 6�Ja�4(�b��"X��\�pN�P��v��c7tw�@}zzJ���~���W>˶�uE��Ւ]�{�������|z�4Co�� �Br�G �@T,�������������_���^�-c��_�6r�,�9��~����Ej���Ӈ�Jg����
Y���_a]��B'�1�C�&���\�MS���a�� �)l󝷹�ㄟW$�ZS��jd0�d[q�����v8���Me�.Rږ1� ���w�˂!��*���!�Z7[�h��O�P�۬���h��J�3�	ְ�a���;%�t}&��͊q�<�c֚������A�})��$_�g�s-L̞*?��`!�ض<�X#�ٌA��j�5B����EE$�>|��[��YoB�P���̨��|J]�I��8&		�����@��}������W�An3н�HT!,]%�CJ�̃ �j71e��
��^?�#u��� �O�߬���`J7�oi]j��������1�?�5�^���S=�r,4P�sX��O���\]��vm�##n��&�ٻՊ�:E��5 h��l����%�D�l��l7��0'*�h*0��*�My�.� �;�D�V����G����~��du���q��<�Z�C08��:܋]׼�:?=�"Ԋ��S)���s^L1)̫�!`�?����}� a/��蛸����Ռ�$ �g��p������y��N��^������f�ի���C�+;^�P<������r��~T��6�LE<7�nq�̉�=���Yc6XkTɖ��-;�DocQlʘ�ݏ����{,��됑�*��#���8��_6PT�B�Zd�|��z��\��I��6��-c=M;�?�{����9����W��Vw��f9 ����,��>-�N�+_���]\��~��r�mە��%
���|$���������s39YRI����p=[Ff�~�_�s�I����c��8~��H��c��8�������Z�ljn�����ٳ�K��?�&;�NOO䍷ޔ��y[�_>�ۛ;P� ����]��՝��?�5��f-_��oȓ'O���1�� N�v	�Kv��@��C7 �8U�~h2�C)�} ��A	��4x(�0S�6�чSx��߲[�@Óoۣ����״(A.�|J�o|㛴��nv��-5*n3��̬���D���HG��0�kכ]������2 	��=b}�MLI�|�Y��o]�@_����jZ5�c��}�Ɣ����qX�u�Kb��q�64�ߙ�oq�k�~�Zx�.Wۘ����R ���?��9a�~M��ތ�];��@�NZ+*��*2b�`����{���
���\Vr�3k6�� � &��!�DV���0�DF<d�t�4�g _�=lo�<���j��e� Xo��0�E������\��`U�2`+�y�n�n�f��^р�H��q,�x�TI�L�<5��lՎ:�#v'��c�y�t	��?��W�����][�sM=Fj�4W�>�D[��̞ż�u��jE�m
;��� �ں����C[��\m�t��zt�3p=�L�,3k�p~׍Z8�Fj��Z�<iuV����ڤ�I��� ��U�����O��JI���0���sK��O?�YV�2Թ��%�)���k�, �k��NIC� k)X�ML��� 
 �+,'3�ےs	8��4�H�a�a���`�G�*0���:Uu`�2$IY��:��c��^AZK�Ѩ�UI��� q�^d��&X
��@�����2\�'����ܯW���S�!fń�X��J	��5��4fӥ������bZ�d��w%Li�;�-�D�����0V@:�W���/�u�Z��[;��I6�b����N�Z���,I�0CG�;,!($@���b.c>n6{�}(�B	�L���^�I���>�`�b��+/�!���׃��#1�iPм|�Rn�Vl
�WiV}8��h�� p�y�B]Q��A�v k�_�޴I�����枵W��w��	`��DbD��Uf���(3���(�D�i3C�h���^��+��XuϹ����"?c��F��UefDx�_��sv����g ��"�4�VM�q1��w�r[Y�Al�z�4A1yQ�1��=|v�3��5�������7<} t~~!�[��;���E���Q��:E���60�F�b�f8e�J��'`Wd�������������*�BΫ����~L���K�W���5x��+SƦ3/�����4i�����A�K����W�p�X�8�C�L�����Cɺ44���k��9_��O�<��'��O?�R?�K����g$ᣌ�/0�.kcL�
fg��h�P�'[�e��U����0����	s!��"���^=�X��� >̊�A�1^�e�uŀ+(1��w�O��y;�j�y�̖����F��1�9ꊅ6���GĒs�"���fX!r`U��Cz�.:�7�@d�0P!�O�e���9��KY�k>/p��9�,�R�;�{�=�˿�>�����/)?����~65�¤��(��y��~���X?�6���M���T����h�ޗ��k]~k]P�������������W�ꥴ�mmk[۾��@�ֶ���m��Χ҉Ǎ?r7�)�죏���+�?59�(h���a��o�Lut�|{?�M�DF�|ͫ�sn��%F|?M$9<��n��n��4��4N��п*.���庛�Nܰv�7�H��gE�����`K�-��;�02�������%M׳����F�Ȗa3�G鯛�^������W�</$�RV�!�p�J#�"0���Ǒ�P�������c��J�(���]*V"�	Y��7`R-�t�5[�Y�䆖D+j�`�\��4|�c�����`�D4�/�܇�P	����?��d�i��C���4Ƶ�*7�n{�����TH�.��_C9���
��&y�}�#W!�D�8�\
��]��wvo�w p��A���|V_�e#o�Y"��=#���t[��$���7$���
��Qv=8�l�$�"YL7����zP���tXml���T`�A��^�XH�`|BF�	_Q�5e7��,^[���"=|��73�xpq  ����9nh����3r"��`ɜB⽮<~�#��t]�M,쫌Je$H��zܤ"Ѐd���7��7y4��3V��|���Z�R�U`�yB ����q��dMa����aW�����,�Ϣx��X(+_y�����{f"�L�������U>'��;=�D>r��Խ�����P�O���I�$��F}�4�A����P������lBv@�E�}�>�.P\A 2�  epE�:홤� f��gu?��k�n��٨��f� K����D��1����p�� H��}<���UӺ� v�R�R�H;����q�7s��pY�������tĹ]i����ϵ/f2i�._�kSxdLl\�A�H� �Дc$\�T�[.6duzɸP�rV����2�:�Fb�9 ?BD6_�7��3n������C�������q׋8 -��$xru}��&�h���dN��� *K$n�О����t$���1�[TV��N���.��(t-�k_F����몑��@1�|g)	�L�{��N�ʃv>V!�x�gm%��h�[qE��G>^,����ww��$5�rL�FEO�;�^��b�l��l���� ѿ��8O�^SH�GBfƆ�A�WS�ح�� �N�ƣ%�p<$�1�觎
{y�`���o�ڄ1�q�?(i\QD��FUa2M�g
��9=;sd}K�/����r��c���

��0�:���a}oVъs�]��L�F�ǣ��x�@�J���N�r?�g��z9S2s!�0��5��*i@��j/sJ_Cؤ� m��B��!�G!�b��3�w�����)m,�D H�x�< `�K��d��ˌRW��!��0*��q�b ���<�^
��
L�{ӁZp��2�!�5�h��'�������L2���R��6���H��@~��+YD��ݻt�����<tV��Ɣh|�7�?�����[|�?8�����j��&�l�y8��$!���g���?��?�?�˿��(�֫G����3�܌�N��e���=!�mmk[���-m- Ҷ���mm���_��_�E2�!�0��o�Z0�^N�g�S�������=9<<�~�k�կ~ɤ��t���gڏ(u{;��ۗ�xO�'���{�:d3�����	����_��%�r��\N��u�ؓ2��w0G �`_���N�%��Ύ�!��� Q7�+=���8�ސ�P0B ���Ԗ�/3�g��|T���q����R._�ss����9�<fG_^31�&7Ŗ`�t���36��~���3jE��dax��b�� �pƫ��[�̏�O��Y.h h���h�#ፄ1�-QmI��$��w$󓘲5Y����� LX��M5t���\�ti���� ��K��ǓJ�$SJ�7�Hr�z�П1E﬜��*�����Q8�z#�mMmY�n��+m�Q�~Oih��5�����R�N �M��Ž���
H3�<�
9:�>�dH����=�%X�D�7���nBγI����`���I��m�E�{�5��}�d��rl$.:u�R ���H`lD�B�[6�b����=BB�[��VZ%L�p@5/+X����l��s@��WM��ݳ� "��˅l�Hw�G$����U�1w����!�d2&d'1V	�I�,]"�K�X"<ZeL���s9;=�?������7��j(K������DL�X:1���bm`<f�@�F\��`@`^q3N�&S)���`���LQǪܧL�%�IǠ��އL��:�������3$�K�(t������́x���dXd�:]{�,�:�BY-2훹o�z>z�?����Z��;}o����T����QRprw��l�x�1��XH��2�9�g�J�������8 `�/'U����Mß@X|C��^]�b>�nb� $�?��=V3�B�/���~r�5��P��D|p������
0=p?�㑄�H�����1k��;�~� �\�u�cj]��iF?�^�q��)M}��\^|y#�ne	m}��|C�s�9 �*��+V�5�?M{d��Ԣ�mX:):H٘�KVe�!�S�N�Ϟ�&&;�L�g�
�M�gS���*&Q�߅4UГ���%:������0qg{	k�U��l�b������v�Q�U��Zr�8`4������?��%e� ���۸+t-����x�G�d�%$�G��3
�}�i�NP4���䪲l�w"�-0",A�&�`�<��[��*d����L�k�A�X��Z������"2�	y��센0�r�w�~��*$�q���כ��ޛ���5�ǎ!�`���oY�"vl���|��;k���8�
˰.w�C�P���k�
�B/t���=�E����H֫�h1[������rC9��c�^_]�����Nf�XQ�,��s�X|�a]\�h8`1>ci3z�ٱA:P�L��́��Q����c ��+��Ln�dm��q��{���+Ƽ0 ��W�20���b.�`W�Q�}+cg0��.x�x4�5`�Y#�ilR���I?{Q�ɐ���	M.
�^�~J�D�X��ٞ��Vs獓���H]��R�������|�P��@��^��t$G���(R��Â}��ե�2�p�����&�V���L6K���rlW�_N(����|�}Y��)��V	}F�uC�o<}C�NN�?K���'��/8��utws�u �����/^<�/����?����~�C9}t&�Η��5��Wu�כ4�5��u+�ն���m��� mk[��ֶ?j˲97����U	��}�������?�Q��͕�^�ҍk$�ߐ�7ީIT�,$=����/�$���9+�>��Sn�����y%=��N��I����X�rË��frh&�H��xmo0���}��y}l�t�#v����BB��Yi����������|63#TT�NQ�w΄�|p�mtɈ���|�X����ӄB	(Td"����S�� �4@����8��%��Lil��%%�L��ǬH���PN>H��(�R7VE�cR�0��
d4��6�v�<�����UD�څU��>Ԯ�RY��(׍d.kY���f�_���VJ7B5���k��w ���U�V�I�x�������S4�d)N��ʺ!K��d'�V%�n��M��t��w|��z/�=�yu��<*�=��,]�%���eܰE<��7��e�f��� ���0�7 �� ��4$Hs�n��ya��H@A�>u�Y����z�a����W[�W%C�����{�> �h�T��Mb�� yp�w�{K~��_�6��}����I-����00U��f��6��@�xn�>'mGO��d���o�V��Ř����� ��혜dz4��b���X�F���1��7�Ro��Q���3 �� @Ta���{��9�8����)���D��&�9M)Å����{Jo9�#�.`�wQ��-d���q�e�?&�U;�_��l<W'M���sجA����]3�f~Y�C�O~VL�e�?	�$��[$S%��0���0@.x�����r�编�|�����!=>P�k&�Rl��te���>�./����Wr{3ј��f��y9t�Pa��;ߥ����#)�7g��X����\7�y�A�t�$cw<dQ =>�;��:		" >a�4C�녗�Tbn�%fkǱ�;��[:c^d=�; ki��? ���
x
(�=��p�r��ư*k�%Um�8G��ڇX�6�ȡ�Rd�1��z�*�}G�>������c&�Fc?X����'�G�bf��@$�=c��y�ƣ�S�иJ|�z�J_&&�k��(�;HP���z����xw��@"�p�ɍɓ���on��N�a?c�}(0�dH��a"���׬+�P,l����8$1KHI��c��M	���1�rU�}��"楱Ʉ��ŲL�Ε�	�nw΂�9���Ūar �Az@ GΕ�0/5�bL%c{��I$a����QXL���Xu��5jl�h߾������P��,���s^\�җ�&���3
<x�	eCs9�k,X��<n��l�Ʈ0�����v�ϭy+ �}��g�Oۿg��� @J�c2�|�Y�2� ����3�n4���P���ɱ��������p��<������-�20m0w<Kc���F��~}.��l=�Nt(	2�.!U���\�o�o����3������˗�Y�^�R��\�G�����!ƀuy�����I��6|�D< p��w&�ruuŢ�'O��ó3��C��y���'oG��N��Y$�ۼX��ֶ�}�[��ֶ���m����G�� �eF��d��O?�X7H]��Ԕ�:>ܓ!���zh.I�-�%~V���w����~,��_2��d�YbӮ;�Ɛ��I��A�_7��D�NW�Tl�ưS�<��&�K��?��@h0k����L��N�@FȪo��x���|~�@n�od	ً�s��x%�^]JԉX9�mJ�8��p�X�s"N�$ߘ�5��Y�duI-3^��&��ܭ�o�fL�II��:	RT��sHv	��,7=k���L- �&ɪ�2U�e��?n����u��r��Ѣ i*�Q�����Íԩ3H�䖙��`�N�����n�ewL=i��_����p�[U��kF�'}E)��}@.�L�C$lM�!ObU�&���d���{�LA�5ܺ �2HXUL@f�}ͤa��L�[�,</���s39�������q�@%�೐��c�l�8s_w]�����7���AR�����8�/�*��z�l���>cB-I,�6];��j� T���{�c�ǁ�㯝̗�����S��N%���ۅ�#�n	xD��� u�d& �H]tx'T�Xa�%�_0&c��e��J��i�$Aʾ68*�e�X��|*�q�H������ʀR~vѸ�o���ig�3I�HSuL����� Y�.J!��Z��_�O j.�n�ُs��2frs}�1� ���o�; 1�T���T��N$_-%�ς�8@�IP���Z�䷐|�i�U��L�ͦ3V�ӑt�V1W�[�d�v?Ē� C�4d���-$I�7�] ��@�m��s�X�Z�b6_���L��P�pf�:��L�
����g��\����^'��&����a�_?��i��Q�D��f��*�Zi?w����{C_�������������H�b^��hs!�s4�n �IRl�7���� P�[)>�N�V�i�
y/A�cҍ��c�KbS��V���5rGH����^���=w~-��w��	�w:����C	N��k��a�G����\}l΋���ԁH��݃%��Uހ�1�vb�_��]Y�蕭��Q`q�K6ր�`L�1�ct]4��<fQ�'��0��ւUC��hL��Җ�ʝ9��~K�,WS~�ymeO��c9>9$��7.᱓;m��d%
2ƃ���19���s��mrs#{�\D丵+qIxT����C�c'�3�B��H�cR�sCC 	�_�R���~Q���%�ôC #�,V̦W"WBY���çϞ�ٓ��P�����s���y�о��@~ȁ�i�g��t��B��9���ٳ;ԣ�v�zb,�$�g��7���"6˼ܡ��46o��c�HakL�X�+��~xև���~*�Á<<}��Ӈrvr"GǇ|����X ������ϴ�N� HI��ø�gr�|{������?���^.���Ջ��V���~"��Fn�3_�g�=��xo_��`t���P��T�}g7�<ހ��h��v�s���,��N��vNz�?2� �����G����#��1�у�a���*��q��Ө��"��a�
���mmk[۾��@�ֶ���mԆ����O��Z"V�-u�钪�d��KU&�� �G�w٬tU�%j0j����m}�����}�yu�LZ`zG���|�$�-:��-�ߙn�Uc�@�������Q��x�?�,�$	걙?#�Z�ܘ�8���{$ӆñ<8{�?����V>����o~%���e>������/�3Q%�A��Í��յ�M��'a��D�1�����*3���%��!�*��i.*� �B]pn�SJ�n�WV�m�����IqSqo�Ֆ�	�Ua�7��L��,_��G�{��L��L��(���fml�[��S�����K�'����Z���7H�J�rX�����`	���x@U���u�?'��<��U�&���̜�@
 >Y�7^����h�����O�{���E�}@؏.!G&E�����"��Sɐ(���,(yS;0���
$�|M����������Fr�W\�/c����((;��wׁ���Ii�Lf��A7��>@�ǉ���I�!q7�\'[�+O�>�gO����o����n�3�ㅬ�4�$�Я�X_K?�Պ��.d��+h���|�6�����&��gNM�Oҳ
d���3����ŖHP�4a�����f�](��	ux~4s�ѢB&�@�Z�UO�z�d��t�������VN����t��e��I{��4���>. ���XQ�iy?��"5�	*�3�p~N�1��4��_?g��IE橣��*�@t�P�����������D,�;0��� ��;��C�L���IV	�T@�@��r9%���8�Ȕ�ϖ2��(����� eȝ�;Ҿ4~��G�J��o�Z�jo���sd�[W��K@Cjo>�D�g�}dE�����������q�1~�G)IH�m�y��ёqf��fI��� �m>E�'�ެ�Mb�.{�3��~��=q�w����}9��l&���L�����0�i],�}'�tUF������C��{ c$r �L�ib�n�2�_ެ	�=�&\Ǳ�cL�X>�2�]��:V�/�gf�&g�i>�f^ϓN����z���bF����>YA(^�K�J�#k�U�*��X[jF�n! U�ڙ�b9>>���3�G�w�.�+�$\�*����pO�<z*o={K��?�>B�y}�����`<|L�%�!�G�������%`��W� p�obNd��^�`V9�H ! H!���
��Xz��d��߆��������fS�ÚE8��3|$2��Q9eQ#g,^������X��yS�������(F�� ��b��8�'�bD���sL��`$J<3��	j�B�+��'���4�<�w���ϵ_�?b�j�b�%�9��l� |��ױ~�U�{�=�������w�ɇȗ_|AF��o�9u��|=��}Jy����I$㽑>�O����� v�����w�Jzn�z�d}��)yM?N����l1�lbLU�\�b	�ƷϡA�N���mmk[����n- Ҷ���mm�����@��D�A�t4���Q44�#��@�ޠ�P;:�q&z%��;RKW�Jv�cؠ�򶜭)�������drO)l&��>��z<$�аQ*ʭi46H$a
�:ҍ�Çt�w�$6�H,��&2B�aZe�OL�
P�?L�$m6�H���uY�z��!|I�cy��g��G�իW����F�d��@����;�����t�i૛?�B�5X-�R,]�Xe6�}��׍���L�t��骧��]��s��E��4�EE���C�y>0Ix�΀Iޘ�d�cj��s@ѕ�I-$@��HT�=@����#��ˤ���'-�K4����0U �,���U#)� ��BЮa�N��2Tf�IOjIc����Yi:�E�X�K��iu��ڙ��zc���	�<2�I3�.�,�w '�^0�C���W�����ʒ����D�k`	YX��[w�ǵ
^�%���嘘<��2XL�8��L<���dv+K4{���� �x����
��!��&�R7 P��eSqkU�H�0W�+�pl�y{�~# FKP�������G�H~�O�z:�^ړ �0��?�q��������:�B���E�����u\�zir,NU݈]e�1�пĒ�Θ�10d〓�hL�+�|�zu��je�,ʟ�η�bUԋWB7�|"����cȧ�)!�)��g�93��Ě䒈I��l�*��7�[��Od>_��` #��H�-fs�%+�����$�jv\?��Ȟ�*�}��Q���|%��}:��(Z��>��͈g`�
��bO]�|��K<!y�%� ��L~Z�4��P�ץ_�� {a���f�dH�LV��.-���2�M��0�#î���q ���s�5N�����c���e��؄l����(`�v:}&Z����9�nCb���M3i�>�IT�q [6�s�� 9 ����x�X���]��|�䗙AG�w)�3'����e#��Z��&v��R�<�!1d���87R%\�pn�H��LU�o��3>^��6?	Y&�V�f��,s��:��<n|u�q�tzo�Q��'P���3���'P��:���S�����^kWФ&m�se&�8i.���L��=�5�U(���>��_ϗo�g':i2�\!ɅxB�NTck�-�Ϟ>��a~бXq\��C}�Zq���������Ť�`,O��}6Z���!|t��/^��9p��i%3����`�B���`&wfl��0�/(�hk5��j2@"�D�P��
�]�j8���6�h܋�Ap�cm�>�A�(�����R��9���G���|���7��ʺZ�*��犅!'1��� �ғ9B������f�)\�i�%bl�GM��k�MIF�8挍;�`�<�ԣ}~Š�Q��}�Ѐ�����3�ƙG�˛�ޔ��C>�;�f e��Y�� q�1�y�n��Z�(0�Xl�)�צ�Z�����{�ʓ����|._|����2ƮWK�Mʮ&��^�1�+O>�.�Ͽ��D�=tn�!\ӓ�(l(LJc��g]mra��Xo0�0�:�cYV�:��eDQ賐�?��}%<��4�^�]mk[��ֶo]k����mmk�����u���<
��rK��DU� QQ��Bl�*nW"n!ǀ$�P��X��]K.��zV���r�`�2�It��xJ���(J0�L��us�'<���S�I ��M`��:�7�mr�K�J.�Lj�9����5�GH��z�AR���ߢ���;ﰂ�o�ÿ��/e�\Q_����f�O�xKN�x��tfէNR� D�$�y�$���be:��}�U�TX	����<L��/���k�[3Q�dA��į'ˍ���S�=�%�*K��b|0PW���aE�����d&���dmp������V�K���Y��v���Ʈp��a/T���d�DC�q�$[Y�f[?�;ez2Kݘ�j��
`�_�{�4�ÿ�{���`��C������>~�*��ǂ�G����D��ah|5�g�pBy$���c���rU��&q���]VG�8FɖD�$E}��Ʊ���y\Jиjj�S��7�K|�ٱ�F��T���}ļF�-��ƯM.�n��ߖk��%͜7br��J�c�2����E2���?��)mV9�7J�Ս/ �3�`�!!fX�rssä�xԕ9 x�¤7����� ��� Ihʐ?�Q9�q�ǽ��iD�	X��[�����6?И��� $<��}��9���}]@�f�N�n�c�De&���L^�@Hfտ3Bg�Soҁ]�mV "E����uc�VH�#����XQ:�#Tk����2���~�h��/f�B-������G�w�y��Jz�l�W�І��F\�+;�`����"�����؅!3G�&���y~�.5U��|�wE������U����͔}��~A�;>f� �V^h�C�Z����c
����@ ���1��>�(��I�a,YL��K�$�[L`v����$&$��۲�7����sLb.c}����x��cd`@4@,c��\�����C1�/�q#h<��_)uq$�2K;�},½�1ټA�1}Ai'���:}��څX��p��7V@�1u����(JR�-H�bY�Z�7��L�u��x��+K'M����J��5c�Bl0�J�����c�u�0��!�2��Lu�G,LI�d�v�����ى��o��\\_���dA�Qz�X�$,��F�(���=;�#�����F. ���-��i��e�Z �#Jw�P���W�1�g'����Ij���3_,d0�t ��Al���}m�bi�
�s�����9�q$�h4�36����AT���/i~��w�z�r���q�R��}�/N�o�A��)V��ɤ0�J2y5άKNY��W6�P8�8�XG��z�6F+��!�g�G��ʳg���Ç���2����K��,�e���s.|�?x*�=!�j���\��eC��눿%~%2�/)��׽6�'���e6�2�`ͅ�:��h �N]k�s���ۨ��UW�#*� i[��ֶoyk����mmk�����WL���n�����}Y�sK��p�K\Ǳ�0`dBE��D�T6�؄UA�S�E3T	�|KV�k���&ܸF.�
�$JY��$t�X�Fq8�!� G��Vk�%�;��n�{La���*��P��tH�����z��Z7��)Mw��F�����)	@��P������z�R7��y?���׾��w����zM�����Z��\�#��5�+cg��D�D�
�H�T��{������֨�m�1�#�!:p�Nl�-1��07_�V�f�IMrl6�Դ���C|R۪]�=�tb �%J�{��>�e�f �y�[�l������&��9����%�+o��%���u�u���� �*F$t��������,���jB��K�Pz	oV����a�s$��W�%E+&��0 � ��y�׉c���nE��Ӑ�r����g���c�TO�c�'&����H{�.��!#��L&U�KXU�b7w`N����ѱ��q�Y8щ���=pC)��DH���� ��B8��4��){m�+��<�c�TA0�2 81�on�e�Z��3�+�1����2&���T�߉��vRg%�&�O��<Uv��R8����g��J(�� �AF������=}�ca� �i� Č+�t�!x���Xs�����.�X@	L����ҁ����ı�r{YT����z�H�����ZP+[<x {�1���qڀy��*3Jҭ;	��m-�)`�`u}�T�{O�F
�z l]��;_J�j�1uP��@��(zWϵB���`rl��/�`����B��jCVF�q� UN����a�\�E�XҞ%�,|c�3�	^�Nf2�O5�g�f��!�6�d"���ql�N*�rC�=�͢	�;��Q`�~�u(5&x�CJL&w�s$�|�qmXT���1b]0Q�#c�)�q���xC�ʝo�{�[9/����]g`��Kb�o�Y����$�}s�u	d)����n��΃��Pc�T��ƢhbW�Ѓ!^�ϳ:bpo7N&������ak��M���Ӂ���d:Ud�yƃ��"�y"y0��Y��������蘷H`�-�cU��P}s+�F�/x�	�����n�btet�J�["&�L���L��Fzqoo��`aF.�"���,��7��8���sp��=��K'����y�v�X����l�wũ��K�R�'a�����=3�eX�K�e��Xզ0�%�C �J��s��C&�<�=�[A�-�3�u�Ɓ�c��ċ	j�ra�0)Q�ǃ����Wi\bL�ЭQ\���ʤ������ �*����5]� Zq��Ƣ�zz���|]�{��o�O�Ǉc��'d3��*��N*�OK���RW�Z���l׽qK�3d��Y�"�쥄�~O��iҗU�g'�-���3�|8(	ۍ�?H��c=�B�����W�k>;PZn��=���r�����ߚ�����^ `�������%2�rt,�g�r����^"��Kom��&��@XҶ���mm�V� i[��ֶ����m���_�]BLL׳%7�����a��l{��%���v��(�_���%����%RǕndǺJW?��|n�IJS�Jr'	��J7�ibCn<}u:4��������,���*\�(��a�	(b2f�f�S$�����	�(��ݭ�sʻ,i�Z�ho,�ǧ��~�����k�ruu�$��&S��?���r
��Ԓ~L�"�_�HVl\b���[vHY��2�db�)�LTlCB���0jd,�oL3�YA�f?���[&L� Y%%�QAJࢢdG�*l��+Ɵ����*�@��v��IڳDT�K�Fb�`�gZҗ{��ۛ��4��>,��RKY�u��]#t�W����He��d��4~���g��24��%�ܤ�����8��<��,Ǽ�&ҞI��_�կ��k_����5 �Vf�]5�8	\�n��}-Q ��v��-�����u�NS��;kP,��!���MR�E<�)<c�'z���Fr�y�x�$��|�3����I8餢�v�Rx�I꫼ᙐ����t��0%Q��%'p�6�~�H̶Q��䖀��P����y92w=E�:��L���.tN�}���
���ݝ�󂉰������ԉ	�/�vz�A�O���<㜧̚gPG��.�x��\�xG�� .#�[����9�@	_V��8N��ȥT:�ד����sE��j߳�������sJ�g�YJ�GL�j #S��I�-�@WIy�����2Ѧ�.��1�I2�N��b:���@&=����T��:ֳʪȵ�7���K�X6�(K&�T]z-3�C%� O��F\Y����s�s�H�z�7��N9.��υ�/���S���@:��+�/�H�eS��~N��8uh0�?��ıͣ��4�Maǀ�@` !$�6�y,���V�*�C������(�VT�ym��D�wJ����]?J��Ebl�pe�c�77ײб�k����ºpIn����m`[�x$��{d�Oм�����Ƴ>�{g�v�l4[_,�.����\y���jJ��8���Yx&��R���\��(���N`��j����������e�J`���,0���͐�t�ta��}0����V]J����������B"�)w�3�O՜��`[-�(�c��o����{���n2!����*��<`g��I;VR� #�h�J���XPa�8k�n�7Ày���X�g����PfK�7z̥������ 	s��alv���@8_9&��9[)Hϔ�[m,���U��k7o���t6׋F򮬍�j���y��Xq)�8|%�i���((�k0��l���[o�%��6�`l���l)� �``��Ӿd�?{��M0��Σ/_�\O���l��i�c�����1�0�=�����|�Ͽ�x��ͺ>����d��G %�{���y}"��83�����lB�e�X������_�;�䓏�V�Ōg��{:�ƃ��t�B�������y�ɣGrvr*�QWc��>Dُ��ϗ���:��UY�����mmk۷�� H��ֶ����NOeruNCCV�%�����T�ǆ�;X��;ݥ� c�d�n~3T>2i����{ݠcӊ�<̳��.��^<.�w?��L��QCZj�* ��_ld�Y�F}��'�����b��3��qZԑU��_ _�T�Cra��s���	��k��\3I��[-(%R�4�q�L������������%�9��_�=�I40A~���x^ؔ������VW#sn��i&��΄��A��uc�-#�)���x�$����M����A#��W!=[h�Z��36������~H4�}�3��D0*���&_@Y����{ ��D1u�i7��Bj	i&��7R�2i����UfU��r�/Ka@�7�FŦ5���)&�j��0ȣ��N�1P�Tz����'5��a`,n�͸�*�qoG����;V#��욙N�J����4rU8Oxj�����݅I;Օ���v�ȶ�O��A���<p�H��NoÒ}������\ x��!ȣ0j�I��gNy#`��A�Ӓ�r1L0��}�4LH�4�1�7�l����֛�#y��w���>�	���v㫣� *��ǃ��8`/\^�1)	Y�R�5��JzD���4��rY��^�Ų˅�:��N����+v��r�0���
t�S�Js�ҖYI ���{{O�2c���w�4 ����8�F�y�a A:�!9���p~Ȃd�9��q�B�Lt<�hXd&�L��"��� �Ȥ���^ӝ����Jj=����y��:�
��7�%%���L�,�H懌��%�c9[h��]��Ž�Ɓa1Hd�5aa]�� �`	���y��s ��t�a�w ϜZ��`�3)(y��̸f?���Q��HA�L�X� g�����>CN�En�8 ��lNv�� ���\c��q`c�
sg�ە�[&�;⭸k�'A��b�v	mcEDNf�`<X��zuu�0����`��U¤.���nNF��Nª�{"*�G�	j�f��:���_�0� *g�B,���P����Wk!������������@�C�&�=�th����́�n�������e=�F�����8�A�u������:�mƕ,��yƈ8fY�@hĳ��k=����\�ƱB�a�g�0ټz�K��>�5������IKT��gF���7 >᝗&�ј`���Ї�bb��7���Z�P��pr��FמM�{3YN(G���1=�z��)���\VǮ�	�2�s�����Wsy�q`4���6�kx��gr��;�1�^��1�_� "���~��v�O����l(&���/>�,���Xm�aN&]EP�	�+��:�2	���`ONNN$��^"�K��K�4AN���k��M(�PLt���!+��">c���3)��=��Y s�!�\z��x���+��}�V����qB���>4VkWcXs��o���<y�P��9p_Ṥ@��W&/��9�uM�T��P��"$�t��p_��J�t���d�>_hC?�<\�kF�W��ё���otm�ʿ�?�7y����:F{1e��k9><����¹]]v�{z��1��_�� !���ӟ�/�y��qjw�9�ذF��%�_+��u���3���_�� ,�2����ɿ���o�����O�u�EQ�����mmk۷�� H��ֶ����B���ʫ�s���NT�����'�IKY�^/�~r�*մ7��Ѿ��e��P�����]Y��d ������G�c&��y}��%7����ɨ`5^ 4E�߇O� �	Y���Qb
	�~�$��"�!F��.��[$���>dBUpH��+V�\�/�0a"���٨".���EE����9?�L7��O�	eB���3&��]�����W���#���z-7Δ=f�3f��G��ȀQ1$#�`�x�a��E�JjO"�
y&Ȯ@� N�p�� ��:�x��;���4���1s\Hh�; �Bs�p+�8�~fUX5peU���г�jKء:ܙa�iw!!��_Ϗ8Sm���K�����S7e�ac�kr9r;L� �0O
C(���2(;����~��W�>��|�W��Ѿ�_d��y#����(�b�z4>�XGR�'��|@��7V�?��}v��MҦ�䌿V�s��������$����V����������+��:���ڶ��^x�����<zͣ�A&g�T��v��;�B���|3P�`&��C(MZ+�-a��fF�׆�P�*v���{�I;L��\p� �y���~ Y�@2&��A@o��I����8��~��̤��[NKB��A"����ƪ��(]<���[�q�FEzd��W�t߃1n@pb��K~y�Rf���4nv� &�c��Y0/hi@č�	<VO�9 	���f�m�{�� O1�����~6ob� $���̲����wC0�d+�ϥ%�Q�Lm2�rʧ���s��[M��1�!y	e�h�y�}&_��i��Ƥ��?�#Y�&s�t�4K��^t$�$�	�ELs�n.�iX4*�sU#�gl5q}��7W,�T.�#.$�/d����D�>H|�?����V� ����laL�����
su6�1�z�:�!�+)��&��$�9�M�=��j�wu�Z졬�=tr��|皥�����x��p���vM�!�-�e���˻&�5G��1K<�@	�.��|�(E�i�mk0��o?v���_j�	�3:�u���LӑP�����ކ!�}�1�>\�'LX(�ρ�@)x1��_>����;�Y����C���r-DR�~6���`�,%<��x}>��q��J�TN��8�tX��A�_5ź���<H��TcJ�WbB��uz!)/�f,�`�ن����R�xK�5�'�ok���|�MRu�X���e�z�}dB�%&�y��׎F���*a�G�-�~N���g�24���?#��Nan�\ݸ�g�28>�����w���2�����5?Vø��ѧ�Lc��A�X�gj��'γ,�3LmkzȺ�� �.d�ɷ�����-}�ϵg���'o���ȒR��!�SO��� E07z�X��#JT~����>��#;�<�J�����8�չ��A�"[,���X�C�Md�,@�f�[��y�PDϽ�w���~��v��1�k[�����/�mmk[����n- Ҷ���mm��6$/�������r$$'�2>�c"$����n����Q7���C^d2�L���}��λ�J /���{>��C�կ#���2(��*7���{��1��B����'OP����
l�`�Ū�D�M!�ڪw��@5aa��d�uSGc�ۅ%kbK����H���7���J����27�B����{���7���#�/u7�:��F7r�%2��X7�;�Sě���	&=s&� ���+�"��a��f9��_H@ �E<���ҵm�M��6�Ù��3�99���[�w݀%��vF��V޸$M�K$�3M�Ł�M+$4���Pis<�� x՝�rfH�5���p���A�&��dv�����(}����OE�7�4�%y E¤d~P��d/����cƳ <#�3�a�a�.���)3Qm�w1���_���-���!����<$s�>����W�Mb�ޅ�7�E��K0!�I�'��u�Ub�9��o5��.�k�4���$a��A��x@�ɠlrf��g%4(��;/����]{�s�b�_�bc����4��dOJ�w/͂j�N�P�bKT޲�W���@et����l�i��dҭR����B�+��|!�|I���2Y���)�/�h��}��@L	��W����{W�q���s���F��Lm@"���y��z7���P,���� L���3�2��.��j<�M��~*�ݞ�4~��d��]V��0Y^,�O`RA�疠Jݴ�c��$���<L;1��`�勭�Pߘb>1mzƗ�`C� j_���[�1��j-Է'L�G�����_� ����n��B��t�k� �(f +/7�{MD d�C`��1�*&_��si����Af�_#��  ��IDAT�$��H�GN.����d��1�I�,�7_�M�
���J3�/Sg��$�l.T�q0Ԧ,S76��|!�ПH,�Y;@b�u�[�7��"�I�ߡ���A^���ïn������X��Ԉ�	�UA�Ćh��&����u��e�'�z�L�_e�v����ܼ�6�,�`mG���"�υ%�7���.�zP���؄�.[֚������^M�����4{��sײװ1�~��R����Յ�����1$��v�ç�����vY.� ����@�X:<<!��˩c�m��z0;�����0��m�G�c�˙\\D�����9�"����Ϸ����c�s��X��?����D
�,�J���Ǭ0\l���D�r��Sk�RT����@)������?�P ߖd�l(�GI��}t������}� @հ@�c��x�C_b���5����U%��=+)��u_�����g������LL1��=��@l���;�ȏ���x�'���_�s�Y��2�gJ�	� ��^'��q�X���+���L@W�@<q�y�k %��s�\��G�@?{K���~ 7w��ʖ�/�Y=*e:_���^���e0��`ؑ�x$7����C<���o~�I�r�Ƅ��ZBV3������'��x���C0� fEpA7�I�Y���o����q+ն���m�?h- Ҷ���mm����nl��>fX7x�����������������4�n��z���ΐ�:;;c�<u��g�tCY!l̰�CZ��-�?�gҘ��H^�	=)�yX�=4�����?�'��P
	x`���vR=n<���.�x*.�p�U�L�;�-$E�ْ�f6�Glp}{��������?�d6[0��\�{<�7�}G�x���?��&�� ��]��͕������i��P��$6���_�R���_�H{Lx�a��Ѩ7�`����`4���N�%MD�8��D�F�lU�iV�\�7E�x$~���p1�K�Q��R��P��hT0�@9�uOy��ϙ`����ͿϤZ�m�|=��[���*�2�/C�0(�����	mj�<4��0��T�*�}������C�Ξ��sG�S�e���
%��ҍ�n��%��|�rU�^p�1i��Kd�I�?�]f������ 4���2��Yq-A���J�$�%� ���7���O(�h��9 %l*�i����UX'����?�4�#���yuq�D��	�P�U:W��{��'Of��#�� �)���&��od��td��0��>Uȕr W���M��+%�V)��Ⱦ��+�G���vd9�9_�n̳�Ы7э,)(uSϪn�T��򊀃�UU��2I���7U�(���
}� �~_�J��s��s���C���2��?C�ç������)��Dƃ�M/b2Yr��  ��&{��v�c�
��� �D�������|�M"s^�֔/�b
a�d��j3�����oL��X~��`� A��.� >��/ ���$:�"�*n�a��L�Uɝ��@�|C�߃"��*�}����`0����R�<f��'\m�5�cl�4��'���S��~�6k���c����4rq1��7\_QiM����F�Vp͆����c��&������)s��������%��!cx�Yn蜏1�L&_���O�r�q��>���k�w�Λ��%��������ۮg��ܛ�A�0l�iq쒽�#�0����{|�8�5��h�5���� �21 �bf�ޗ4��yUaܔ_c,o+V�7��?��{:f�䋗��,q'�Wr{{��V,���Ւ��"�j������	m�U$޻����er�`�����%	9NЧ��{���������	�'������w�zS��~�]��tb+|jܚ��������VH�e���5P�e�y ���cc�1��506�'Ӆ��67ʜ����ɡ�3$���F���o�У�IM
��	A,�� ǖ:��q��~��ۯ����#ςۚœ��N�殆2W�<yB@k���A]6� ǳŚ���|z�q�?5LI0��>cnA>R�o���7#}~) hK༌t���+�	S�1���[O�z�=}f��4���L��2����Zq��gQ���/_�{�� N��3��Bc4�2��`����Th2{�5�sǾ�N�3�U�gӴ7��_�������V����ߕ���9�U��ֶ���[�Z �mmk[���GkH���}~G) �� ����3 q��w<ps�DH�/�����Bu_�ۧ�|:wF�V�\����|�Tx"Y�D)�$C�I`$R��?;;��O2A4�B��E��-̍9�$�ZX1Q  ��1���ڼ B�F7��I��F��VT��%��(1[�u��T���2U?O����&��V4D�;ߑ�����@�4�ߟ�<������P�wr���^�5v��IDy �:cc�{S]  �8wlcX��Aɤ���`��J�eF��Ie��]Y+���	��l=�L@��0�W�O���P��������\	EL���ӌ�Mbƪ�~ Ajz虓���z�h�h�߼/�5�&##��H���i0e���<�ƽ�;7^{U0ɝ:�_���|�-���*>��x�eի�)����`��ښ~[�ǒL��� G�O`b�[����̖7n� Es=.��J������H��4����|���L�����M��0�Ǭ_P�D�}�D�������X���ծ���籠Y=��Ԯ;��KI�a&�u�t{�վ�dn\[E7�,��ng��=G�!s�%�rH��d��	ȃ�s�T�#��u��8������?I��jvT�C�'����VFSN)2�i �%�� �i�K#���`�f�bR=
ٳ��?�����׸�fݡQ h\�ZD�5������}4��x(��1�l�:  �F0Ù�t�eጛ������	4�فa��w21��AU�K&� �C��3?/*��W����fV�J������$|�^���vɼ9:<���=V/6+�/�H�ci�󘂁%|ir��L0�o�]�%#��r�@o}dRd�1B^k^^�c�ŕUuL�����c�������F\���g����H觱!��r�Y.U�|,�� �t@ b,�IY�5ߤș3����L��蘼AJu-��{�a����K���X=���9�:.!����g$h��ٲ[�g���u�"�L�y2���AD`��띿���Ս�
��z�d� ��<�x��c��w� �+W4��7� oL?��(��T�x_�spN�oWi����A���h8<��{o?��������R��k�}��CHn�6hW�w�������!������6��3�a�૊5�߅�荞sU@�*����s��ѹ�w�"��������@���H��S��:�`t��%�#k&�=�� =����<�ϸ�e��'d���6 >�o �s�}���Td�������P�>�����O�~vG����%X��X���L��Q�N9 I� �I��_VnLW&���5�h��!K�9�El��Y`����<#�`�����3��cl�8����<��kx���Ե01���d��� �QL`���M���sJ�k.XV���]8��~O^>�R�7�:֒���ͭ<��5ϞH��ѓ���^r���^B�b�; >j�}=?�0_p�n�,^��`@�<�ɂ�zC&Y��NI�O~������^�?����mmk۷�� H��ֶ���D;?�d�`4�go>�,U��+����qc�X��bqA�P�{��B�a����N��+��P� 	��rō�z�r�������q��"��?xx��| )h��4��� 6�777@�<�����&</��H<c����i�v�f&�����O>�X�2�$�ʫW�rs?���nbKWO|���2` ���}����I8$G��|yyɿ��	�")���P�V��O0@�UݩK�X�t*�sT����2��Jx��a_��R3YnF���IVx�
��gBN,�e�ޤa�@.���AJ'�2>�ಿSL���β���l�%7�ܘ T���}���w����kl���6ڂ#H:$;��ۊ�W�3jʅ`��V��R���v��NR�k}�&o~����pU˨��X��T:�V��1�C��q�J�E%eV�K�b��̏B_�+d=���2�����.�	��-{��Xm���J�Je���8��l�g�*��G� +�����^�KPF�$ۼE�ẗ��\5<5����H�DN�"#���*��e��0�,�|��\���G�3ҖFz
���XqJ/  ��?�9uX�|���O��Y@�;�~\T]3�L�:��8�Ri�2C�G�a����(#��ZK���d�~vZZQuX2�3\��(EV�
l�? X`9�R���zzL$��
Ygr��J�%�`��ޞ�v��ar�!�&���;6��yxP�
���L�z/9jx^P*J�M���%�-������\ԙ|0�06��,	�@�� @,H#����`�6��%i"����� &u�t�U��V�Y�qSSʪ$��J{�K�xi�F�ʳv �U&�Eb�S�82���v^b�6�v r��q�t��+�I+�	vG���g�\��L����?�čǁ�����B�엝�d=�vVm_S�׊dw��c�#�`�Z���gj��^��ǂ�����MU�0�<Ȁu�_��8�3����[��T�6,;�S��^K#���z ��o��{]��y8@>����Q�w=�|��ĺ*��.�' "e+���>� =�c�d�����P��C�9O1<��^�����u}��#p����^bc�8@�?��O&���~��%d��bM5dn����9����y��=r �`���wޕ�>7}��gP�"�$�c�|��}����FɳX�&�-��г8�=����1�)� /&�sx`D��b�%�~s7a�8�?����P�y�m���
e�r}�}{w��xL.�Cq�Ҫ�i��9�n�.܎������}���3.��_آ� r���ݯ7 :���0��9.�}�w�E�_�� ~ա�n��C�L���	���ɇ��!�j��8q�4+<g�M"-��@�Rj�y �x#+�?����1�t�ٳ7��v"��7C>�u��ȱ�>z,��~Qx����p��rZ7���Ic���`ú\꺿�-���N:�լ��n��~��j�mmk[����h- Ҷ���mm��n�Ic���ѓ'�{#&VV�⅜_\��})77w��2Y�73A�+�#J���G����/��X7A��\���K�j`���� �枉 m����3JI��Mc�1-�*`��[��⼆�Cn�Y	�\���Ȥ�0�>$F�������+�������[����z%}}���)�vD �	7�{�Cy�g��G�r���L����ϵ,7k�zLڡ:��ZlrsT��m�#?��(�g +(KUY�׎�i��$# G�$��[9q�(l6�L:Y�L��ب�r д�⊬�oK�x��R�bk�Gf�	����� ��D�9�I���-����Q��/m��dq=i'a���+{���ZT�P��눭�Ɇ���盐>2>�[��aT��!s�y�U4S��u��x���Mm\��@�g�A��p$��$2���i���Ɖl�{FUn����`߽�/�猗M�+��yq�*�CK�2A�N��|r,�N3��2`>��d
�H��<�����R\���@
����C2ժ_k�{H&-��qcU2z�،�W�L(è	��j΋I)����_ -I�d�v�A z�Iۀ��*�+���P����1���C�g!��J��j������c�f�FB�=���q.��s@J�|l賁9Rj({�i�c`!��	6�_��1�>N�R.�ʈ}�㖕{kp������X�[j��t��6W��%��@81 �49�(=�!�X�M��g��qԉ��_.�D��GY�,!%`����Y��_@ٝ`�M�r��5�(�2�(���?���4�Ĥ���sJti���T��
c��Z����� L��x�~~���{�2� G1�̛�k`C)L��c�>�+�`@%�I[���+����`���� 9|j� "�`����#([����ѐ����)�� ���G�����uޫă�X?� Y.Lfmg=���Rm�W�cWa^�L@�[E��EW��c�u]���s��Q �ث�l��yt���@w�T�(�8���Z\�&��ã�%�y�;2E�$����y8�7v���K��l�+&{�46&�n�����u���{Sc��6z�R�4�:	�)G���a���J'L��h$'�'4�����ө��M9�	TW6_9��X�5�M���c.
����w�|��Lgs&��=�ý}>ӽ��;�p��W�4&����م1k��+ ��s+�ԡ30�x�ĠT2ly��5���d���w��!��H Fsc����8�����B���x3�5}��#kz��)�`b�F�s{<b�< 3!�3���5�qq4n�
��6����bgm�̻G_�)�<}����χ�+���:�9&W�&���LJ;>�:���nj,`}��s����QZ�ʪ���ρ4�0��]��,5��\�:�m������D.��3xԀ�,p#`c�N�̱��	����s��ޒJ�)ؼ���'�`N�����nЕ��% ��Ϋ��!^>?��?�X^�xVW�����J��k[��ֶ�}�[���mmk[��A�~/e���Z�us�+$�Þ�f+�x�J>�݇�_�F7//�_��lI�,��w�9����k�B7�� F�«����Uf4}�2} M0E���Cu�U����悔���g4I/�f�{��33"��g�g��֢o1�����(�/Hj �3�s���������|��gr{sC��x|H@۪���''�|/l8�OX
��)V������n";�����n��rzz�M��ze 6���|!��L;�{�ܻ'?���P7���@������|��'�����K��J�v2�/(���
S '�?���zEP���8��f����NR�^���W{��<au�@�8X�$��N`h�[�lZ�Ϩ��BdK���]j�%��� Cc R�r�V/5K+T�V��$�N��#�@c�����-/�	����2�r�`͐�o�gq�dˊ��7�M�u�^po�����P��j���+�CxFZ�|`*[#y�®j#�@2�ҡ%��@�4(��#��*w�$T^[�7 N�W8��iK�d�^<�3���DP����,>��Z$+^���f�Z~���*�`�}
����o� L���u�����B�5Ak&�+[p]����Ђ_?����!�Aq�{0��&�
ZT��w�da���zc��	(ej=ߺ02$�s�{T鸏-�9�������^�����B�AK)��Ѣ�_�&Aw�L�Va��m]��'R�F2��֕  $hq�.i�����Ȋ��`�A���,tP=N��%�G�@k<�c��A����5N
��Ǆp���E�B�mby3�;�Z[��H���s�)�Mo�t���g��Q�0g5�G��@���� E0�u�O<�B�h�A�Z�}�&��<����G;QI�8���"��cE54�u��l��&![A��q1Ir~>��-l����)%�鵯	�� �"��
���(��A� �畔�T�(��Y�@f͉��tiOF�e�Y8��O�kԔ�e��M�'�7a��T&��**B$2DZ�����tF��	B��w��V��G�u��y�i��a� ���$�:�U�>PNr����c@1������-�h%VK�c3!/S��a�T�D}����.����-0-gc��h�= A�qN2x��w�W�e�n�۷�ʽ�v>�? �2�!��N��!qu"���:�+��j ��]�a�6&�l9%Xc0��$�>��?�T��'mI�b���Wk]#[;�����{�zC	�c���H�B����V��@h���W�U�Q���ݞKL�;i�);B=��}ÂZ�a�}��<��Nb�я>��v-/�y�����O�V�$w�(��g��(�Zq���~-��O�X�:���J�(��_e��n[��r*�@L��o<鸡j	*]]�|2f� v�$��8��e�z����u⌮��t;��c_B�?qŠ=q��ú����Z�B��#(G*'A����%�P�y%�=�5�q���
���ʔ{�s��ٖTG�`�H|��s|z_�?g��}@R��,d�,�k9�6d���_GKW(a��"7J��2������q���3�w�@��_S�G�����Ǫ� �c��&����<���/���ev�燋����lh�u�؟3XuA!��s0�Vkϟ+w￈������{����́�І6���@�mhC��~�m�m-����k(�?<�H��Ͽ���Q��.��ӷ�>��������>�}�󯾔��+�"�
�Z��G �������������_�g��o��]7�)dW�^s�u����?9e���Ņ#��c =v�����p�
��eLVq/n�����rx|$�#�<��9>>�{�'��Új���B�1*i#��ђv��U��|v u^��o�@~��O-�A_{}#ݔ&"=�ۛ��,�є�V�	*.�6m�P�>�,���������T7���H�,|҈�=��^��\7�s���]�"��p�����@,�V���������Vw�	��Υn<������P�l��U��,��ز*udA���=�!	�Y��&i��o�?��'9�A��}��h�n-Y5z)����&���
������8�3s"A0b�!Pi6Ff�aD���ۻ�.����*(��5@��_��	* G۪��6!�9H�0b����
k�� ���+Bː������UH��F�7-�3hlc@���z�7Vu5UJx��xN"X,Ԋ�`�����5mf\i��)��б�[�)n�]X>��
v\? �P�W��M���E,�V����/��[�ғ�������=����r�j�
$Q��%�r��U��ׂ�fv9ȠhXm<r�.�X��Y�l�~�χE��t]m��a�BE�~�������41�r���HB ��y�J���L�굮��0���[�ʩ�TTЊ�e�nי�>��  ߒ�����- Ns���H�Io�9�q�E�w�-�5�T�
sp:Y��Sة�5����r5�Ω���F�7@�@|L�ܡ����-#'#;�"�~P�Z���&���h<��a�s�UN7�+��D��*��p7����SA!e��q�Vvu �l��!��O�p���D	Âv��nS$ϐ-����������O �I��՛�m�dиF�xʼ,�Sno��#���
����k��>�X=??׵ֲU�����ܔl�68Ae���gGs�l�`���J�7 ��vC��$z�W�$��d���qo�Ȁ�� q\Tp约�3�ѹվ�l=����:��l�L5�~e�+� q#m��	w�[�9U^PC@9��� ���eX������
uT�3�}>�g��!ɖ��+lP颟U("�6;��R�-�	�ڦX��&S]��9ET_��(�y�`RJ�ܔZ�� a���ѹj�!����j�'����$�� �W�,E���+}H�ffg3y��3�c���̠խ���<��]�s�O�Ӿj�9�'�t%$ͫʔ��er����l��Y� T��e��b�1���c9<<�}����~"��1��ϥ�b���a�~ �Ԉ��N�b��T�@��X���}�Oi 	+f��N��� |�z�`��1�����Di��^��B�S m8�*�c�����2����QF��9		�k�]������:��焪�H~��Ü�>��Lu��euwg�ہbM���bvİq��ei���[�ߑ�)v�Z�fU�s�	֌���ʏ��GO�Y�HƺFP%k:�3�Y��3�k�����JS�3V:�����YN��5�q��1��QTz|���=��\��F._˱Z�ڏ5��Mdg�>���3��?�C��?�S9����9��*L���ŷP�>���J"�0���F$=���s�kS��jG�긓mhC�о�m @�6��mh��@�Z7e�ͦ��2���n)7Ww���w�����g�|�*ۏ?�D��-�y�ÝX�n�(�?��m��租}*��.���o�/���׺q\2�tv�ĳ/bV¢j^�����`�\i�!�@� T	y*�\��;&�A���V�`�X7� Q�z#����\I#�D�r��ݤ-A!T������)�d�EU�t;e���~Ό$m��)]Q\\	����&@	[�0Ǭ8���d׳*����a%q��7��#9��¯M� ����n�M�)> ��e��{��6�aN�����J����Q�M�uT)�B!���ٸ���px����݂�������g}_���5\����"�S��hhY� ���*-C�3�)�B%mL��*�3f��^�AU�Ʃ+�6*JI��@h}��10��[nF�X�g�$��d��HV��ʬt5���!�,�u�g�������@�y��
�
h��~<���^]�
�bE �m�b����A#ڱ�q�c���!� +ޓ�:ؽ���]��-±7�:�����x�*�z%شoc�U1�c@|c�&M�#��H��
}�='��:�+�@�����=1:� s�d��애�HS���IFS�;�kXRU����'���R�3���,�FR��C�^/�17`�rp>�b�jY�ּ�k��ٰ�i���\��b��;��"�����,㹑0�emԶ��7���;mL�a�h�7�� )�k@ �[li�+A��TK伶}�f]l.�}[4�H�q{2��}��X�9,���x�.���Z^G�����*�x��!0�r�!��̪�I.�\w��l�k9O���Q�'�[@���v]e�Y,\|�b5�����X�;���:��0Pޭ�"n�b��S}�cIn�����#��z/�Vo �򹮁Px6s�
�Z�����7�'���~�ַv�]��'Z���S���SS����ĵĚ29*'\��f�@���m����X0{�-����b��5�gB�`����բ�����F�cN
vYF*������G��!�e���4�y)|$1�+�H`x~�Hb_[��/2��>	��q�q.-�F�c,z�h�5I<gJ�%�9�</q �!�?Z���l�֞]���[�6��{T��͓f�f����|{uc�C��:x?�,�z��		��rcye���,�l.4U�P�27���l�b���)�\�
	#���.f.��Z��e$�#��O�7�k�Z�m�����[��r}'Wr�����P��H�����˫k>�@=�g%(.0�L����H"��
�X�X���-�5׮�)n���B(\���$Lb<6�݄���xa�c�a��������;^��Uf��r`��T[�����Wm�?7u���3|����ǙgW���x�-�k�F��!o>���/P�n��A�A�4�T��y��lqq���%��o1�Ƒ^��~�dl$x��AA�=KB,�3<�b<����W�����S=����ޛ����?<��?���2��mhC�޶� �І6�����b��|6%8^�S���<_���X�9�Z�t,�����������kto$�O��������~͊C�Wc�������SѰY�Pmy�[��Fi��1*R��~�j�T`?�M��=��?����l�*ax�=��MY�B�;��k�^ �dR����k�C	��ܻw"WW���2�y顗w���GX�mFpb���Z`W�c@c>B��.��3 ��� ��vG��n�拎�������u�<@��;<+��������:��BǍ�>�K�r�bNva� b���F���d_����B�쏐��%�1���VP�`�c��v�� ���\�H����ĝ�MM��I����ɍ} ���k�w?�kܽ�_A� ��`@�va��k���FH!Q]a�-3(j*�±�c�U���q�۹�O���pL$�O�� 塜)A@v�	^�m�-�M"�����=X,d�c�[z�� ؚ�恿��y�4_�� �XK\��sI��X"d�$��)��!WFK�[�TP�=o���)R3XbT/�!]E"4�	���A�%�eqpH0[�S#���nL�-�5�D�$�8>OG^A ��ĕ۪�� �*�vy�=��UT�W�5������T&un�$A�E�Z 9�l��vr����	��Q����Ȃ�S�<������Ee��AeY,���-�[����k�.�cC���Pƾ�1ǥ�5�+|~*�
,Iv�xaJ� ����y���ZHwΪr(I� \9]���b	�a�����jf��-����ʧ��m@�@�%9�&se"S�d�ml���~-��sNך]�0 `���[�����M��ѶƲg���" F�9��I�0'{�W��A��~�䉇F��8sT���:��j0�3�'�jv@�y����E��r5��U��������ˈ��a�cJ9#+���#WnD�]sM�ߑ}@"��%����ޚr�k 
j<Y�c���d� ~i��ڼ)��D���禞�`�M�KF���P�a�58�kr� �;k���?::��$0�ui�g,q�zɲ�ʸ��_����z
V��:��0�P	��-߼�C�da�����E��=���R..����Ih _u������i?�7_~#��_���m�a?���F<��0��mʹ4�2��Ibg�P�J��:�a�\������π�ٖ�ƣn$�
�lB	�PK9�zM �ϩ�S��y�t�yi}���Yb
�0�vF�&TbF���^1��E��Bf7������`��X��0Ǣ�ϛP�B�׸��l��777-�nJW�q������P�NO���)����A�u�
Ȏ�sE���<�"�s=�H��Ơ�s��"����綈jU�°�����t$��1���;o�㧏��ڸ���7|���-��3��C�� �2�/9<�&�>�s]��$9_nF�~����;��[�U:��mhC����І6���wުj%�*"g2��Γ�����������|v(Ǉؐ=��&����)X%<y�H�{��pTۍ|��y����,�X�����W����Rk��uQ���V���M6Y�h�F� *�{^\��b�O[�2
6�naM����,g�=�Hk6�����g�ỵ�ziU�׮+��6 zL�m��+�ޜ�����(.PX�� �l!��(�����-K#ଋ�Z'5�4�K$M �Y]��6W����k �42P��i��7�Ty��R%�`mT�o������a�z=r�4 P¥��q����,�����L��潔��������-��r�,ɬb��ɉx�����}�9�4��l�P;U��L�Tx/�M�+/��	2��(�·>��0�W��� ��@��f�:f��]�>�ß5m�	B����*k#��`!�-�g�~��	F6%Xo� ��*&�>�}pJ#ف�����Nި��ɡ�Ο�����U�ٴ�q6&��Fk~>�b���)��P�J�U� QՅ�WK�%1)T��ke��$�0�y"0֊[���Z%ɡ
�iP��ƙ���}bppg*�,;�-:��L�ձr�i��ёd�̪d=$�:�r��l<uT��p2t��f-����ށ$"؟�|��xr����0L Y�yfAEP��/s��П_���{O��pƾ~u}億ϡ�Ki��	��^�>��@����+�a���B�����mP��zn���<�%��L��p��n�>�X�{�3����W7B�a�ɢ3��w�j��50�m�~�*���$  �%��i�r���
&�Zlc��/W��$�g��|o���1�{PL�cW5�Cu@�ʚjō_�]�x:'x���9v�#�
^�x?�m�B_�q�%�-~����q���m]�ָE_�J1�;��(��<��X���бr�p.x���
���@�@p�y������K���Ɗ Zs��瀮k�y��㮷ė�±�������k����ؘg�G���RЉW�>X;�v�����5�0�8��}y��ocl�
m�������x~�s���F�t�a޸vO<:#A��M�	t���*F�� ���*��|OY@�Ȏ�$Y�Ъ�>���֟���<|�P⧩���>���z�:l�Y'e|~��	�$3K���&�ce����n�� rf���.q��n���aח�����7�a'I�|S�͕)�B_˦W�T�[aE
5�Ui�t	�M��kf���:e�
��R��d�Z`%�쪖
�Z�^�J�B�$I�Ԕ��F��:�}�� ?Z����-��q�B=���s�G�6�S�J�g�,����e$��(�Q�ϮwqO(����_�c�]d����r�輔�8�\���B�xv!��pq,g0Dr[�$���_���s<������P�s@B6���bx�x�������v"G��t�|��;����jL�l��6���{�dhC�І�{h ����b������ޓGܸc���b���>�H~�ӟɓ�?�?���-����z��1� �ֺ�~��[�!�Ǧ�/��/�n���O>�������us�vH�A&��-�c��r�m��cOJi�8���39Ʀ_�ǆ��
s 8V�k������ӷuc}+�^�b�c`aO!{A�MdJ�[���Um���o�ް�o4��|���6�eC~���bm��@wuý�����4TYeV���Q;��N4��Í�hZ}�O�5�:R���&jݖ����n�1e
�P�*Tp �����F�BW;��Z6�n����թ�ivXA	�oU�O��;�@�6�ā(SBe�>�A����ł�]Լ'�ޟ`vY�<���^_�*}�&-� ��6dx�6@,�2��q4�88($��� ���I�+/� .�Z��F�{ �xN�k�oqO���Q�/ )؅j#�Q�^ �`˴m*�8�{�C�2v�Yյt�"c%2��<-�`��������S����O0'�{*,M0g�@��D*՛�$�܏�N�_���
Ѥ&�A�: �P�:�L3�R��W�*��^���=V����(��s�S5A9 �J���`1���5�˒8v��X��W��=��G[Z�t�_��E� ��,��	�mZ(�x�i=�_	���1���\�'�O�'TlX�L��֕����\[�G���/����hJ��իs��1�)��ǧ�q�ٔ�p��A~l6N\�;�#�!�_T�{�k�
��a���`� c;t'=L�aa'B���>�О�@�N	Ċ�$4[.H�A>��!)܆Y�����7v 5b��"z"�r�N��4��q��*39t"�}9PW2 ���Y̺�n������2����@��=�X�@@y�K�XK&X��-��5b~���e�����UT�`n0��+�ͷ�	\�y��5e�RBr	�"�dG�#�|��/\�P�	��{`�Z������r)8'{�I}-�|~i��/��U#R�'��K+�����Qܯ�N0��r�ɀlZ���k�/
��P����,���"K+���kbjqU�שH���s�,�z�����/�����}�8��[}fZ����Ǧ�E�mĲ�P�鵀
f����!o��z��O�oi널��tN�
PNO�qMĜ��3΃\���03vJz}����x��� E	Xb��)=�x�_#^G�}@pQ�1%�N���N+Q3�D�9�:
����/�H��Ʀpcyp�H����u�1C���*���̇��b�bK]]7=Qb���+--�l^��,ۂkK�q��>[��t��s�suoӉ�C�JY�3�!r[p�"�����q�	�9UyQgV��l���6+<�4fs�k�[HP��X�#�#=�\�G�##i����-���mǹ�6�h�/�~�-���+g�J6�1��hZi�������"�����/�2{0��y��ZB���l����=9<\���L�٬>u.��+�8�v�����\lhC�о�m��6��mh����m'DoZ˶l�n��t�0w�)�~���?���?��,ǒ�RGw�'ˍ�����5����MX}:��5���$a����y�6J���ol�i�0t2���=�8x��Jyl� ,mK���FݪK��Y�Z`'���(��W�%��'��C5_Uu��&� �t�	�6W�~Un���$	 7���<Ѝ�S���� Y��ۗr��̪R[�݆Z5)T�����q�AL����K�z^�z!����Pth�F��Tg�mKӶ*]�]���v'�ġ-�+��zl�QK��1�&Tn�����Jֵ��3S�lZ;?��A� B	���
7�z����֓ n�@.����+�zP�r@¿#Z;��x63��[ÄJd#i &�9���!�& uv,I����p��,��_>('���L���*D~�>oʏ�vR�}�=�+(.2������e	���}���{a��h��`ٯ�fU*+��Z�G��rqy)����M�;��z���xU��džNP��X��]lǔ䲮���{0�k�tIz �,Pޫ�ᡒ۟]|�-� ���Jt>���!����1��[x�vk�>��n��1�u�>�#�6�d:�7�Q�8��ބ��-�S),m���{zz��<wB��k{E�����j-XX�zE:�m�c��!�me�.���<�͖c3�A����s�BV�AeZ���y(T�m�6�� 7#�Y��=��o
���W�^_^�U���hB �.*#��{�bۏ�Z�\q���)�����=n��<I�.�ρJ�$${��{s�iҔ0G�뚘�{R��2`h����
�]Ph�ma�1PS�t�8���8�RS��M�g&�
	J*΁̜�Y;a�� 댠�VW��'����ɹ[�}E}k�BqT �W�	3��^��3����rɵ� �\ˑ@?��b��c���'��V���#�C���p��ø+��1�,Y�aD�}f�N\���]P�k�[⟃ף� �MKMW�����{| �xH%�O��	�
x-�ݎ�:bʬ��ae>��?c]Q��l�'��#�[6�{M��Ҕj"p�Y�~F��a�C�}�s [dڈ�ؘ��,B������gg�:���-]��%AD�f�Z�A�a���k#�Dk6[�錤<������ʧ�}��x��>�ʣ���l���!�|}s�"��U�Q)+�lln��2���vn ��o8>	�w� e��0 >�]��4��)�pb�4�(0��5���ZA�{
�ԧO����}��c�c��+cW�u>����0wāL�~a}�e���b�)>�N�?yv7���s��Z���^7Eg:���y}YSE��mI�E\�u�Y������HʚM-�&6�pmnw
S�cJNn9��^��%�6G�/�N|u�AfǼ]A�8�g�,����g�XX��3ؾ��׿�_��o�7��ryq����N`Ŧ�a<M�nA�1���'?�C��>�llϱUQG��"�����K��'�mhC�о�m @�6��mh��V�M��Q���f�%MQ6�����LG����~�s����T>y"e�tW��U)��j��au ��E!���?�06���?�_��-�+��0�%���F�*�(c$H Q�s\4=����ؐ���
�4͌����?��ܰɢ�ҖP,6���A�<A�w����<�`æ���+��#�$�M���@����U��_^�x>%��F��A�9�ɷ�YD�mN�#�"�n״�2Ia-3&h�m��G��l�>�<�:]��]t7�wߘ�z5�<��Y�V{D��
ce^��$L�U�$�@�P����0�3Ty���V�~�X�x ���?������s ������qO��gt�v����m�Ze*8�	��+�Ce��^��8 ҹ���w}%�yϖ���Ǆ����z��8Z� ���&�W�a�� �1({<�6 �A�5�DUC"���R�/���Cj�??�8�� ǡ�z%�^7����L�YG�L_r�w�Xe;+�a�=�- �����.؇��������ߝ�� ��,y-ұv�['F���O*�W[�FXli�
���I�X�9X�̞�)g(4
3�<�%�P1�����3�&�p�``���s�t.�׵N��@�5� ʰ�c52��3��dq0' �T��?`�zޖ�Ľ
�8������1碂�_���M.2���t?}$ƽ�[�I���X��)$Q���@1f��+��E��|m��SPz�98�f��b������6^ ����
*�|�b^�Y˞�A������@NX�Ft$���x73���w���$�ʒ�-��@�;ZSt$IPsX��y��_�۸�Q�6{u���1 �e`��^fo̖�>��@���}�e�D�j�~����\Ӊ[���{��������M%lS�S�rˤ0�ES�`<�ny��4�0�ŋ��-X�>�u�Df�1��'�����7���j�`?��Bu�e1��x���ށ��3�x�Af�+�\�{:䠠�yJFV�{��e}��Th�Zf��ơ�y��`��[j� _�>20p�H۽ut���l�Dq$}�š��������B����nY�ݐ��OH��t.�f��?P��R����{T��a���I��W$~�S_��T����믾��r�L�-�͟���|�͗�ub.Zj,�9kBC�'�U�3 {���^m4�9���"��hw�)󭠟��)jq˼�2�����I����Ձ(8Y�$-�tX��FJ#����}c^ՈNƈ[-z���8��r��uYә�,��@.͠���p���^���z�5O��Z��#%>���ϒ���H0�P/�5�5�E<������N��� �/�������z>KIU��s�"��YoK5H�"��
&� ���#F�
0�?fs�����%���uu�Z>�����O�����Dv��-W�Z�`��x�}"�K���kUy��Ε����<l�@�mhC����І6���w��4��It]��j�`o��4ݗu��goɣ�O�?��?��-���c'�T�Y� �%8ҡ��26�A���Uۭ,��?������o�~����h<a%�$���s���� ��@U��q9��Z"����1��?D#�Ǡ%Rk`N]�`��W|:�7�6F .��*N��$�?;�2@�\_\ ��8'�N��@Ԫ1��P� {m Q��ցp���Tu����@:|%�FMqE��X~���}���Y_����:&no�Hl��6�;�bI�ٚ�N��#�'a��}�n�s@��)ZUPbU�ٕ�����גݏw��G���2�#ة4�c��'�t�X��j�����@��5�7�ok��zH Ȩ�ɳ� Bȝ	��]誫m���:��n{{��������K���P���wB�G�s 5he���O�k�{�����B+QfW���y�U��� �K�@(q�t���;}_w%�N����Fpo��)V�w"�W�b^�]Lb *�r� -퍘qa7�M��'�FQ�X6J�b�߀��I�o�}�q �y�R%F��I��HŴ6K?|`��d"g�N���5���l>���T��.f{07�B_���#8����1[� s�-�sY��D%=T,�q�N:����Fڄ@a�VWh;�eFT�f��s���P��J�,����~��b���ϖ�3F�9n�֊����.�����ȯ��<L�x�F��x��jp����@;��d�j��V[�Wh�I-����0o�d <l��x�����5�bP�ECd�;�T�L$���l�5���?�*ĲG<nu%ׯ�W�spgs�(�M���6blX-mV����u`HzB��Z�����9s��T�̬�9D���L
����&��@��n�϶��37�Kӏ�0���0��j�����?m��R��a��n�R���� ��}��E �y�Tn�u�0�{�@?�7�/;��?>~.,�<3�������]1�H��2/<��|f�����՝u��ݞ]:�Y�u�#�P�QY�Z��HԵ�0�A�7�nol����ZK���μ*]��FhP�:���3K5j�^a�ĺ
�+���@$�`���R
}�A���u}���^.湜�z��jkj�/@��x����Aa$6��\�L�rcd4�@*����tK�Ɲ�5!x��H�o0��`;��/z��r�����!=�\�C
A� >c�o�}_I<�)�wĉ���1��`j�=�_$�����J	skQ�3Ĉc��I����](��g$I��=�����Fү١����ߟN�^����3G��j�����@�9�����~SrM�
���A��v�Ͻ�93a�w�:�paA��<V���u��n��/0�k\s�ڔk9?)�>wv�\�6��mh��6 C�І6��Ck�����R��Z�Lg�9��?{<������O����X�:�,���f�lf�ہ tl�,�����+ZI�n!���:==��vpVi|�8���� �7�?���5���I����>6W�s��(�Ϙ�6����`wb6���i� f"k�A#F8�%)��Ңiv�\�n3��s���0|}y-_~���mX��p�kTs�[�I�9!�mY�� N�r#��R�w�ӝ�;����p�W.�
���P��¦�l	�n6G�T ��\��Z����k��4�`C]�IH�ԝl���P�n�-U) LpmQ���ڦ�������Y��hBjCmܖ��  xMӼ���jr�9^�W�
+�;���X!�{�r�5��P 7 A$�{���,0����G�����q�8��xm�oT��t\GZ�$�gy�T*����n"��^�&�b�¾�d;������!w{���k�j| c����¿=d� �M0Ӭn@���c���*���e�mv63 g�E���͚G*�ϦܼA� �U�f7��U�[�+�\�{,du{�ϝj?�l_�`v�M��i:������V��X畔���TB��b��]s���P����a�1�_�	�yo��z�s�a\�C�����~���?::��ٔ����d>8���'g2��Vz�ׅ��
�d�3z����;m����HG&���΅�B���Z�L�����؂�?C�iRl���v���a�5����L�S��h�ކkf�mK`�u��	̦￴A�)���c#g%1�a~Q��	��=�t��ۗT)$�]���MOL�n�\6���#� u��w�B�f�8�}/�]��T)e�k����H����AB��K���l 9]�}���,��ӿs�
���,G	�뽅B+%\��r��1��������fnc���[���ڷ�ONt��g�}.�^�����Z��~Ȋ� ������G��T����X�O��kHH�v=�? ���X�������}�֍׶�y���k�.���'��`���3��[H!L٬�F=��Op�_�(s6��Q f��Q� c�[�*3�0`������r�E�<<��|��>��L�i�A�����?v��s[̟s&�~]qNMFsS�%�3�3�	��*Mc�o؀$�w�Gv�3��,q�Z��:W�=JY�{=p�X����% �:?BI�s��v��P!��+y��7��oy�O����=�S�C�g &֛�����<)�1����'���{��V��k=�-u X��i]�*eo7�ί�8��X�}�g>��=.��mF�z�}�J���@͒$��cA�)8�V���2�}㞅��o�t�7�'�����g��y�`��-�8��;�w��kTG�E{��������:�n��#�\�}qa�����PG$����>>����-�l���(2���*<CC�1'I_0�Xu�Ssq��]Úd5�]�̵b	rD���J./_�G �ӜE ��O�8
�SIbM�&���T�����oQġ�uv�P����L&:��u
��t$��mhC�о�m @�6��mh���o����ſ�7��Y��/t��B�[g��[<x�t���[�#��d�Æ��V���Ky����ח��yE�峇����Y 5�ɺ���f���D�=}G>|(���C����k�0���Mx
�ju���MrclJ{�` �ګ��Y�D��C��ѯ��R#�����T��!I�Eʭ�M��Ky���q�+4*k�9�a�sx��!l?3?Q�F� 8#f;��6�T��7����~߲*������ot��I_��6╵b*@:P����������`�`�
*8�k����8נ���7]oEIQji��A@��!�(�]�`���x��c���s��Z�e��챾K��}8��j����6��Z���`���UP֞��Uw��������n\�]�G�W55D��dJ �D��q k,��)/jIo��v[��	
��{���W��f��YK�<�@ʄ
�W��qL/�Mp���5�?���}�Ǚz��~���-��f)��c$:�7�7���c����T���Y��F�F~�Z�i�o;��]cVͣښ��VQ$��7t[��z���^���娠a��7v� v�:��\�v�"�z|���l6���?id�Y�ߝ ��a�:w� pF.oK� ���A �2 ~��Zq�Mij�P^H���3fvȶt���B�'9I�U�4}���k@��jP 5���# �ʣ}��?̗IR��G�W)�����I`+]����\3��T��aN3B�2����7���+��a����23>!Sz%:���s�Ds-҉+{l@4 ﴫ��$i�c�������)�����ÿ�+cޥ�>��y��LX�8w�NP�Y���� ���y n	�ϋ�sAu���忓AN{!�'�C�ٜۢU�8%7�\K2kW�~�
���	(e���_�����}uEP���"ʥ����M9�9Ȃ�j�q�y7(FHX���,�j�/�Fk?�<d8��JS����8���gv�A-GK*W4U˵:Ƶ�v��$tt�v�<��(�0�"�GjF-�1sBп��\Hk)�da0=	��Lpn 0OP������jg�죐�c㱅a	z����AXW�2�$Ɩ�+�*r�u�{�t�9���?���[פ=h�4��V�Ҁ�M���޺ �1��TQff��Az�O�xi��g���n�j�0�)��	<SL0��׿}HX�����v���3'9N*Ŋ5@�m��1�"�Ob��d��Ǆsk��o�!���u��Ѥ�I2'��b���X�<���3]n�����}����9I�@:���#�_��N�t�sv��0%���g��m6�cf�\�_�'�|"��Cy��)I��t.���|�񧴊�����۳�d~�w�Fa$���ӵ�X��g(��>"'f�����ի�˯�h�z�Nm�m5:��mhC���� �І6���^Z�v���y!M��g�N��fE�]G�n𒈤�+��?�����A<p[��g_���Mt*�G���b��Ǧ��wޑ�l�X7���B7�#~��+�6!��n��6H�CU?�ֺ���%P"�&����u���l����<z�P�%�F�~���:�����I� ��V~s�<��c�Ʊ�iG1��X� �@��v  ZA�P�Y#����)+t,�%	�òͽE���h����,�(H����⽭a�3O'����3������B�U�G���g��A�1 h |r�`�ہ(Y%|ʟ�M��Y��>5�)�"�����^|읥�~fl�Wx�8�oᯥ�@а�'(���F����z��
X�H�A�Z
�A�m��,zP�����( n��݂�YI�@�P��-�����f�U\���h܃|�G������٠����M��(͝P,[�n	�H�����e���&�����L�i��8nW ���� ��3��~��!d�hߑ��^ux�?ߵ�AVH����78���CK�ĈX��pϓ�Y�����d�������J�mI�Fъ�Ĉ���Y�L��a����"�x��8�̗ԏ�|��7�_?X�A����3U��}�j�?�U��L&Sd��m�o�I�̕52��-A�)�ו����1�M�e����� ��;n� :�ʄ�v=����l��!���¬��g6�b$v���0f�b6އ<K���Yگ�z��D�>>A4$ubEc6@�@�RQ��6Z���ui*T#W�%Oa�Z�[}�=
��BrK��&� i���3^�G���B�v� �� ^x�5��m��s�ƲHk�����r���������.3�6F�$X۠V��
�Qo����-�h���J,W"�ȃA��c[T�.֫��銘��,�0�1�ʀ�b��XN}�A�zUZev�w�5"n<65����c�C%;��c-�s�#������u�D����Y����������� �޺�.�7[_�\�6ܳ@
��iߢP< ��lN�4Qe ;����'�5c��7��c�ezc�\��������u�:J�rS����kw����lM���`��ɡ>�,t�0E'ք�6���.2q�j�h��8�2�W�֣��T�0��ṗ��ҮUbj����r||���m�rmd7��Zm�^�U�
����ǵ�-N�%��`��x�:.C��[ّFN��-�m���l+	�v�Db|V�}=����|*!��k�l%ɔ@��ϦB5�Y��6�܂,���Qd�a�$a�k�).�Laue��1`~g�v(��q���Z.�^���W��3�ص��x����H�B�k~C�x�[ǅu�I%^i�HT�Xum�`ɇ�������?^|�\^�s��ٙ=��}����_���<~�K>S@�:�b�#��{><�gO���+����畄������>�B[�u+\FQ��X�6��mh��6 C�І6��K�w����������8�.���}}񪸾�j	�o���:��o��B~�W#������a�/�ō7d�M"�͝np x��3�裏��=��f౹p���WMZ��@�W�X �=� وLT��5 �`K.H�Q���V"	�L��Vܸ��8�J����H&��L���*���q҃�!O���&� �0��;	������V���ҟ�I�4� ��?h)��J̎�$��6��w��ӷ���� �ƶc��RV��"�##rh�R��a}�0<7e��0N�0�|��.QȪR�_6�_�O�pv�/	8'=��Od��7[��?����(786�G ����(T�:���!XL�=�V�����*����ҍz�T�.�;���'�1� �A���j:x�Ӣ��S����ob�;o��)�� � ��J���@4eǌ��U8�p�  q�'�9�<���VIn���>��.�3B��3"�v4!�%O��V%^;Y�Jd:&13�g~�Q�� $*z�BƋ+��(��Y�DIP;��4�Ǵ�� ?z}0	��~�
� ��{x�Su)�Jz|�`z�cn]!��z}CB�le26"p�����e"zʨ�J��:�{��C��X�똭��O���ņj�mY�H��H�� V +��u�>���H/�����۱���#���h�����5��
�؜p�2A���r�y���ؕ5�˃Y �d�����H� ��˼x}uI��N/��Nx�H)���65�[�CN���CIU�^���VUn9��q?�nv�2�(�m�{�v�'=q�u;�#�SZ��r$�b�Q�#�A�F�^Jx�X�]V���a�!?�o F��3��Zצ+�fP��όP�`�I�y���7��@C!�s�[�1s�dނ����4��`F��1f�h?�F��a�>�����DZ��}��-��>����x�+�������֍ή$�#@�yAݑ����h�LZ�ۃ:-d6�W�2�a� �c�*���/�=z5]Me$�Ơ�D`4��,*+�qbJE����{�I�k#^S�܉����Lݘ�� ?�+F|��ޯ������]�Z�Ĕ.�� ����k��3 ��=���䦘��0��JK����@�_��Q��{���o�1(pi���/?�5 ����5Ǉ��B��d�[9ᙠ�Xh����h�ϖ�Cۆ�PS�`RFP�ڪ�<��'�����{��@a�X���6�����Ҹ��(=s(�����6kI\��`y�k�H��B��p�B��JbS�R�����ڎ����^ۂcϥU��Hx�����Wgd.Ӻ(��)�?���l��Y�b.��+,Y� �n
�rQ�g �S	��젭g���/���}&���~S�;==�?��T�������ua�IE˺���e1����!�3�{a�����?o!�����z���fU�І6���{�dhC�І�{k�8߬�r�������O����u���.M"J�G �Y���G���dNU��՝mP#�{8:<!�tu{+��W���f���*7@�!�B�T�@j Ea}ӵ"����
�a�m� i�r����4"b�����Grp0��h<��+����n��/.���%	�vC8���#V�e��<�!�461�ul@��Z�OF:�+���*�U��t�f�"HY�"P�J����#���S����ݭ���P�����`mM��k�j ��\ � s�4�쏘����%B�ad�����۩0�X�7랻v�JW�r����K�~ԍ�z�۷��>	¿	H"}�q.�.�W�D2Oe������fV���|ԃq
ݎXʨ1�W�vC * M �`�����i�_7����z�g�F`M�-2"��U��.< n<겷p�)�vd^���e���EAK�գF�>9=5�����w��쵩	���;1���K����`�aU�mO��81��߯q�3���@=��91��w̢J���v0 ��ʫxݲ��Rb�c�Y�i��?���G�v��<�UǴEs�
c s�,���Y��-l:d�@���m�3< �AMԢ4���*�8j9>�8� ��)���byxv,��	�8ܟ�+��N�`�YE8��;��R����d\�A�����OyBn�އ�v`uLO�J�a�_3=�_V�G��岔���=,HX�;�= �<������NZ�!kB8���<"�+�-�$�v��9W��g ���N�Ȼ|}Ū_��N�	U��b�ϋ�2~���y����ʭrDLt����o���r��@�����`��8��,\�x�o�ܤ��KP��$&�1a��x:������X� x�;P� '(�|!|�\12pW���U0�^�>�G_�z��0"(���"�+��Bǩ�KlT�ņU�v�H��^��a�7�O"X�A%�\W����l\3\��'~�1e���������>�,�8?F��6޲ ��mӷFQE�[a�nKGf����s�
۾="	��_'�_���}n���d\kq�INiߊ�3Y��Ξ,���"q���ǜ������[)���VePj�i��jd�Y���V��Zףk�g�C�w̩vR�M�<���Q��.�u��<�@MX[Ş�6�Ή6vJ�����S^��������''ǖU�_P�9����W��z��n��@��xc�DP ��u�~�}���\���7b_�}�bV���,'v�ӑ�ر�N��R�������j�c���f�ge���qi�\�ϒ�9�G�W��<_a^E>搛�>?���P^���Vk>C�ss���)�`�
iK[@SU]_]˫W�HL,�N��zIҔ����3(l��c���s�+�=b�+���7�w..u��b�Gb�lX��F�����dZy}~!���/�~H;6<��~�����Cx���g�r+I�9�
z���¿������'�|�����w߽��w���N��mhC�о�m @�6��mh����K�4���F�+j� {
�$-����G�ij��䲯���~��J����BY�IG�5 3TQ��@uyk@�fca�7��M�t2�Mp��ޯh�(NN�)A�'�2��믩rhۇ�L3rH%�RA����J����Vu��+�� Y�n��� 96| ( ��j�}�y��z���N��#����m �xB����)x���Yzdj�b��n�R^MI�!"�`Pl�{�3��	���|���ܫa��?���@��EVl�ة[��Hڠ����쇍F��Ye�
6���Ո���77���MU+��`��P�~�ǭ��4��Xe�Q���a<��S ��|[�i��32�����0W�h�u��p�+�[��遶��a��DY X���E���� ��v,��@v�x�� ������}�/��nY8q�.6 ����*Ҹ�cL�lkx����΄̃�0��/��,=vP܃�v�<��2��(���G1m���'6A��Qg�+�3��P��6] �PQ�#t,����F 2�� �_���$�9a�Y�W��<b�MbU���;��P]�s��͇5
T����A��L�yB�<�&��ñ$c������y��9�p8�(�+��@?z�G����IB>��������R��|���Ӂ
�� �`����rD�Y�AA:��kh��
���W+��w77���_�Z�l�zPAـjrڭ������\׈�;�%��8h��;�h��9�Z���9bY�{�6Y�)�@nAaU{Ɓ��Њ�����l	�>o!6{@��>����-�qf3�3d�ɶ��R�<:��!ӆ㾡ʈ6U�)���C՝(�Ø�oI��u��|��r�l�	U�$\`?��28\b���9�4�r��7��Ά����t��N'��������0��y!���[�S���3�!��������<��+�k�n�9�$wiYBP��1��#I���E!�)#�1�9}���Q�i�y4�c��PR7f�g��qh��>v}N�7ʨ�1%[�9
�ǉ���|�{@M��C�W7|���K�曯dv�`��8�s�#8���AQB�����3�y�󶚠n���s����Q٧��`<�׋�\������e�k+��NN��J��j��0f���nM5�v��Pl���uq����{�&;L[�8�P4��}�2o��Z��� gLM��. ���2*@����<�2ĉ�I�$]ޓ$�m��>���J\�2�uσ��״C_���:�^��zG��;!a�5"��7,v��<�>~��
>�E㑯�֯A�wz\˕)Hp�p�p���	Y_P�!���������Y����� �A��Xi��:��Hv����흼��9�B>��Cf�A9s��cPx��3D� �(�B���|f��8��^^\�R���k���［���ϗ���������\�6��mh��6 C�І6��k{��W��?|�;��V�_m����N�7��O�Pnn�I�F>IYAZ�6 ���RR�X����ީ��޻!�o7|���MG2���I�� ��� �u`�XI �v!�
[d  �`�x��ח�I]�1^���)�T�&� :�� ���Ͽ}A(؉@0B<����u ���g=�2�/��U!P�\��"C�$3od4��"D\�W���bJ̺!` )�s�5�¬�`�R��VK�FB�����'�c�6�@;��E�<�	 �(I��EE�m�kV��~�z�!�o9+�]To�VB� �[� 0�*�no�7H*�V��AGh����Y�@t��w���^�Yx�ǅ<=Xe�g9q@x{��V0����Z����E-���b;����?�@�(*`ƻ@Z�`!��>]P6t;��c]mi���]Q�wQ	���Af�.[��}U4��t�~����]�{8'Z�$F��㝗`����#~����$������~�I�²��}84mټ�U�Vi^��8��lh�a�1�kr�!�{��7�AVbK.�>��:�z���❈���4C *�֔W!���]&�3ɂ�o�neq7���s�Y�p�����������}L�9��<ֹ��|�&��cvo;�F��m_�NUC]����V��`^A��G�:<:�/���v* a?~���8@����5��K�Jb�	 {��r�*(�V �ˊ�>�2H��W��0�ї��� H��u�u���,ǬX$�����b�c>Mv��1Ȼ4�bʌ{���B�F�{���"�*��60�u��8O�x�����-�ď��#���5o� �A,�!� �K������k>�|��-cS�H�j����͊*��cc��tJE_��cc58_�q�&Y��,'��UU��'�X����TP��9�}�J71[�T��k���������)���?T���3��* ���!�*���r����pO�g��c���na���yw�y��`x���Y���ڑ�a-����H�I���v�bIۺ���Ui�b�ǺvFퟓگ�p��(ض�Z�j��CZ����ȶ��y�(nn�@��[�<yҫ��� ���<��s��X�V~����4�ux�'jC�-ۊʹ��Xeg��)w��r'�i?����A��u��F�=4B��F"��=1E�M'�pf\���NX`�~��8K���Fm����kk��9�i��
ͮ����h�x�z[�y���� �$��sؓ�<�6���0Xnd���d�3��N7:�b-x��s[�B�ϑ������:�{���-;*U���kP#�x�\>��39{x�ϱG鉓�9�nY[��"PX��$�+�Y�8�C�g�ϦE���3u)�rwsm���X��F
�Ku�y����÷���B~����铷���GrxrO�?*��w�?����Ye���+;Vz�(��~[V$?�Ow�����'?������[�o?�����jhC���;h2��mhC���O?�-7�؜��?�tcj���nv=z"���rs�����c��72�e2�ͯ0�\7=><`eY���_<|�r�	��I��K�Y�����Q��r(��7�fl	J�=b��n�R����r���˫sy���m�u��ʹ$��3��r���d˄6 ���Pܭu{"�E$c�y|rD  �� A��
ʖ��dy���Ѝ�(����_� �@(0`�cn+"�C�Q 2rG5�Y|��rC�gv�_����Ō�.�ꎹ,�ojkӮ���GY. 5(H��`P\� V{7!��#P�@0*;����mۃ j�ݷ��I,�T�6�!w ��GAlKg��H:�%�K�`��Kz @w������&�]o���T�$�X8y݃h8�G5{�k���Y�t=� � F�� ��T����&dct�
$d������Hn%� �����fp%聮.(_���-=x�?C?�tT�[i�i����n��D#�vd�d���$��ӫ������F�ҵ�Q��Â����i�3x�P��*d^T�ٻ ����n�3�!��u1T��a�Ce�< � �������`��y��:�#fM%�N��BH�T�:�oί2�k�cn:F^FN����J�- ��9Z�<�x��0v�2^^�M �+����m��UU�ZX�p�X�\�%	�p��O��~������$�b��[=^�i�s�_�,Xo��z��f�n���r��J��k�*w�#��,8��|��F�����b[�=do���>���:>F` ص��9�� t���;�LI�WF�@9��y�=�O۴�������"�;��c����²��-��%� A��2_7� ��t]�y��|1'yq�����vM�aQ��l uԏG󀋨P�j��Ú���S���I�C�k�|C@ה f����2��\3h�ӄ ���#k0�͆sX�G�����J�x��gJ*�6i�]fAP�IP���1 ��N�7dh����A��H��#t�:����j@/@�M�~(Yٺ#4m3�%�9.��SC���ˈ��2�p��N�n'��Y�����EE��z	�X�p[6˵��zE+8f�D#�),{�d���yPa$�i��ŚDJX��X����N鼑�!�$6�/ﶖ{��T]���A�'܏��'P�y`:;����^_��/^�=��]6��9;�b:L�:�c��zi}$%���/8����%QN��k--�Lbk~�{�:���cvS�S��n���Ж:O�r��[�����p���
S@�֞k6�EW�j�k�J��KZ�=xp��k���0 ��XڬB)|{s�kGI�!V�8��ϛ�������?�%�٦`����u���,\���33�MPK-����t:7����3��'�η�������]��s?�}�6��<�]3&�)���[��_�5���'����o��������}!ٰ~�b�7�̷#� e�����ו��o?���u�kw��}�~l�� :��mhC���� �І6������O�������Ź<8;#� ��t4��~�3������Ms�o��n�Y=��u#��'�җ�@7�_�9=�ᑍ����Rк`���Cx ��j�Y���il���<Y�[y�\���Id���Q��m����5�` �d�;:f�B'�)l'"y���'�;ݔ.(�?�ױ{��@���U&cT�1 �����\�p���@6��&2�F�a���܃��L�jn�A���'�]�<���MU̣e��6�otY�?�ɒ%ɕ%vm~�����J��Vw�����)䎔^P(�)�s����"�Y-$���	@�L$2��1y��f���ܫ�^d�p�%�i�>�g�LM���9���� =�]�����}@od ��ߟ���z��9�G�6'ࣚ�-A<�}�(�
�1N���saw0,NT�@�_PP�T
͜$P p���wK< Rd�*h�o�U�p�K��j�[���J���ʐY�e^�&�����=*��Q�ѻ;~7L�ƿ��*�bf��xgFz��- �d��=h�	,x^�m�4�{��"K�u�@h��Un"�{Mf{"�y���{h1���|D�+�oo_���d>[��W��ao�T9)��;;I�0��@J��$8o��8�$	^�������N�����j��k�
�(��Mjď��t�GGN0d2٣��/]�.p����V����>�9�p�{P�<���͊lb��!�?��<.F�ZI�M�}�	A��l�(j��Ž6��^=4<GFr�Y+��bH�&�]?en��k ���YT�J�,�?q�W����ײ\޹��{���d3�s	|!ӻ.׏�K�	��)�ԍ�hE�}8ؓ�C��5�H��_Ӗ����bU $Y����(H��*� ���Dc�x����D^����o�U���蘙���5�nќ�Dˆ���I0��I0�k�ʊ�.��^���O%��_�����^��rBr�8�d& ��Y
�94�,�o�u�����'T�B*V��U� �� ����aCH��<���ҍyRD짪hH�a����xuкx��\* /.^u`� 4$��lk�T&_�b�$�
=�s�e�S�vT�X{�5c٭	�h���"���~zz��ءx�i�%|i���Yj#v]�)75�<��ƍ�� ��NX��.:��yV���Y(F�M���"�j��5�}d~��k�wa�TҚ�GM� 1F(1&V���̸�j�hD� @=*��ܕ��C�k��J�t���VA�Vam��K��,�n�o�*˅1��'G|�d�+���5s�ķ�����d��ͭ{-,�����5�tf�S�SP �>D̰_��x��������.G��ȍ�vհ��r4��zۺg�����i�g��%?'s�i��C�p��͓r鞘���Kj�q�p�o\��n�$�l��7��\i��/�ROX���`�m��zu-��ǽ����;���C7�Wr�w~����ெ����Ŝ������Q��`Ř��5?\7HC���sѡ�o+Ƶ!b<+�ʢ�?�<�b ��Fc</)���IV�A���C<��?z8YLӊK�k\�Ál�?bRd�<~���Cuޏg�ت!I��*)s�I������v~q./�?�w�~��@{�!�t��8�$��=�!���X��������}vz���>�X^]����kV$��@���­k��lU±K�`�@�uRU����q��`<�Z���;y��[V�Hü�Q��:�x1��V�����<��!G.���}���#�7���y�e�ZD��ݍ|���Ǐt��:����.]|E<���?���OҾ�7�o}�[�����z�o}�[����6�6 #�ч��fRT��f,L4��_������>���hb�����L�Q6��"!M������+�9����� �:�w-ݦn�XJE qIo���L2 �i��j���m��%:4���2ucnBGو��Ay��h�eN�F(S2�e;f06�� ��M$>��m����r~�B>����`i��|�\ @dƢ��";�Apw��h����^K=T����u#��OƔ$AV.�y�o��lR�xd�qǄn�b�ljhK� ���P��2�N	�uf�I��vd5�2%=v�����Q���:�yzπ��Uz.��G^��m��A}n��7��+��:Oo>K0"�Tp�I�a ���j�x/	��4p�`sF����=&Ȉ�E��
؛��'B��eQ ��j�θ���x�ͿaW�����9�[��pk�^�$��U\��(Sa ]TE�Id��;^��$^36�8|&�{��x�����u��"��Z%��So�.1�T�P/?2����{��R��,#;5�s5w��yf���jR;1u�S�W�%�/��� aA�d� 71���s^0)�� %m���rU� VG�D4���4�)w���/�jV-��R�~Vd L�l�����cC�' �(���.�An�� Jb�떫Zn�3��RV�R./\Lt���za yľ�7PرV� ������J}�HN�9C\ 屢� }A���F�I}y���
	r�~N���j�P�Q �a<����(�pWd��b92}k����w[г`D3��*J��$� @��̇�!�Ϊ6�-�S��	�6��m��+�y�w	1�s�]?����MO�3u?6���/��Z�}B	3���j��Ȭ�H�3S^�+R�e�h 6[v�s�B�?@0�F$�?�ܘ� �����a(]l��ѐ�R�*C�t{�jC��q�ts���� �
�6C�Ak�@�q^1N�n,�Y�1���U*)+�<x�l�=$��X��ר�J�9������*���&I&�(u��O��
yO1N����ܽA����į׾���R��ZV��{	R�DE�'���1�TZ+z�T��>���ѹ&2���X�]J2�-���W�`��U)�uK��#-��J@��%�:���)���c��� �q
�F}�Gذ��砑�����{/RB�b�ɯ�6�R�s�!9�����m�2D?B:	�q06��F�2�����V��&�Or�(*ڐ��$
x��Gc3�˘s�����of`�9M�Ýy��`@�H�;8��n�(��vQ���Ҋ�5�Je5��0��sP[��h[a��(�Ub�V1+Y�nu�V�@��QG��JBo9�E�H_�g[���=ϥ ;�xC�
��_����b�;��#�y\/U&�	N@v���!�ɁL��$��<~�j��WW$Sj���ET!����3a��V�*楇���;�s�ȝ��ݵ�VV�y��!�P%Ap��F*X}s8r�x><�Jٖ��U�x6��Ps��1�P��;�iG�!����7d�#�׷���o}��i=ҷ���o}�B[Ci��m�
��O~�6��u_��2����ȃ7�pw���&�4ē$�j�X��<&�Uxq%/�?���Kf{��P��W!����@ܫ�kn�����j(��rn�ܦ**T�'����Δ zQ�x
�L�=#(M���@� �#���o:҈Y������������|����@�rD��fy�>#u�=J��҃>6�Yո>L��<��Mw:T�������b�,Od�G�lWP�0V(�gȼ0��d1_01"�!�^.y����HA�F��!�v��Yhkf������⛚��HVz�a���7。�W �������� �:�;
<l��	��`fF]�:�ϔ� @��N��D���u�2*k �Фf��3�7��^_,`���3/��׼�����N��U"�D�����K�5 u�4逋]��N����K� �u��.~c&�5��s3oH�y�,� � �L��.��L.�-J9�����|�>�k�����$�^�\��`�f�Z����_�G-�>�-3��Z���X��Π�3HVZ i!"�D��XT�_O�w}�v� �U���(i��0���j��	A�2����cőe''�ϐ�CV:�}���^�	)�ȐG�*w��}�����t-7����ɛ���/��6+���R�+����Ci����$6�;���B�A�8��M]�Q���/J���Ι�8B閲d����<=M��)Q���^�9CO���Uӟ� !�H��X�"�sS��|�>�]�ǘ��u��;j �C����z]�;cuT�$�![1T� C_���3'QoxK���X.�xם���E��A�8ְ������xh�R���a�j�H�e'�� � ɼyvG,��*S1Aw/�W�� UG����\�{��VA�xL3c�u���@��f1	 � Җ��Y2=ؓ�d�q	`2k$TY����t���E ��>C��q	:9<A%~H�Z��X���S����P�3��V�Y�;6���}�"�* �Q���e�v}���j�(tk;*�HP��p�)J<?������s�*��P�?f*�)����� 5�O�} *w��c���,^�'��8��?�Ԍ�%��8���4�l�H�
��ra���u`m+��Y��;>9a�]���T���<�;rG�.��FV��QTZǬ�q���*-��P�3G(q��y^S�)4����v1冾j�߻٭����G�� T",GUA���'��1R(����I�z��^gq�v;\S��J��� b)��W]��ܒ�4��L�i������$��;M%�*���8m��⼎S���7��Ysxt�u���V�>}!���X��q�e�F�<(�sHH~�r��*�9׈��A"� �D?����=OƜg*���ƣ	�������CV}�|~.�����\W�2�d��3�(�$��?1�U�Wo���|��w�q	,<�c�[F*�
���߿ϊ����X�u��썆���9;����{��?��?�<�X�޷���o}��o=ҷ���o}���rq��F���U���>���l��ԃ7��7t�QH�6y؜���Eq3�e���|0ݓ�W�?�>�@�˕d�4 �6t�����E���r�^{%�������NJ�@	��5P%@��3�5�2�)��ֵi��D5P �un�@�����=bh�G		�l0Ѭ��^��᱂�-��3nX_�|&O�n�/����g��Y�1 p��&���I`���Zw����Dd�
���$m���|//��̋��� U����ͷH����d9/�f]Ⱦ�C;��A� ЄM-�[XU�|��sM�3�{�߮*h���5�8����!W� ]��9wզC���Q�Ra�cRT� (��"�b y��ll��y� ��nJ8�j2Q�ݍXVx�BɆ�����y3�����&=���<��l��+C|Ň�ڇ!�K�K�z�:R�j�財��.�|�m���5�`O��<5#?�yz��6���a��ԯDI���2��̍I��k�� '����	�=�(bU2��{��\�9�k2靀��I��"&��	΂Y��fg�A�L~Hܔ�	B3�E�g���ρz��J����#�e�iz@`��AS�|-�\�B�뜨:<p$TO�x�VsY,sVp`.3��*fJ�Q9�M�@XD�]C�@/�χ�=�y�X�Y���G�K���T�� ��z�Ϟ=a����Wr^T��AE wz��±@:h�OH4y �$��}�j ���v��?�99�X��	�G��x��T�A���:D�Q�@�C�����nB��G!��rc$02�	���	�%Up}�X��`Vȭ�wOPMi����H�c���q��oJ(zQ,�yMZ}�aՋ�DHYq�}[�?�����fQ!��ǋ�gɏ�������
%f����8��VtP*���
��UT@�Jc��Q�t�@k�-�Uׅ�q�n����y�e�6��*6�q��>�R��.#��hܞј��|�ʾ���s���:�%��>���}��)�/J��*��
�0ƤZ��y3UuK�{��9Wp�F�+ Y��r�����xQ�Ř���� �X���*�UM"�|tx"{�}�i����\��>������L���I������D�z����l��yu ��Lڰ%��+H�y��bp�%LY"4��*+�%i5�VI�B������QݔUd��:'��+�3GE�<�øw���,ݘ���~������d���F�4ЪF]�����՝��s<?��39#
�|{�Q�+���������Fxl�T>s �SZ�/�c�*@��b2�*����x�E�˅�����ݽ���*(������8� �Ɂ���������A Y�;�V7���w�&ٓ��=�_=
bU��W�	~��F������|��QɃ
�!e�P�je�{��dT�܋*ށ�g{����o�����/�7��{!�ڲjٍ@H�a�ܑ�C"$�� �(�L��h���	�_[�[��ַ��.�� �[��ַ�}a�������r-�>}*�����q_~���._�ʗ����mv�r;[ȳg�h4�rY^c 6~��[n6_�x��\�=y"U^3���䣔��Q°kl:��qsu#S#
��&�Ǧ��rj}�n�7��X�R�̖`vi�Y��@)�=w��G�z�$�R�d�b�wtt$I�Q^	���Xhd���~(�<z$��Ăؠ)n�����،��|"7�xmm� W`H�RV�=Pn>_���="�S�q��|3�яsQ��3�BF��rv�_�i�XM:��ww3�`��F�J� �Kh*<�Y`#� ��~hѸS�@�-B����-AXV����::jꞛd�7!���㥢�iW�X�j��Q��5P�U#j2F��5
ή֔9	��H���٦^�j%+��V�����ש�w�cF�5{�kQu�+A�ς� A��e)��`N`�IɌb�^��k�I�<��Q�I�3@%���%h�U��@�fCG�DGfz]+�QUjt��.%A64�Y���x@#����ٱ*quxx��|>p/�
&b�)Hd� /�Tn�kH�U�m\<A�N]5-�EA�
-z�8/� �����7�?�%ӊ�cD��덬3zVbDd(�l�U��J��p�H7jL�d�� ���K�/Wn����2Od���� �H,��7e��N�u�,�125F5���	��ꩻ{Ŭ{7��V�� �N��ŔƷ�{H�$@8ڕ;�	$�b�d���_�n"�7KCVkэ���7^'*m69�:Tvk��/G�ޮW�\]_�t'�H�� �=����(ϵZ	ݞ�����0c�Tr��afF�n��7F
��e��*�L_�\�V�+ �b2�Jm���M�2ܩ�x͞�D��wm�hUPؼf���S9(tΞ[S�I7�*�'�R"�,iF��
R��7^f��Cd�g���d�(��#�����/��O��>ʅ�M�UJ��A�1	�5<���5TH��-�}K>�x�0�͛��m����8�Q����TC��b1c5#$6�4�I����k���*'�k#�ٚ�s����A��L�d����U�aU+`(i�~O���Wmw��Z+%�mEiˮH ^X�D��������)��Y�Լ`Z<�2��8H=r�3�N���G�2f���3y�ƛ��M�����+7�HT� QM.� I:P��R=obV�)��jK�AKB�A�%<� �I�}�U����u�-�糧Ϟ�����0�Sʓ� CJh6���		�]�똿7�х {�lm��Z�Hp�� ���=�hL� ��}��VQ������!.�\�%�����X!�")��/vq�U�5�!����G�)W��HT͐HQ����C7�\�	�*H�a�Ab,���G𼣤+<p�#}ޞ���3ٟ��M_�CE ��Ճ���[+�n-fw���!��CJ^-\�ެ.��G�*�]܁��fS�zc77Q��+��|O�|�m�?<����N1@�D�z�����RgH�AJ�kh�gn0�c7��ַ���o���'@�ַ���o��dL^�x)��<��o�����r~�-y�wH$���׿�����?�@$� � ���a6���r�Ag��6nrA:x�la�<t5�:��������A�t��i���@C�6�ө�`�v �	n�%���"%Cj�?�TǙ �n(�a7u��'�?�_�����W���̀#�jV�j�G�]Ei�vk�+ZB �af�ʊ����@�lq��2Nu���ǡ�s#���Xl%�C�)���ZJ��n��U��	� �ި|Dkf� q2zf$܀��x!�Q��0�����W ��MoV�Q���(�U�\�%M*؂Vl�i�Hhr 1M��b�@�O����Q�:�4�6�x%�R	ُ�sȽ��#"���J�݊T���/5��ͷrN�� ��k�����ǘ��1>;ٓ��dP<�%\|�3�ﳮ=�K��t�)�܉��) �`��祯�Ќ�P�3��-78�gzR$�� �hm�z!��ß���v��Tnh$��\A�%NP!��^�(�J۱J
���͗A8�����w 
S�<,�6r�7jz^��Gh�;�����n1	3��uX�9�*����14C�R 
�$��# ��"�"���є� 6�: "�@��	�Vx��%.�E���/���\�BZhcRs�\%��k��� %@�M���MA�	&� �Ѡ?����C,O�k�H���b�p
 ���ѡ,ҍ��o��*$mRL1�������n�Y��fQC>f�j�C�Qr)7�#b��:��)��ޓ�*��� ��~��� ½j4�`l�]%��۱�#jo��ЩIX�U�* ��~@�7Z��	xz���b$��
T>IW9DrU���!����r���g��HJeJb�̄����Ű��2�l���A�1����H+/6a�~�3w��ƂL�,^2P�Jz�BKz3
��V7[�#ۼ��'��rsX�R3Z�8ݲ/!rc��Kxe�VG`�o�.^�Dc7�y���c�RF�td����k?{�6�G����b�X��p���$][�k���_h�f�3�5J
FV	�u?s�d�7��*<�0c<�ݭd9�y�.�$�p<��D+\��P5�O�R���C9:>���#w��j� �j�u��)�3~��Kl�1X4V�h�G$!W(�r`����1	�ED���ϔ�JX�իs�/�����x�i�ƈsT�1=�_+�x"y�
/Oc#�!�������{-��9ؚ��鶪c��LH������v�v�;iLK�?|���-$lÈUg�F?6A§ɐ��O>�����ÇC>_��ߌ��T�y| ��1�D�E<c�~���Z�G���\�|`vsci<P�;�q�
�G��/�9��k\�rkg�7͟$���Ӎ���3�z�����_����˷���\��C�@2�{�xGB���3i�}���:�jB�(x)Ӗ�6�[�����_������ҷ���o}��j=ҷ���o}�G�(ɳZP� ���Y����o>v��ϗ��~-/_��׭�a(1��UFe�:㔓�&6di �g����z��J��dQ�)���n&7��$��b.���NG6�nn�LZ��D�!<G*�#��0e%H�z�ȤT�7Q-�Z����,�;�Rn���T�+����?��<~��U~��<���%0@H@SМ�%j0� >=>p�A�}]�2�93�V�J�� ��+a�;җA6 �%��M����H�ÃC���0)�.���%l���%�JQ�Pu��MI��U>*��RT���^� ��h[�~�����2�Џc�n����Һ3:W�ƲP�NQz@`<0��ɰ3H���Y��Ss�]�q� �&˓3�\ɴ�@�* ��ߒ+��`W�	�.��z�p�LZ׎G�6�4��4R$ 1�QQ�޷�<�cWVK���_�7�}���lLP�o��)sn3��k .E�;��}�t�����13N}x�K��8�λ
O��LT|�2oH�p��1d!��m�.�n^�;�n�`L"�Q�ïA0C�W�(8���8��Y�aM�B�0�-s��DM�y]
|���lс����k�m��֌�������s�T�Z�ā������`"��N���M�gY''s7������u���~&o><�gϞ��-̱W�8X1��H� V���M�O��t�k��|M�)��`N����?8'����2��g���XAR�u�ZSHձ2C�Z �J�5��a��0�2��Ay�TT��
���U&��Q/� Q/!��U���oȴ�����X�n��� ��#�(	k�,z \����cJI$���	��n���a��DZc�#�� 2f�����!-h��� X� �з}.T���f&w7�ϭ��a���*�u�%�5��	��H�����D��Dl�_Y���zw�|�����Mpޕ����K�G���0�OĢ�0�c<q����FUV�E��S�������r'��W�jzD�4Q�e��&��� ǽ����m���_Qt�'��7$�[��J"
�;�2��RM�r	bV����)�����u˴O5+?sc����^4�'Q�{S���7��}�A�q�+9�k�LNh�?�p��3b��9d���Ʀ�}� 3��!��n����W�Gݥ�]��6����\Qߊe'+��)�rnZ};�l'�clG��(y� �UZ]Xғ(��#�<�>�U��ׅ���\��q�mW�>O��ɞ���)���WxT:��o)�ߝ�m��w*�g�eQd��6+���+�>/FVMY�5M̓��b�i�4�i7�Q��D�8S�/eY�<v���ƣ��x�~�1�Qu��I2%����	|��3-**A����!C7��H����F>��c�B��/�T|.����5GTä��{��|E���oʽ�{2[,Ԍ}��k����a�t�{��9ޛ����$���}w�#�IH��;��?�/��Ԯo��������o}��ow�	����o}��ڰY�ˊ��zőJ��D%)W)���K9=�G�*_�d�F�����P�Q��٨,P �!I0p�3d����T�y��t�d�|>�w|�k^_�PjSn�1>�� ݭ{HdqGɒ��/���� B�0Md��f�E�"C"�:���FD�(���|?�L~��ȯ>|߽~�6���iB�RE!./]�؁��n�U�uj�ۘD��Rހ��.`��o��ez�-H�o׷{{��o(����W�GЏ��
�K� 鉪������J��x|�->:�z���Z5m��Q��x�f���� M�?<�YtB�Hl�Hb�f���3���;��V�H�`uf}�Ɲ;GJVa[�4�Nr������I�l+0n|��' X��*��RA( ٞ ���	�oWw~����z}p�KH�f�3;w�fK��zb ��Ŵ
0a7��߇�9?gdY�j�^��hY�	��VMuT	 ��g�zo��3ü��lm8��3�z�.Y�;1ocJ����4S^�U4��(�$�V�(�"$ m���Wc�p ��LM	����)i��%�����Y��k��i��j�=6X���Z^��P�*�N��c��p4��9!0f��ˣéL'99>���}ٟ�	h����h��n9��<��@'�k$gv_��P>}�\�>}&��Fp��jM��0�N�� ����P3�����BAe=vm�/��IUƯ�j5ȟ |����W�� �Ч0�FU���BkH+!ۛR��af��'CU  G�L3����hLRɃ�$b�ws�|F·����X� �Q��bU�d�V���HՂ�
B �c OA���VQ)��!��v�`�bQ�(�2��곂�	��Y�R���蛵�ӣc��t�@c�p��q|:и�*���@l]��Z������}�4n&�f�/*j y��i2��Vl�^�u�_ʦ�VZd*/�9:��'��/��9��ʛoc~O�)}(Mi�Õl��Tst�����A�1�[�$��Fd�8�O���L�Jr)Y��	��Ϻ&��]_X��X�J�a���]�P�p�Q��WT�Y�e�*���Eu$���^��n9rs���ت�Ī[jJ����e5-�tR'��c�CJ�H�K�k��Tf:��L��	���x߳�����*K]��S����(TG6��k+�捃YQ�}�ԘK�_v�[�K�ƽz�Ԝ�<�P�s��W$��x�Ƒ0���e��6�$�8�B_��ugm�sV��	O	wJ>�iL��{�V`���� y��R����6�*MX���ie��q�JN�f�ӣi,��C�4]�#�bϝI���ń�}��p�7�Q}9�wV�v�x枘�V�kh�*#'��?{n-�'�\<�#~��_��¼P��F甒,%+�A��^�ч����=˾ ^R�T�KcGw���x��X��ãc�KT+q)`�p��?y�H>���r��1�
�.��i;����J������x���hO"��������a��<��o}�[�~�[O���o}�[߾����t��1=*�$��|.�7�Q3���m�?�T3*|�̗� 0d��	L���m���`�)���[���1n�52E	^���� _��Wi����˗/	�@�ihƮ�,!(
CbT]�b��
���6�n�H@)�U;�ifk�$�@	�Je42��M��ǟȏ~�z\_^1Y #�
��$ @4x`Ee�TB��5 �@%-X%�*�AA�L�� H�(7>��2�k3,%� (;rf�C����J..�)���T`�G{CI�;|dOC� ����������a6W���J̨�.K��O��_�zZ�L�.��W��A���x�u�!����ޣ�����{1��a�}���+� ��
d��H����7�k +Rz6(A�I ��#Cy�� {O����#M��d (��lA��$��	"�ӓ �?����+o����/���v���㼕�R0�n3�V���be`�Iń��Ɋ�(%��lW�K��>��������g##U+��#��2���r6�Œ�kI¤ÎX¹L�
q*�W��"�����Ʊ># �
c+4Y�1�=`�]��I�Ea�����`2���\<C6> �����;_��s. �B�9 s�W�%9=4�u|49����G�?y�� �x�����`I[J�2F$�f7�*/�i��񙁀U[ �N���K_~C^]|U>~�|��#���4{��C�ó*XU��^ã
⭇�Q�	���(�		���
$��x�5L{�c,����qLY���� �_�<g<cL�R7M��*3���g �Ab�ͫ��ן ����(�0b�f�8��l�dq��¡V"��*�T�[I�L�޺�=v�ƕ�� �]/��b\'�r=��8wO�)��D6@˅[����x��ù��1�f �q �k�,�ro�ɔ�z��Ǻ[�_[��O��AT�k�ϊ�iM��%�X̄	��*HRP
̭+ai`��(�n��H����w���I �{�2���H��Z�J�z;�R&쪚��bk��k��1&/�Q��U5�����x�B\H�)��I(�G�8�	UxT@�����a ]�ޏ�z�	�m��.5I/8�H�L�,SC��@����Xٚ_�:��*��(��Cy�����-�&m���Ǔ�4=��]��a�j�*�$�Q9<Ĩ�j-� 2�ѩ%/��Ǌت�XU���Ua��Cu�Z��.��ػ>\���x���!蚁�E+���� �fO�	�x$@�<=9�3��eJ��{J+J@��WVmf���/�` ��p��Y�����$!+��Au(ϓF��RrJ�$����}`r��J���h�I|J2@�?,�.2Qc}c��Ğ������2}ZB���{{{�{ߎ+��a�� �g��oe��.�K�H���x�$�������jJ<��ܽE�E*ǻ[�RxC���
&l����\�򽿤_��ɡ��̯od�����m\����'�������'b�'1^���擏�'?����?�O�<���c�r�����<w"9����y�k+�Z��[�*&%��o}�[�~7ZO���o}�[��Q4ḩe�Md5n���92�Lǚ��-l�7n�T�U" �CT�r���Lr�!�wV�o����ov�$ �@Y��Hmj�'d���֬6�� ���cnȰiÆ0�bf�Lm�Σ���Y��8�lyQ��K���L��s����ߗ��7�����?��O�6��|�\��JSw��=�s`+�� �ǃN��,�D݁� � �r�jӅ�J1�R=1@F�4����32ݸ#��Y�O��2�H3�sG߁Y��:�,_j�7*����GɒX����z��,#���șp����K��ӣ��?��Ȥ/�K��8Ѭ�x�40�o�n�`�5��M�9�khZ�Rٸ@õx��53��NJ�g�������z�'��
��a�h�{<�+�̈́=��U�I�%c�Ϟ����P�bk��K�����I�'K:����Vc�A���ᐅ¹�W ���ͤ�m:���ր��8��N��W��<��	IL��@yT	�� �Ȝ�)��t�Q�HBf����3@B.��=v�BV�	��Sƙ]�[� ��Hk�`���T�ܻ��v�?�� ���"*-*�?�w{�1���ݭ䋅�]L!鱯 {cf�V���PZ�Ra�L��S!�0�QWVL'C���z.��e�6��8�U�	d-*9������z�P��`�D���hܑ��^���� �@t�1��43��9	Ű�0���+*P��L�`�x{.N&L���xyAߔ��c�H�_��&��8�l=4������Ul�}0��.�Jp�\�R%n b&�U���U\e
�����)	���a���L�2Ī�B����<hy�CT`�֍�a4K��cT�Ћ��N�noH ���v�]����U�yzsw\6�
�]yE���~�xJv*�P��%~p�)e}�s��oI�,���3�� �g1hWb�W��8����HMҧ��L���k����*���G�n����S�;���'��.�������-I�ϳ����]O"�0RPrO%F���g��U� �A�b���(���'�}M����Y�YՌ�+D�gI�j+�VЈUr�x9�����$�d'��
��u6)C���3�oT=m@H��V�'>� �@ҮRƊ<:��'����
�IS��D����Vu�2��d��͵J���S��dVv�Zeۺ���7�1D��#�����Ph���ʩ!L(�����Z��X����99+��/�;/I[5��k5� zsZ uDZU4$V��RUʓ��)�-l�@��L&6\�*����l3�YP;�b	�y"c*�<�}>�܂���Ze���X-�Yj�>$��g$<�=�\�{�=����\^^��G�(D��`<4�?o$��J��{<_�MկJ���wf�^�����駟��fƾ+�\��#N#Ơ⋞[n��\_h��[S�߇س\�|_���Z�ҷ���o}��h=ҷ���o}���ά�]��@�6bȞ��0Myu%����F����0��9)6����)51 +[��хY%w�B�2o�!F��6~ I����ͦ����zyq.� !``6_r���ރ��T��$|%� #�,U��%�&�L B��8hx�,w��dP�M�ӧO����o����!�L �h�4�� ������U*E35�0�D��Z54� �,
34'�e��-QPSѢ4b��C+���r���q4L����sI�aRt�J�$x���Y�P��G��Y \s�+&@��|a��x5@JAQ 5� �{=ű�8��LM�d�������;"d<�0]9=�f��	T�	}���
�@kͿ�6�@e!�ɕI=AJ�0�wয^�ۛ��-���FV��yw|o~�k�{lJm��y�t�D�ڪQ諩Q� �J�P�*SSU�:�uG��J� T' �%b*�#`�����ɻ,�Y�- Z sp,̷�r�z�$2~&���y�@cD�F��k�~�>.Hf HF3�Av��q�!�Os]J�Q��1UCQ��m�1�D�I��![�]��C�8Jl%τ�m�^3� �~�!{�ɎQ��ͻ�3@��|��{/*�����ó�2�������M��ޗ to#V�P
�>QW�sz�Gr�?��١�ͮ����F5R2:���1pͯ�/\̼bf5�R}�li���:�� �yr6��-��[w��i!=srrL����p�R��� �<_�{|N�eZO9��%��X`e�ϸ�� �Y����V��f�\5*��^�g�Vs?��ts��|�h�xD��V�J���}gAz�%9�Z�8W"�Ķ��e[�dT�����fT���ℬ�S3{f��@�t����G_�]4D6��%�oij��3*�I���`9??��x_lX-Q1�#*�!�5�����-�.Ә�WF�r��76�D��Æ�3B�8����l���O���Nݽq S�\%�FZ��E@�8��|��Pe�Xa�D76p�M��+	ц�r�߰( �C��0� ~�nQ.ϭMia�M�FV�X<EB�\�MI` �`>a��y q	_�՜��(8��{������+���ѡ��Vxd���=Ƭ���T�[�)�~K�!>n�o@���3�/Q�{Zה���ӡG	�x��QZT�H�*[��q���ڪ/����1�
�&ꈒm��$��>�#T�,Ga^Q�������J<4����A�Jrbl#nSB��/���z����<��'Jd6�� dּ1d�T�����WM���C���m��,1?O�#f��*l"�0�RF�A��P^#@��č;�:����A�y��Fn������n��g��A�	=�L+�����5�0�j-̝��� ��9����TN�ڃ��x�B>y�H~��ʏ~�C��O&�n�Ҋ <������[�i;�VJ���j��=k�q����g��ѓ�2w�T!�
��Dv���=�#C��_�����sV�?x��jm�r1f�*�����o}�[���[�z�o}�[����6d��ڣ�c�淿#�n�6[�������~,�7�ь&S�(X��A���ҁ!�2��a�"Ȋ�d�����K�|u%t�݆k<u�
�]�x�v\*7 ���\��fc�qh�La P���}y���~0����J��f���&VU��X���f~�����'��T���A>��c9uN	���#�)�B��,)u��0	Tm3Scf ��Fu��@%d��*��1�%q���\JWA0�dF�Z� >�jM醒2��k�D�6����1u�D��(���>�@-�YB �gG7���Y�� �{ 23UQtקV��-b vn�N:j]��E�Q���l�g�0���j��n��nf�vM?��`�
��z`�]��v�{_� pYߪU��gd>����JeW��g@�ʌn>A�	?�=����#v=>|5^볉�T�K�O�t��i�v���D��V�v�f������Z��`4{O������ �������7*�x�l��T6㯲�$�lK�Rk�H���jFwH��twj�+Q6�Y����{_g�f�b~��n���<�o��W��xՊ�،E�2����N�Q��۫k�1ʬ�_��˙�S�k!Ý����B 2���1Z�� 2�)iP��% � SaT{�O��Ŏ�D����N���fC�/���	8��������$j2T%�9��ō�&&8UѧhC��╻K^/*8�P}NNNF� �#�����qV=rrf 49V���nn�H>�kY�x��y�
����I�%du��m���@Z( @Q�D���@��N��xe�; ^A� p�R�*_87-�����$��I�����?�,�'���;��T�o��F���#�'���q�����$�nn�\�P�����9%SPU����� A^R�-G�ĺ�?$���8���*6��c��-�\��
&��� ܀D���
�*j�p,7<��� ���h��UL����+Ə�H�]C~ѝ��<>�#����ೲl��w����d�U8��(x���!|ߦ|�� �w���!��CME�o:�1|��ָ�E&���9��7��������k_{Ӎ�9�	1K7����	c�H�,!
����0e�&֗�I�<XQ�0� <�kv7������0�a����0����/n,�x}'�W^6N,���X���G�QȵWT�Iu�v�?<Q��,���8�����u��,�9��&29��}G�X�-�F�"^?��n��0�"��V��4�X@��y$��}C]�@�"�Ԟi�Z�Us�����̓�*^��
���Fj#��}�h��kFeۏU���٫�&���e}˟��p��D�SHB��9wtxL�(�� ���=]��35M���ڸ��S�^�B���������ϯ�GCE*=V�5?W�MB�L}��Ϭ��ǈ��_!�Vi�{�36b'���5$̌Bl	R7�cխD��\g�����yU��a����/���?�W�)�c�ַ���o���'@�ַ���o_X;<<�j��mʱ�lY��{���|��o���|������?��e�.d�)I(�̈s�Ph������Pb�������|Ib���X�����;_�f�W?�����J��ԈNÌ���򂛮�U�>E����Kn�j���-����\_�M9.d����&nSyh� w���t�L7�^�Z�J�//��>���g���!�=�'�������}s�Q�(���D� t(@m�k� �f5o�p��U�� ���o��
�=�k3F��YqIFC��(A�R�ؽAp��/����}[�YΘA��P�ȣ*D�C	$Gu�`Vh2KХ�x��Ɣ�G��`˚&����?���>�����YB��ؚ��=Mˤ�f%{)Bf����~l(D�Q���d���G���`��U��A�5��|B��MsgEZ�G���� ��v��mo��?k���������5�ƟoК�Vt�ʪQ�G�F�&$��U4B�M����0�����u�1�<*LrC+0<q��Zq�5M���g
*q�!��x�e�m3���*oGt
� Vy����-���u��kS͌�H��i�$lM��#n[�g�д6�G��~�R�&91oiJ� ���Wsy�+I镳7Ƚ�#9;|(�$��%��wY��9w1���}z�)&����_�+˘3�{�Z2����y[iEK4$@.�A���B��k�/�H�}w�9�hT�%*�"��n,[Xk7�,#ͬ�/��e4�2h>�q���o���͊s�Ƚ{ǔ��X 	}�ީ���Sv~ �n�o�!q��&���*��b|�����TJG�|4�MiI��`����5�$��l$� �̯VK�y51kY�j���Ӫ��B?��U)��U+�@�t^���6L�I�~D���ވ}��}&��X>y򉜿z���c�n�3&	;�g�h�RhX�JV�2_�̬���QQ�&(J#)Տ �����r:~�q�5���ɍ�OHx+�4���aoZ��^���� j���&(�/C]�E%��S���F!��H�h1�p�T��W]![}�X3��a��u�Z�hK���i'6z��n�����L�8[�j=s���	Ȍ���F.^�jN�J�����O�����{rp0�WO]�)��ų�*�`i[��ʋb�9:<q_�g�� Y�/����i���/���xo��5���-t�{%��*ӄJ��H ����F���[[	JH�IToID���`����߱yi�$3Q���1"1����︿j��&xOc�x~��R��n�\���c:Q�
	$x΃4�r9c̎����*��Mbd�`�q��V�K�f]�w��3,��r#	�*LI̊'<$���M�dk����QW	�7{�娤|u�>^M%nb>ێ@�A��g����01`^Y.�`�+#���X���l~+/�?�G�>���[�H\X�,Y�ݻ4𙱅�;��r7?6��R�ڠR).����!��=7!�歇oʷ���<}���x���J �9[M@X�%ɚ}7�����eE/��sĮ�k���K��ַ����H��ַ���m�I�ߓo�;r��rx�<���#�r��m�V�����c&Z�~~y���8���θ1B��˗/X���o|]��?�S�ַ�� 6����}���䡝E=��<b���P�i�~��   )��3d���`p��%���^]��޾����χ��hd�!-�1#�`Y��\__�������F�<yB9l^��w�N4��M%C���ϞPyE��j�¯�,wl��c5F&��H�,����a/�D����F�B�N���f���h��/C^V�0��d`������Y�Q�ݦ�ԩ_���@��o	��Z���A��H5�ٵ����DL��nNC^�=�P�����D��l~��,���b-
�C��^�8��ѲU_ �D��c�����jT�j�K� ~��K�[�04��A!�f�- � �z�<�9U�z6,�ߪ7|E����?���"�\�����s��f���f�̀��;��rÁ�|D�2-���- HP�6�A�[��c�'��A٩����r���X�� ��&Q"#M�*���w�V��"�G^ӿ?�?r�kT�	D����JX��A� �b��J��:�F3XCp��O��T�6f�[�@h��^��Q����l��Qm11 a����73s����g�dQ�2%	�i>�iE-��
�2ח+��f�"c�tc@u�1S��;MG6M*fv����	�rݹ��9��h�w�g�lG��DFd�LD=]�D�ڙ�n���u�>f0�,��A�
.�F�˂�+��� ;�k���� �Ļ�!2	��R8��0M��A��y��ҵ�8m,���dxa��� 	-n���P�RV������SB3c�*����	�e�P	�r�t�\Jii刂��ŏ�J�{�P�����Ige$p����䇏s�#?xM)	��x4 �W���WkV9����VY�91�Qdb�c>v���I|ƪ
̟{ �4��'a�c�t�HsO��4����=/gWw1��D%h���V	aE�v�	�{�B�����P�v%�}5	�K�S���e[WVA���cW����!Η�\-ǎʳ|.A�(�x^�h�����n��5�?��?�?��"S�I���-�ٌrCs7�������T����H{�(u�g�.�&��M����sӊY�}�fn��\^�yR{�
��1�P
�K��*����U��I_"�OW$�ʜ�$__�� ��ے4 �6d��<�M����T��.�Vfn%,� ���$
�����D=��Lk�R�~je���qk�I]Q�k�M���� �Iam������!�G$@.��+O�x}�P��Ⱦ�-f�JbE4�O����M��H�I�.�I��u������|+�O�W@~���Y6�8��ˍ�;�~q垉����y��\^�����|>c��+���t`�}>k�D���e��bm�AB�jI��o�z@M�Z���}K���-���D��'���|�����,�wﾼ�֗��蔿ojM �w�׿aD����Cu��ַ���o���'@�ַ���o_h;8=�o���q6dy��z)�龼���J����2O݆l$�w����%7��''n�vJi 0_�s��o?��|��������8q�O�2���qg�!c����!0i��M��bICMHd1$�9+@�	ܟ�a�d<��|�eb��5j��̋�r�6�7�7$Z(	R�4ΐ���W S#W�v �E3O)��ꆸ*U'�?�!�-TG�m�[ݕ�n���q��!H4��U�Tw���f�B�F5̅�#~�lrfԹ󩓊�; �Ѱ�O%	���ۮ: �7���IU��=L�Z�	 �6T��樱E��cI�5�;D�I~��
��0ū]��Z̛��D�8TxB�8+jn�Ĺz��Ie���f� ����t�����p�\�����-�R$P�O���8&��w���x(�j�]�s���Խ��7��,���T��ʮ��ቑς����QU�������Pߗ� ����FNI��H=с��bF���%ZX�X���Z��=xO���Nކ�^�Q�ˀU�^e�����4$9�gA
h��*:(�asJl��=#������V۝`����`���G�P��	��K��b�0��>��"�\.no%�����P�SN�8r�F� �;�҃DԊ˭�X]m`�;2Px@���J����$�*VDD�)�
�>7�A ���Ն��h�������Vխ6|�V�)0���3�^���M�]Y�������fcH�>D2�Pb�u�lq�J|�&��"Z��@F��V���Rc#އ{+�J΀�"��ͦ��ī���"N�)�V
ԕv+ԓ�&�\@�M��D-4�,�zz�T*#��XM_�6 ��1�7���Ӥ�H dd����D��'���'�)��1�狹�"����O�����9����vAhp��)6~O�2?�C<8<�oL��$<満@�����1���-%cV*}��\^��K�,Z�k�؉���j1^J�`܋$����=���^�y�;�I[��ʜ��6%y�Χɯ�o��>�c�o�U��d,#)��h�$�>徢F�g�o|�������䭷��3C]/���
��>��ސg�%�r�*�a&j/T��2K�yGh�z�����W�3�������q�)��ƈۛ+�o��X�l�2�_�Z���� ��ć��|�D}ʐ�����[����l#rq-IA����$��A�+q<,�Q?�De�`�m���� N��S�"!R�_A�㱡8�w����R��F�{�����ohCe��S��? ��*1Ҽ	����o���,�Ă�k�8��	C#mt�k]�B<��q��/dq����[�������_��|h8�tO����Ŝ�l!�.����B^�����;}>��U��*m�%��97L� �ZQ医k7w�z�|�ڑs���3m�}��Z� O�˃7ߒ/}��2��O$1@�v����E���ߔ�#7^'r�(���$��dk��ַ���w��H��ַ���k��lO���w��&��X�@
}A�o3#m2�tƹw�MΧ�<�����rswK�rx���+�~�����&��f����YV�W�Y���T�HA@��Xss�����E���B�C}��e�s�9CVdj��
�^]^���5�:$#̂"KX����4"���X��@Rf ��A�T���`u	��������Y�P@Z�_�b����� ��I?p�ña��,d�v�L�;�1<  ܋(Z�B�6���%XڪΓ���w -�e���n�߸sl�է�����H~��I�(�f���yfGC���l��N_����5n�(�X,��W�O����΀x�m������z  2c!� o	�>�~eEE��n��������(���Y��ܸ���I��f�0C�y���3�1^�U�{�w�K�x�п`�73ef��;v��� �K��$ֆ"���
 ��$�<9���j�)oaRP�!0Ȳ��0eq��[�p=�¬�v`d�j��;�i^#��VAġ���H�b��sA�c��Ě�H�M��{ 9��h(o�s���{�׹��6fB�>@,}t�jĤ�"� �U����I��ިր�_R��D	Ff��z��J�<!�����V ���d��$���9�g\?�H�dO�s �g�2���}������f�X�5 ��V〘�����a���{�p�B��  ����)��@�f	�TQ�q�x�Tl���DǱ���e�k�U��VH{�7�a�Ѭ���늄͊q�˙M&)�!�a̽���l$�..^�[o�M�hT��V�2&�@��\� ����!�2�qo��*.,>0���� .��5���q
���������5 j����T�e# �z���G�Џ�&��V�x�j��c�<�b @t��n̯�!��G�|��0Q"~�ϝL�d�`��׶Jn7V����Ҳ�O�լ�������'�������a��@����KV^�n�6��R?��B�)���Zh�ι�^�
�%��s�j�J�%%\��t�F&����u�2��Þ�F�G��4%���G٤x[e����b^��U����w�#L�pc�W�a�F|�<�D�㑻�k!Z�����K�@V���_��o���ٟ�|�\Wgw3�Y���+�����t�o>��HxTk�@�� ��]U*C�����zp��U��p�
Ym�t�fBG���!<2p��6����3�A��1� 3*Nm��2�r-f��������2���*���g.ДM�B=r'���>���ݘ�~A�P��<��ׄ��(uU%�U��9)"	F�R���*��*�B5����N��A`��S	R%�?_	�z�s�!�ߋz���J/e8l�QbR�$H�%�9���+oi_�/T�� ��V��$ժD����'�\_/�Z���ITC�����щ��\���t��t)���g7c��X��5���uQ������!�ϒD���l������O=���cw�"ӣ=VO�e�y|z"��}}�pk�װ�m�/	��ǇGn�0�k��C栋�W�N�ַ���o�{�'@�ַ���o�(��� �7JG,�/Vk� @���Jf~�I(��2C�8�jlee<t��Cn�K�Y- w)� �T;���7H[�N5���ڲy����5�� ���"�z3_�|~K�Y� "	�
$ H��܆���r��  f�<ȸ�f���QIM䅻>)BY��2���ά`���_}>R5č�k Rf%2���� U�\rJ7�( ��q��rzt�XfY/ ̸2�� �㸍t�^�IK�ٕ�ՆY����-�	� ���]�!b6cS4�"ٸ����Ii�V=C�3@Sh` ��hdL�Z�-d1�p.��C����B�1*�Ka:�4a�o��G��X��0R={���[�+�Rf��$W�n��M��Ͱ�2�����Z�0�x���\���X�4��H%7D_�	 B�(�5T� I���[3W=���Bl�-eeDG6�9Ѓ��?�[�P�қ"�lؐ@1�e�13�����H�ܚ����>����
V{l��Q-t`;���(�j�
Y�ͺ�ڒ�X��~T���g ���~�+f0��Ai٩��ဦ���ߔ�X�*' ���k軋��]Sk��Vrs����0s1 W#x;�I��%^)9p�X��˂�"$@���č	�d����$�B=V+�+#$>J))�Ҷե�V��P4;��dx�X���D!�d(�bEi�'���͵4�|_^]_�;o?��o=t�����f{�����e�({�*yE�Ĵ6`V;+�Z�B��S����Ԟ��W�qsq!*�*�"g�g��Ky1{��K�x�.�@&�DI�@d��ӡ�~h���A�D�g�UzM�: K�P��T�}��kd�{;M��� ;��6@_%�w���e��:&��C
&"�"�Ń��<�C_	�.��l�?*q��	�Q�k�������Z��Ød;�z�&U]���Kd�/# \��N���+������f�JǰbgI���h8��MHܜ_^��/������~�g4�AR�)0ւP�/��w^W�Wn��5t�1	����6$"'������W�y�ф��zw7'�	� k����� O�/7/�n�G�8b�jB��؍�!!U6 �[H�T%�,>[	bFQ�5'Nt-A���H�!�bf�Z1/O �P���W��o8GTe���j��[�J����0���k<���=�DU�τ?�o��!&�5d�Z�-rs�}5�R��}y��@�������~_+�5���ɕ�Ϳ���/*���?�w����ÄL�dF�9=��F�)ىX�sBE)� Vi�c.�:2w����d �W<�L�.�v�aN����L(�3���:��8�2��3OmZW�F�THH$��ҢC5�����#c�)}� ̒��Ӭ]�EBF���B
��\�G�[s�sIO!U�9�SV[.�yfViWSvL���Pn�kX���\�����-ɏ�G�	��������L����wĭ�X��R�U�x���h�F��"}Ր�bRV�%J��jkz�(��Wg���Tr屋Z��R�K����q�Ʀ��ۛ�ܹ>���(X�|�������·2�E��DÑV]"v�V��gd>b;�Q�ӛl�1�u8�O�u���M� Ԣ/�3��/�o��=z!�d��[$��V���"+oAN�s�0΄���A�Ȓ��]|J�����k�?���{�%[��Hl�|�̓Ý�
(���D6�6�z�L�����E�7�d��z�̺�&�1�1�H��[��x����Z+"�Ph��
��]H���s�İ�������ş�Ԧ6��M���&djS��Ԧ�ŵ���UY����_�����Y�����"��Z�
�SX� # �.��N�P	{_�&�{ ��wGVv�i!����s����rи`
�9����*,��} �T����} �%a9�X���"0C����X�yX���y\?�q�  �������� �8�f%-*`՗�b6	�
��1�R�c�Z`!-x�kN��� )�}�@�.k�5˕��J[��W�D�U"�T��Qы�0 b���E�����(��)\p*�؇��c��3VZ��'�l���@g���=� ��jNR*�mz  Mk��9�ʞؘ����0{Bm8W�螆��2�V��m��V�q��_p�e4�X�� ��IX�y�'{9���T���@�7V����8Q5�#j��Zf@E�VJ&I_E�^�C�jmYUo-���S�`!�m����}Bx9.��2h��=�wW��Jī���$@� ���i6�Wc��3��	4�Jn����j˷��������x x9KsV%�:�ꄖ}����1�J���F5s���V��^� 'cZ��')�M ���@�B8J�Z�)�,$��K�Jد��)��p^:�U�wj���5�)�i�����g�f�(�\C6� ���_���!@�\��:��~���u'��F6[�`�䜒��X]Q5 +*��3����l����,� \g����r��8�S�F[d��5G�*-��
�տ�+:9�����΅�t�y�E
T* ��?n)���U�c�i�]�Ϩ��qQ���~��C����|?�~�\$ob�*g�زv�����������<�E��U��
�l���82ՋZ����m���>���z(n��Ҭc.���
�p�O{f,A-�std=���L�P�9���|��M�'?��υ��%��,Km����:ǜWi�|�O�깾FI�$H��vu.�x�1�gPdU1��v���Z+�1�"ojq��TVz��o��[ľ�c8��X8'sf���\}��_�NJ�#t�$��Dkk�#��e����\r�< �=��S���s�P�Ý�]c�3��}IV�b�z��`�ԁ��#�5'��4�S�c
}��o~�=�����2�*�?�����'?��������������sI�ys���I�̳Ȕsa���	*8���>VG�N;ɚ�� �+�é�����g?�ak$�Y�F�9�b�f(8��fRI���M?��un��`Tk��v�����AsД�V�����D��*Ec;����dP1@�+E������v{�X�X�ܟ��
%�C���M̪���mj{�䧵S��p���(:�k�1Zȡ��� ڏ4o	��\�����`��5Eu,5�(���g��!:��� 4��hC�`w���π��=�U�e���� 
x�JhwE���N�(d�q�a��@p�j�%�%H����б��m�I=�������O~$�����|�ߐ�������Px����Cf��b����ԅ�S�ע��.�����g�&l����NmjS��Ծ4m"@�6��Mmj_x{�}K������]���?p���"ٯwr,����_b�t��@�%�E�R��?lI��av��yX,��\����g��òUnY�����;�-H�po�@�E�Bf\ �2�@,T~WX��3��f�����!,��b�(��
,W��]"��J���Q� ���s��fD�>4� ܇ݑ�ZlH<*���s��j;��	,GI@D�bU����h@�!�SQ@�g�e��],5��c Nh�i6�2�G�Il%5�PFU~�dE8�Ie�4@ี�Q�@v�X�2_�
s�^�3�͏%*���F�ڏJ�S���R�ie=�u�����-�50`��oN�B%A�s˽�z;V��:��Y/��"�>Խ�|a�0x?*+d��
��$�9m�r�W�*A�rd���ЊR�\��ā�%�5�	��2�^�d��*��	�+��.��x���7B�A!W��� �Y�A�����Ȍ��!�#1k��,[h��XkFBeD���*n3������dQ+1 �+�jg��8�fe�`@�S�&���O�����#�?n��Z�,$���Z��Qu��q2����"���
۬
��X��in���y�������w�	����Q��|&�WT��f�\��N�`(mUv�X�p̵�"�p�>���$��o�1�o �6/T��]��e��N|����J<��@`����4��2f+TIT��7��,��ub��|���{�G�HL�:�lZ�ƹ� P��E�B=���R�Un*p�x��qK��I&������y��Yo6� �:V:ZZ�\3&�������N�"�F 6�����:�#�������۷a^����ן|"��������OͨоN9�ͪZ��-���2"'���5�l���Ȝ)O��PE��%E� qx��2N`C�a�*��m�Z^�rT��9N��2Fm� ��
��y*�yY����$�� �C��	|q�Ɲ�e#��S��T�ϟeD��/ `��ٶkS��/*�'IZ�M*f#�vK�Y1�8c<��f^JxB��7���������o|�kTO4��ӿ�����}����<\�R��rVJ��+�����9#|F���\�)��&��i%@� ��II�z�_s;�����k����~/��cf����U��L����|>JX�1��c����g&@�>E�E8��+��X�,�j[��g1�E0\�(�vSj��S@W|}���c��.#ܩ�ev�)�T��٪��M"6E������!�c}~T#������|��l|?iu*U�2c�U� �A@7�Diz^ڳ��Y��|�.f�+��~���b��*L�u�Ses�Pm�Pl�H8'v�i&:��>��mx�<QuT��|�N����(��lJ��c<��I�
4�_��±i����������ų+���c%'�쀢���3�雇-�8��a'}�������|�!	�o����?���
djS��Ծ,m"@�6��Mmj_X�U;�ZC���(?��������5=��?�뿒�����y�����aUt�pO�Xo,=�YE�������	4���$���{6���-�� t4�.4)�a�V6�Uv��"RP�J_T���,��k�6��� ��X<ܲ!����&�\AT����
�)��H�P�uA�A������@��5���ǧ#���쌋~z�WM,	�I�^tAJ����D#i�����Vb�
��d�Њ*����w�`~jzP���T��ZQ�*�۴C,��h,b�_�����\�3�-��Үn`Kl�%G�Rz�aL�hU�{�eb@�z��޸�e\t
�Ű*BEs�՟�P���c%�#����X���
p�H~����EJʀ��r� %8]U���C�����;��d��8;d�E0�T؆�C�z��x@����+�\��>�N�(���XV�j�h�F�U��2�ÁL'��#�d��D�Љ��S%�J���N��n;���U����E�5�ׅ��N�'�'�0e;�L`�����G�O�&�%�`�'Z	�`B7j�}�>�ʷ���Z�%6�{*Fp��?�>P�r(�*[��]�Tr����f+�o���W/������Յ�.� �m��鶴By^d���@YW)1V��X,�e���̬h�s3���r�H���֪hv6$i���b��3�����<�q
����`ղ<[���>X��P ���L��Id��(v8��f���̛N�U��3��~�ź��{ e�z���Z%�9	
��GW���l�J��b�}$N�V%�&����=�o���|��$�����A�@|��Sy�{4~mӠ��YF�壟s�
	�7���݃[����{"�*�p͏偊�x1�eq֏yU�y��4�~%�aw+"�h�������Z��fxzgj���t{�\d_��~m�F��c.�=������依~~0��H��u���>��9]��Vx��/�!�X2�����H�����:��b�U�?�(y�+��?��?�o~��T���"s��?��|���\���o���|��mx&�}�F�}�}k���g�V��b�-�p/*5�'�y��cŐ��a������s���<>l������Qno��A�&��ۓf(H�-zH��/mߟJ��AI�!�ei?�@0�q��ZW�f'��r�h�$�����&�ه�I���J�/�f���9?��J!���5�1f�az����z�"ףV��$�q�sK��X�|:�kb�.k��H����p������U¹��
1��K�<��o������>�e�Դ0t��W��6�{AT� �.Nyl!��)3X<G��(��Jת
S�:��}ط����XI�H��s��&
����=�R��*�S�Z��'��}�������׾�>m8Aj����&�;R��z��݅u��a��½���V�~�!s�6��Mmj_�6 S��Ԧ6�/�0�|ح�?�k������'?������-�W��-z���C����\�duK�FN�9�t�wuy-�b�E����z dEX�=�z �,��kRJ�	�Ĵ8�B��z?�\d��.IN�@k����&��j�'�}N7_ �	����ʃ��2,jg�e7�
H�1Ê��Eu���������N��D�BUP�S���H���"��uUk�cD�
$}<���TZ]��b&��Q��!#DI�",��(m��.��h3��� ����礮]=`ժ�U�6j�R�j��B��Ϙ��ғT�[=XC�$@V;'��C�4C�~c����4��r�]��C�}8&���U���b���{��ۯ�IK�X���" �0Й��UC��2��nU�|1 2��&����clo��D���p�����iܡ�a�h�ev0^�W���9����(���`A��a���Њσ=@B^�Dց��~�m@G�H1���*_Za ��}S#�]J{�:��4����L��~LO�3�s��  ��IDAT�\�p5eNb)�nWD� /B�͢	c�x��[�44��'D��"����րu� m �%���n�=	gr�W���H��e�}�x@>x�Ca�������^%��r
����-�[pڗ��AEm��Z��J�c>V�f� @J�"���⒊����dxfTH�r�%��Z�3^����� �I���XI''[���a�����'J6A:�6|-�mȏꨖk�sX~�\�#�$F��Ê�F�	�����D���W笆ּ�gM{��~kVG%�Nf�e���`)�k^����o ���Jx>��##�b�L�^T�Aȹ�� ۛ��1~`At�8�}v�M{>)�q6��K%����M��U���&lw�A�Vq��N(�%@Ѹ1c�����9vn����������hO�%T"�%��@�$P#<�����Ъm�.��3ԊP%]�p���y�,�ϲ�'@�-����ht��R��m��5�H���W��ܩ�1kM%�p�\M�s26����II�� ��5+�8j1��D�a������&���ר��E�6^�}+���w�?��_����-	cE!on�ʳ���=�de,f�����B���Ph9���7�Uª��/�~)y\�q��	�+�<�X�F;s�wD�q+R�임
S�5�Bř�H�Ш]��T�}�����lS�o3{1�I������{$!c>k���7�/��C�����f�\��0����&�q��j��p5�[d������������VR��V��ż����Op�� ��l��9,�g���Y%ߋ<�g�$N#���(~_�L���w��FΩU'� WU�V��--�h�L��BX�
�!v��4V
Hq>_㿺���C����F<�B�$��r������{+����W�J�;<�><��s���yx�^�s� 9��|�8�%�>X�5����/����?���N�6��Mmj��m"@�6��Mmj�1���r{wC+���as�
5T�������a!�3��9r:�D��^ǵܼ}#?�������?��` �#����+�t0�nVv[E" ���Up��"0��KX(��lɭU��Z�s��*CU�w}})W�W��RC������T��`��� �Ċԓ�0@ ��ZA��7,8Q-��Ŭ\�/C���V�@
���B�2C�Ն
����V����7Xku�S���2@h�����)J4�^�y���Z[xG$o�z�}H �ȅ��%qՇ�y\?U����8���p��ؠ���p��D32�P� �7� V�V��c�Ap-	��"�I��a�fyk�<6��6]_
@/��h�04��z�}ī��UUD���*����}Q9(�y������� E�D�؂���	��@����  d�0�C���"�gJ칭Ve�쨡�l=���&=��j�.&��X� �n�b;KU]�y��2:�¥����c��ځ�Td�񪗿�`���zO�
��R23����r�9i�T�T��*Vًw�ڑ�(��
e�+��K�~z���Tt�*��0S���I��B@6H�2\�m���Mm�J9-��__�����r�b�Wj^��D�����E.���q�L
��/r?�5���)��66N�G�<7Mη�"p~:�݁M��X��Cs�M�9��}�<�J�К >m�"�P��vNm��H�WJ�w�l�ɏr ?�����x��;�1�^?J�+,�@���c^�Z�����,���r*2�C]��ߙ����H��
A��lN�.���w ~�p~|||�	���3S"2�Ηgr~~Ʊ�"�� �gNuE�w�]��G��	}��9�Ҋ������ᜠ���ǜ�Zn��n�.�Jת�s:@ʢАyU
`�{� �Ł�v����b�;Ҹ
����L�jN�:�Kҹ�z�X�:%�%�]�}��J������8�~�@s5���(Ϋϋ ?\��v4�\eYN�ەd���\S"D�:_�|E�����>�!\���'���|��k��&[����8���|�y*M�WҲ��H�J��s�m#ޙ��bG��[��Ta|��Q>�d�y�;���0O�,���e���^q�O�H%ᶕ�!�"����S��~@a� ��sE��$�9W�h1�	�\U3�5�K�Q,��jk+'�΁�#��Դ�#ӀΑ `��
Ȏ��#��L�c���d8��#���D>_�cs��G�R��^l����~�/x?��³T��+<l# ���(E�E�f��@5M�畹jlDy�N�ґ=7�KE�@�s���1^�}��%h06`��ߟ̮��BiM"e����jaaɮ)�C8�'i�Y�0��sn��1A-W��1[Υ�z&�� ���;ʘsRbn���o3���������m���;��Ԧ6������ ��Ԧ6���F���Q>�<ȧ���뷯)�GX+�k�gKY]�HjI>���v��EVH�X��~+��@�����۷�� F�1���X0f�L+��W�<n�E��j0-2.�QыE2���Bn�;P9��t ��0=i4�<y�|��Gd\]�����U	��VTx�����ͽ���P�k�P� <@.�-*�@p���j�6Х%�@(��a�	Z�Y�-Ɂ�] 3���w>��HՊɎ  +�	JvR5�n��� �*r��i�bW���_uk�G�<E���\۬�~䢺1��X5���b�s��@��+��c��n/\/�~jS��j���i�b`�m���@fD��j8�@�,�+����!�\I�x��8؋��'��a�GA�$Jf�XMS�$��H
���ǶOzN��u�ȫ=qƁ�M�����v1^�$�oO�%�~�)5"E�~?BM��f2�K�����}qb�$�Yf��� 4d(H������gFXvcګ �պ&�}���8F����<#��D��� ��ׄ�Tʈ;��+-Cd�m��X� ��T�0Tbgfa�+�F˙�G ��0v���Q�U�����j(�0r���}�%��B �'��JyR���������HV��(f)_P쏻^����ϡ� ��Y�/ L�܅��͍�?�+rZ�̬�u�U��n�=�1�������~�3�ףR=�\k̕J.YNg�R��Ru�P;�x��H�~U���
+�S12�Uz-�e�9���
��B�]_���_�H�*�UU]b��a'l����J\�fȁF�����g5�i�>���������^ބ���p������ ���J.//�"|A��Z��Z*��Gyx���Q�J���YK�Wr<�U�r�϶J�b�s>-�چ�q�U��=�L��3f( ��a�h�a!��5�R�bn+�9(¶�s����Ґ��T\Z�N��b��గ���f�,�Xr뿪R�׌DB�>�[�)�ٚmS֫
\�W�N0��������z��Gh =��V��;��ʈ�?���;�������!�%ha����J�/��Fp�½�O ?�L���n1���q�~�������b���B�!/_�ùu "��V����$,��|�Y�=�@,z����m��|5��Dr��L�O�/��t�L�P�=H�y��jMjV�v��`��/��;�y�RKS�bl�@��JG������qR��)�����3�|���K�d8|-����<�"S(ꣁ��T�T���5\�vN���,e�f^LI��7��E�Ke?���FL�1��ap<adQ����|/-�bIC��H��i�L)�����:���C�G�Wy ���k5��=���9��L ���� �ʐ,}rΘ��w�ɛ�U
�p'��Б�p_�o<��X-,+#�O�0�;�k�����}��������MmjS�ڗ�M�Ԧ6��M�7��.ι@Y�7�~����8[��Ҫz � �࣎�r@�J�e	�� F�;� �ZT�f�qD�l!)�xA*X�wbA睩0hF��X3<������Յ����U�j}�X͵��a�?���^6�{A�z�A� �a��B�q�f�/*�@��<(�s~\E���[+�g�c�
ے��,��]'�z�$9+h�◕�U�.��<�}�.Y�[��X��J+w-+^ҩY��Jv �	bWZ}	� ����,�#dA���?��f�0(�����3���c[[S�����A�C�*�W{�N�o����c =�38�
҆!�n�T+Z�{�w�UIj**��i�����Y���	t rd�Q�%4 �k��2����3>ܮŉ ����a?��ׯ��;@zF��}^=� �+�}�������}\)�}SpRA�Sy�	l��$�DA���L�V8$o��Vw�.�e@���̫�IH-`6���-�W�~''8@[C�+�?Y� �����U���yUR�	�aʢ�o8^��p>[U� H=9&�"'k `�ZUt���������R���.�qz�a��x��4c%~�j8*�wUH�pY]^��4�Y���k9�6$�a����y��A��f��> U�-��?p�0�Ζ�T>�a��w���]8�U��Ø;�rvq%K���� x��n�(ǃ���x�������#�\iƼ��1T$j���FL�(�\�9~��e�I����E���ȭF�0 ��O%�3 �bc�1�/]\h�9>g�ݰO�g�w�b��v� �ZO ���+�4\^-}�\��x��Ȁ�EO�����ww��͍<>nm>�9���p>k�ˡ�p��.�Q}�
�/�Ҹ�+�|�wY?�e�a�~o����H ��T�׃|^k��1��T��y#KTOUa�ާ0�$1-��v8GT�T�]A�f��`��{�
ZB�Hxpn�a/u�1]���=�	I�圯�y�9�D�h���N`;i�shf!�;��p�u]*�I�F��@���,5�+��휆�,���,���lq��̊���������}_�yP���������pF["�M��r���dQ��-6������.�ق�n�{��{��<��c�{��>�>��3U�4�5�E ��OԚ~b?����^Ho�՘?n���<
,���lD�8q������#,�x8�
 *�)U��B�0�)���h�`��a�Rmn�X>a.��@�%��"F=	W�+3���U���Y|�Ts��mmnp2 �zB�5�0�-�)�za���Lf�u��� yљ�/�H���R3A�S�
�ڬA=�'ͩ�B�� UO:#�]���,�^,+F�L���i����}k'�|.K��L-mc�HG0���ś�a;�ȁ�G�V�w�ө��D��}�K5�^<�㜔GU��g:�L�b���6��Mmj_�6 S��Ԧ6�/����T��:��.�Y���2g@,�<�/�JV%X`����eu���	*�X�m�����X�����u�+Y,�	���-EB�[CIA��f!P�-��w�"�Պ���a�`^��v���>����X�ɧo��q-�+y�����cx�f ���H b>�Qy��:�b1GK�$�C� ���J�cTՇs��q�
����a�N�>������$��=N �k�w@�e=(݅s����P�
�T�2 �^��Z�"NҊ��, J�sN?��� bN�$��*H�����*A�+��a���ev�X���0,���`Kn��W:�]sS������9�ϞXDy��;h_lQ�*��	ǟ��	�!��Z���Lq�0������)�`�g
(h�����lQǿ鮸e��Nm+v�S����� ��N�A,�xu��لc@���Q��	'nh�dV4<�T��8����$��WU�t��T�Jb�$g�:y���؝����؀�ga�rqq��^{!%����X>K ;l���~-���%�vG3#��v����=S�כ���U�Z o��"��+j�Jx��ZX��^Z�#��u�Y�,�� j^���2�ly��=�p�����s����o|�}����]y���P�>Z�(�*�9爡� !�w �m���Fn��x��9�b1c?��1'��,�۫�A�s4}����X]�@�`i�tҠp�o�WU5TQM���H]�#lW��U҄�k����_M}���ZI_x��/,|�-�n�Ga7ER�(8o!�=�>��CL5Ȗ���Ʋ+ܚ��0�,��h������i��Y�놬�m8?w7�ч�s�ZB?�����o�7Gn@�@o�gr����m����M��#Itlf>��6Pz`4�������*�{���)�jC�����=�V�^�R��|�p��,� 6�7��V�'$�5X�&�����sM��yo��͇:gx�jsV2CJIY�i񹡱0s\gZ�%�|�B���[#1�	K�B��N�#���N���K��M!�:�?��,V�,z�˹,Cxz��qZP%�����������ܭC�_\�☖N�?���)�N+�pn���y����͢�+N�P��)o5��V{��f'm�8L��1����w�o��F?��?h���#Qp}V̕ ��l皡ߘRc�3/`�UD�V� 
��)���ϕ�b�e�����L�X�G�>�����b��)� Q�4�s�Gjv�{,.˘�va��Ҥ 9�v�����pe`5��B�^��lMk�'��7	C��>�ؐ�<e��³��6/�/�I�ML����W�M$?iC�V �7�m7(jK�n	�8΍�Q�da>�J���0��Y���Q u���DH�֓�\,$:�w�4\��ω��f0`�0�gbӕ'̐Se"��]l��(��s�Ĕ �ϟ���7��OdjS��Ԧ���&djS��Ԧ�����Q�W�\̵"�� �8,�Q�3A���M���w��Qb�����V?�%_hV�Zp����ڒhe�Zt�)��۲>�݆U�\������"|�g7�a��s�U_�G�$U;*4������ݚ� "�@kXP�ZK��S9��D�,^ �q�V�" �z��JX��o}�1���|�}V##���q��.��6\ ) ��=��'O[�*�ڀ��zR�:X����~Th�:=&���z�tJ5�)XNm� Uc�&	���D�%��	
�O]�DI�Xp8U*p��z��V�ImƸ�2ª	�Tѿ52l�����{���c����dhj�N���@�R�GG�<�V���aoh]��QA�ؼ�+8��Z��QZ���lYR�A:�� ֱ:D�e�^�1��۰8��_�k��۩��r�|Wwx_v�W]knI�WsS����|?Ѩh1"���O�ь@�Ď+�1�΀���L�qk-�&��}�I���ɩ.Ax5�����Q��f-A��tP2�\����ʓ�Ζ�m����e�t�sT  �l	�.@@ ���;F��:b�K��8��Vf�$TҬQp�N+���c�Ԭ�?H������u�L� �0�*O�|��+�A�<�� @X��m����zX�=�j�S�L������=�e8�Z�`���Xt��8gI��L�e��?^p}=3�Ck�ܮ8cU�Y
AA��/ǌ�3w�󢖈�]d+��6���
9⚷�������΍tV�*̭�0���΃ȝ��$���cn�p���留iqgʏ��άB7"� ��������Uo޼��mO�^s�����A며o *1O���f+�cIз�xU~��0���	����P�$I�h.Wr���0f@�@���_���ɳ���0G��^�+��o=T^Сt�y���<�Ϡ$����= ����2�P%O�^��S���Z֧>��a&�Y��B�*�������/�}[�9.+��9r��m��kZυ�Yxp��Z��^���F��o~$?������Z����-5���X�6�ny�ѧ�p��g�/ð~j;��+�>Wr�X?�r�$թ�^@���R3�@
�97.�*Q[c�F�F�M�{5�.ے�T�����hMՇ9�U���3�>�YW|���W�(@���]R��6�G�ċz5#��1��y�h�w��ò?t�F���@	����?�S4GM�{F�����V�9[}V�Mu����<�j/���0�#��0���l���#i|@�9j�'F�_ا&|^��|�e�pY��sA�P��uka�PB�rȜ22�?C�ra��ϕ|�Tf���S�8�G�Oj�)����ϙY2c�{l9E��C_�BV8P��x��ul�*Ψ�k�p����Ԧ6��M���&djS��Ԧ�����e�~�Ӆ�Iá��oaQ@�U����ch�A�mV����ڢ��W<���>X^a�=?��zBkY�aT��O?Յm��v�7_?n������4��0�Ԏ�|a��<�����/�p�����ýlH�(�����%�c����6$hZ�������,5`�U�-�o^���|~Y.���m�������m `8�
�kQ		1II@ �C�W8��%�ҤЌ,O"�V,�:���ma��7p���T��%QA����ZQ�iN���`�n�hv�UT���uQ��v�JH��0��w���PZ�(�U,kAA5(�+*_���Y��
-9~��5%I�O� V�}?� oÿaݦ՝U_]�vR��p"��;����=^��v^�į�[��mT�W/�"�ϩoq4�8��>���F�����v����W�Z'<����Bu)�Q�6;P��(Ò���U'�h �Nmi���d U'�<�K��A���أ���x
"zJZ�oj�� �<�ԇ��T�F �+%K
Vc��M�+=	��KPq��k�mI3Ȇ���2�rf�U���xSˠ\���$0�T�)���hN6 i ����^���׷�w^��ס��h� In�ٳgruy�kv���.\���N6a�BxC�C/���%�-+�� 1��XHs�+o�� ?8N"Z�/X?�<����r<9�q�psl`\�U�3ĭ�0j��ԶL���2A� �q߀�����2��b3KU��I�ټr��AԳ�9�Կ��R]G�Pd�2��IJre�@V�%U����G���ן|����3s�5bs1�t�� '��[���v#���l��RP��1�9��UU7d<)(
B ;	�p��'3�=��6P\���*5��,�4�zP;`{���N�B9B'\G�	�L����W��JG(�j�wa&@d�(`��� ��Z"gen����M�צ�+�^����Z�*ȕ}3���7�� ŵI�ν	�:��pO��~.Ϟ�ð��}�o���?����o*�}8���4�7����L*�O���J��v��q�wZQ��0T%�3h�d��)�s�sQ��x�d-b�O�uSN����5��6i̫���Fՙ#���m<1���ZJ��Hz�T�Y-ƴ���HO�����J�������=�af��3k*�I-
�m��e\���������������s�{7���@F���=�x���f��a,QR�$�����$�"�O�c�5��@l8��V>� �L���~�*����ߦ�Rң����m^�w��w�������<SF���	Ϫi�����8!C��\�H�<���9d��

����buP0ז��g�L���'�B;#������MmjS�2�� ��Ԧ6��}���q�J���N�]����ii�.]7���Qy�^��i�b���Z�����
x�6 ��>Y����+N������E~�r&�O^w�$���͎�S������� �kxQϔ���p�+�l4Ä+L%N��|����,ԅ�f���@�y0�~$��&��]�j?0 -���h��L�a���d�-���@u$U�oݯV�u�ba��B��J��~��k��P���� ��F��z�,�I�Y`7�*�.��ȑ���MWK��9�Ze<�M����^A��yN| �]ķPP�lE�3%$�Wو��B���N�C%�,�uO����G!�-�� ��)���4a�>>�����Q��*K�B�r��8��u�L0��B��:�d�rZK$O�D\�����}�mM�b
�T�DU䐃�ܞǳ��V�j v���g��F����?o�Z�/�c�E��*������A�v~��H�`�ڊB&��j��cK2�r�$��y7��MYU���j���z�ɛ4U�:I�y2��j-赳�T�%��۾Q2��l�8�,��T]8�0�_��K��"p��՚��'�E7 �PA{>��\��E|���$l..o�ŋ��㶇���dw�~���@�U�� �w�:�%��m9 �b%���+�c��g����q�J�L�bؗc������w�k?�z�U�!/ڦE�lfV'Ij���n��t��yf ���J	�ZIڤK45�,V�wzoQŒ͝ B[���,�D�� Ω�N�#Ղ�aMX��kX��T� <���[�n�y��D�1��t���\�=���e�`j�5}���qGu��
�����m��M�~�ix��r4�Pj��X��64ϟo�z�T��y��B_NTYcdw�vL)�3+�#'W�b�(����)��s�_'%�L!��=]�4����ύ��s���?c�@1���=8�}ݛϕg�;�gB���9��fT�P�̉m�$���3��|�;%����礃d��
$i��u�AX�,�3��,g��@j�8�yB��D:�@�J�*�J���y���8��m����Lj��nB�}�a�1�(�U&��DM���>�Ls!��������O�~��H�]ט������(�H,�Cǟ��0��]ݏ;����b@��T��N0׀��܊���so���!���N���K	R����0ø����l�(� ��`U~F�:�$���� x��=��{��[��D�ѿ��-��O�d<�?����m��,�Ĳ@j5c>>�f�?�c�XAC_ca�f@���������}��3�z��ZI��ծx�7��2頖�DI���������ܫ�N�S��Ԧ6�/I���MmjS���T�U���m_�	��6TV!��_��ú.c�6Aj���Is98���*B��� �����ɒ��Ay<P��&���-<�62j�C�O���S@��U��UJ���-���G�`�/4�a�Y�Ġ�,hr;��H��gg.	CJ�U�`t�lI�Vu�	�T���އsx��	!���þ�����<^4�y[��k'$G���`�.	�t���-<�
�x5Z�` ��ǉw�݇m��8Tp�X�ZXq�U	�K ��*]�y&E���1��.nI~��YR�	`����QC<?[��@�[d	�=�*T��8��p����`��T�}��T�A݊
�,P��i|m͝ �; \I�9����|!�ż�|�"zM�)PU�w��S��pb�;�����������U�jѼ��3?�<����p�W��,��vg��}��cx�o{��P�W�{�9L2����+�*z�-��`S��������0n�'���{d����P����UK�p�tT����
fô�;8`�?�:ż�X.~�a�;�����Ȋr{$z.@�CN�/(�nk�۝M�)����;�Vb�v¶�a>�펲\j�7�3B�s���O�I�s]��d���&����Z�l���?���%� `M�F�5<�+�0��ԫ����r�X�9�cF�a�㵟ϖ2�rd�FI�6' j1�ho5�*aڨ��	�ϸ�R��]�hH� �x����2�|p��������V3�����������"�¯�q�����K$��j�GB$��~6U=��
�y��,o䣻G���OI��37����5�O]]]1���w_�k�$=���d�n��p� ձf�Mۖ&�K�B5 ������q������]���e��m��A�B����/��lw�T�!�*�z#�@�)�;T���D�t2��p*���0�Q�L�%�8�A�8��̊�={<��nq���1�P�9=����uxmޫ 0n�H��q�:��C���Z���DIM�,��tᘎ#~=<ne�~+���k��Y���LƤdrj#�� mu� ����Rn�ò��/�Ixb�VyI��*M�,����<4��uNX�
;���yO�+q&�����Q��#�c���%�':+n`�gM0�d�*�|$D��%,T�iVj��*vv=�l0�Ϙ�nFE���0��C,-����`�Z�y�5�Ͽ���=���?#f��Mm^ñs+�Pbǵy��Xxʥ��`��m�l���t��S�c� ���B�b�L� ���X���l�2H�Z��<�s[�"���H��l�������|��* c��ǳ����㍍gU{.���YdjK�M'� 1�W���gׂ���7ٚ�����/��;?�P�6��Mmj��m"@�6��Mmj����L+�iͤ�'l@* q��3�DV��B��Q�[T>X�a%�� � �3T����7��X�C>l	��FUn�#���C�A�����L�*�ժ 8y<��2�)��yX��:��eǞU�h�B�̆��$�[���C����a�}Ē�y��@7�T���#��v#]@�Iڰ��4�r!XR�	�< �����<�V7��QFȗ��l��a1 ^H�gd�}Ѡ�ʀ�s��Hd�	��$�k�1����K�NG�2��/��}��dF��3XD�;�WI���D�~��i�M�,�QQ� �80vl�p���#zX>�(ۣU+�յ
��j,��z	N�6��P@\,�>�'�*� qb�		Wf��b��.Ɖ��nՂ��m��n��!����ɀ��y# (��+��)$7z��|w���D�
�n���bW��gd��?�ɁHtW���;����!C �E��6]���Q�� Vf	me�g���`N3 b�ϯ	�Ci��&����x�;@�#�s��B��8!��P�}AI��̒c�I�Ss-6�Q��@�Hc�B/3�  �ֻ�Z�Q��#�Y7a�D��P�`>�v�R�u>k1[�W��srn���z����,���J�}�<���cWUT+K��_\�l�����ۻ;��*��j9w���1�8��;i���u�<��6̹Jd��X*�|
���"@�BBr ���y����76�b_����+�ox�Wu?�|.��s�����Ҙ�O��� q����ln*"�ȏ�on��_|�W~�ʼe�d��ju)��|�B�=��ɷ��|�f�/�܅ؔ�K�IMw�n���r%����8C���J�T�z$�B܆>w���$��O��}~�u�\�@4��,y`�H8F��m���*2����=T���ү��������1�	?�s�طñ����=���%���T�-4c�Ʌ�I�m Nn�j��f�r	��G}$�?~�O?��ݜ�c>!k,�)���.f�4���"��ju'�*5h��t��7z�B�@�T�S2n�9a\�jCE�g�FHx��SW7�m��jAbc-����u���H]4��>%�]Y�6���$�7:�P�y��`˄g;<sᾙv�����L�^��X�h������@|T�ɶ��gD�����i�̤���I��[��6�D��N�:�0n�w�Jr���x:"˺��WoÏ��f�?w�(�cP�T%8��$��W6x|djQd�L;�3Ezp�ӑ���ڸ�e���H���K�|�6g�y���l'���y^�Ye�Z3�W\���F�P�X
m��LP5���~�WY�$��Ԧ6�/K���MmjS��oD+f�0XP��|.Y "�B���#3*��jh��>0 f���]z*�E�UHǭ���g�p��>�i<�Ow���a��*��\M� 5����N�
A��� V��-���=��8p�2Ҭ6�
����hPM�\���BLH�b
V\$ZVh���[eg�`�c`z�*gHQI]v�50[� /�;_�v}�/�!Z1�F���f˄y]P��<�}�j@�F��_�L,�r��>���m���2ЁH�o  	캔�I@����b�c�����P��c;l}O�8@􄌹&��� ��s�Kiow�Zq����}�� ��"Q 
 T>3��1�H�-��NA�!��Vٶ5ϋ�@J���"�pt���~0�y�}Lt�}�wD\������E׃ax@G/f?��m 2��"b�<� AC�� D �jU��*a�5�վ�
��F������`u�g�u����$?�:���ר�~N��}��\�f4�!��9�y]<P�5�FD��p���;4p�->И�0W^ m*|g�~�!ç$HU�5�+��S��+x�WC�q��� ���>�yK�Z8F̛1-��0�,e���N���|.2�p=01�#�$r���_�
�s8��S��~��e���2��C�<�A���!��c�-�Ѳ�40�\#H�"g�=���t02rN��X�y)��}+�$�}����}��(^1��G Y�,�[�t~F�r�]n����*62g��8^M-�/�k)mUy�]�R~�����g[Ӄ��c=?_ɋ/�w^�˗/y�����61��I6������
�D+�ծ���*�D��96��w
�����΢����%�����#;>��l��Ά��cSŵ�_8jſ)G�0w������ ?2���F4[D-�r>'0��9��<��uc�Ω 1'�@0��fzM�:�`g%9��󱇨s�6��8��( �{3N�fj�Nt;ؿ7��ȇ����=�+��[�Ї��,̃�s�J/N�2��_���Ƶ���ߓ�ͨ��%�J�V��128��֊vw	c�_竔k��j����qu1�R��=��H��VKO<ȶ��z>�Q�M�B��H���+H�BY�i�|V�d.�?��B�#�:1�i!rqZ" p�=F��Ɣh�i?�F�>Ga��=��dU�O�It����N�6��&�yPKǲ?W H�eDª�tĤ�$W��3��M����Y�sN;2iz£��>�Dځ�a1
��Si��fؾ���HC�Z�Z�Ԑ(]�-��M��Юm4� ��š|�`�~̴�Q�`<��1�P�����Ka#���E(P;՚�ѰP������Z���r%��}W���)wjS��Ԧ�[�&djS��Ԧ������V�b��!�5�U�B���"x��Ӯ@I���զ��U�u�ҋ��<�q�e�VQ��bXw����g��`EV ��α��P��-�ɧ'��?p�
@"��J˪��r>+%1������Y-��ӏ�n}��fa�aU鵅B
��Yy�*d�]��1^��f�@�{z,<���̂�����]
��Py�ϰ`ezX�,�J�ZSEx�̂����k�eĬl'0d�pT�֍�fA�PJ�u;��!P�~DN
 "T§�+ěNm�pW��v4vѰ/��  �l��7��2����~B��Hm�@j�O�(�1,���̪�T;B�0�)`�JVUx�}��Y�	(>R��1ÿ��u_�g�5Ȏ��`	3&0��c���5�`p��Yakċ�*:fBıY�D"=�[9���Q��Ȫ������;���j?J�F*�s ��$H2WL�H�%z�q�Y��c���*�I	Z9:ퟁ�9T7�c�*nS2��R�/����/Q�2�P��I�2��)O�q�{���sZ4����# �
��g��X�%g&����'?����j6P���`)05�J�(#[Պ�� o�-�B�mRm�	����5AL �y��ܿ㑯�]]�n�� Q��}c�p/w������=�p	���͛0��+_��f���م�P���$���p��}+��^�0�`{����f	�$+���AJ��<����\��zj^M�\ ��oX{�� ���1�$�9��L֭��Nژa���H}t�U�wJ�3�D������è
�S2��ˉ�b�υ��(t
}��t'������%j������<������ʜ�OU��CfԚ�QP̔fQGw�LX}��#�Mb(�é�Q)�YFrǑ�g�{�L�5��O�Q�H�7G����ć��a�x�
�cyT{(-A�����z�UrFK5�9��̢�a�v��`l�Q�1�N�V��(A6���y� ��r�A��[R�>��k���d.ދmi�H�+'��K3�58q�>+�t�.����}x�8�p-r*��0Ԗ�qu���{�=�z�߸/��C�G�S�=>�d�\�4?��nȕ���!
Oj�� ��5bdO��,<���j%����O۶Qq3Ryx�Ij�;iFVXc"���*#�C���\F�R�k�4N�5��X3��*3աf�Q5��|��=��j�N�
C��<�}wPop>G_�-fKPrjQ�j�H��k���q�n�L�;=DJ��|"�0Q5�ZC�p��#�H��ߘ�ԉ!���G��cdo������H�N��R��(����'�zB~�4T��%6[�h~W.�+����߶G%�#a��g�{Aa�Ǽ�\b�l�
��4��gb��sLf�kd)������Y ���Jb���̏����B>}��LmjS��Ծ<m"@�6��Mmj��� ����$���v��H��b��Q�r課�C��;�E�j��o���H lc�eX���p��,�k�x�@�{V����|&�b.�<!P�������J^\_�W����9S���" ��gWr}uŪB7h��}��9�9����e�ޑ�9�DX,gK����mg��]<Z	�oY�K`>�j��St o+��$�y��j�%�d8�� �VͦR �	i��յz~(���+<b�� �:��֬n.��;�@I�!��1�Y��.\s� ���k���MI� Z%[0+%e��U�B9SW�8��WL���%lQP��p��u�r (�D�h�׷�:���_DX����_p�-����"\�����U&��͙y��y�WM13/����
�f_ ؾ�H�Q�Q{}�h(�ok��WEJn�XI��d�[���I4%mr@2�S���<vP�C�AֹmI'*��𾹩���z�5��wʚc	 ��Lm��p}��v8�ma�1�p�s*`�Y�35q��Ta�4�F�,dI8���� `�xNKI`�l�b�7 �O���zJ�*h�̘�0��	��UM�W�-���z�c+U��;~��`(9C��[VBP+����s(LE@/�$�3"9 �0�m�G��ɢ4��I)�V%�'(ɒ�3t�A�l�ѱba���F@x�m��� ��S��*�|���pN�:(� ��j�<anQ̠��Mt��S%�M\�pz�}b>���c�*��b�q_3�#����|��i�kvۭT |*��	�R< __^G�n�~���uuK� ���'���ǃ��wj�����|�$�����#��
YCa<S�<�ϡlH֠?-�p~#�4�[S{�Jr�"ނ���U[��0�H��VtJz��Dg$Z�9ux?r�tX?�x��nǀ�BKL�q�����G����ϥ,�v���n޾e�{��S�a��|��9B�ֲS0�]����}����
�v��X�*����?"�#���Vk1%���r\�x�øK	���Q���.Ζ�zϥ½�s�\�� (�.W�I��A���9'�5���"������a��
3y`YV�y�A��A|�7�~~&�hN�xOƽ.�J��ZU!�d���syxhHJ,ýkq~&�C��ox�y�/���|b�<������+
�M���(ݩ�����B_��sͱ�O��Y�i ��?:^��K��x��*$ʝ�ۇ�����V�53f��>�]#Si��WIf�K	���6�x�(<�4�&Z���p_B����Hx�Q:��#��g�|b��� ��xG�wo�1Kf��Zo�cx��YA��lU���lN*M�>���7�+_������������h*�p?��d����+Rf�T�y���gR��½�����#�Hӓ\���EVmV_9Uy`����n���>>ų�L�����yv6��7���������5�%�(A}��y�3�Õ��CeQj��*� �P�C�$3�Ԛ��Gn�C"�h�j�$�v��׾�RU�HH��x���</��拜{�^?�v���ZF�XN_�_�>�
���������k�c��G�$�����MmjS��ow���MmjS�������"�P��M)�<�nvw\�V�{�b!W�Z�h%s�uE���,�@�j/�^�$ȸ�U@8#�D%�s�+%W���d�#�ϱ0[�r 8��Q����þD���W�r�o���ʆ��y�3����ʂ���~uq���yQ�_A��bgo��&h���ʖ��q�4�PxN�4,�����h���dq҆J"1�y�6Yf�R��G4�Pj���+��V�|qN 6j�m�����e��d؄ϩ�/�"��:O%�%o�S�疸�Vg��{J'qb6j�Ek4 ,�P\�/����� �kʃ�@l�oU�m���u�6C�U� ��Hz;'������z0`�
�*�T7�����!p�-��3�b�l@D�+6�>��p%�+<\��!��}Fb^�yO$(84�V2Y�&aւ.�u��m?U�H�"�C�A��R��6�݃����+�������������2W�xh�Xs�wk�d��N3= 4j�N,*jk��E�<Ɠf)Q�2p6�H�p>�W:C�SV�C%�qRGv]��59Bn#��������]�S]�D�VNPG4� 8^�����O[�����%W՚U�*ly'���e�$9./����uԑ��g#�%K_� �G ��d ���}I�ǒ����Z��)�����9�/xܰ=��7Twe in�N��#�IP�hf��X��/W��Q^#���������{Kj�0`?��fG�l+U���l�Te�W�7s.RVE��2�/��h��$D 
�>�>�𰓛�[م�\Zպg��JK��������¥�|�R^�z%Ϟ=#�r<�6���*u��G�_�U��c%d�6s���k�p_�JEIS��@r�Him���� =R�p��}�V8�����4d/F�:.���m Uy@j#RP��=ڕUr�J���z���[̗�ϜO���C�O�����pef�͊^�֙=UV�$k}>C���')â�c��Ui:��ZvTp�?���}�,%�!Bͧ�'2�����5TJa�i��w��0I��XN�JH7�p���(@zY�YK��*	��;Y�/�<,��:��e_�����^�R�m���b�=�-,4���0����E�sٕ���/XH�fn�钩Hz�g���ꒄE�H+*S��8=*�r��9�15��6y�{ݘ�fۙ���f���K��r*Cp~�a������eI��_��~�g�75��ྟ�}��l �[ys���C�[�����/I��8�33?L����Xc׬O�x*fU2*��i-�s'ɗ�fn�>��X�@H%f��sCn���͉�~ ��v��l�h�*E'vJ3��|�WQ�$��#2�\{�<�U|� [,�dy~&���0�a�߄kMU���≚dXM2
�B��aN�~v�}<�g>����迕_M;��Ԧ6���6�� ��Ԧ6���F5,R��K�_��.��U�dg�$�#�,�-�B(,TQ��*��YX�c��X����g�oo�d��S��S>6��������pg�Wv� L�S��D��Q���xO���KZ�`Mwqq)�g�f����wV���g ��n!�� 	jT+3_[���vh��jk�ƺ��"���;:�!Tu��Q�n�����T>�MB���k��$Pl`���KA|]db5���H3A��T��:r�շXfF�O{E��@V�{��Q���P���0�,�3�/�5CC����K� "�sQ�9$:�����Gs:AH��Dm~��s����s� lw� pU�i����[��V*v=�P�M��qXm��b�I߆_߇�,�|_��˟<;���׃y�mX������~��?����x����z�%@�~k)ڵ5��hQ(��D�x��!�:�@k �8� ?6�S��!D/����SH��)9~��d��cU���-����ٿ���o S�����Hr�Q��L���Y�ǨF5j��|��A�T�G�+�� R}4�M��wo��C-�4�`<��ۓ�q��x�ʼ�i���q| hҸ��uT��n	+�g�3�k��RYU,$[��M8Q�,�Nn���1J�p�f���Q�A����p][˄б��B�7�f�z�B�������*2��"|^G��j���s�2��w����j�B�N���9��<���ٴ�`����*�b�Z8v̙�W�??<��9�����V6�R��`m����O����J��zF�ǫ�/8.qC,]^�~#�ͽ�w{V`��0+!|��}��� ��џ�Œ� v��v�7�9U�E�1s���p,��*dJ@K�DF�(��>���k��IZi<��S!�m`?1���;�.N'�:�林"�{���1�y`�1��R����_�t8'Ǒ�r���=�}���0�:z�HTyT��"k��e�.m�j���m���:H�{kN;*~�шs�>�PU�M�=�Ҍ2��$�ےHE_,�P�����i��i���Ԓ���b��P��|��owt*����16����@"�
���(�ra$��+�߀E�+�g��of��"��(��l�Z4Ph~	�)��a^�! ��.�*��e�>�̵D��<�^�	MM��e�v�g@��3�G�6�Z%���R����[e�}��������?n��j�DSAV��V�y|��`��O����J*9���h�ϐC���Ҕ��/@`�&�R��79���f�K��(1�v��`�^��+1�A$7�AՈ�Ø����2~V#��	�2�ζ��G�(���Z[hO	r$E�X-TM���J�	�+ZP1��a�[R�@T9E��Ԧ6��M�K�&djS��Ԧ�� z��W��;f[`ɇ*E-�N�;�����S�A	( � ����?�P޾}+���X(��C�Pe��5��V�P61$`��a�[��ã$}�a��T)��f����[9��A��/h������l���",,������<�}5ݱ�<z����U|J� �T���YUb�$����c9�BP� G�9�Ɵ���g)�4 z��� HҰ�qP�4v-`������T�h�b6���P�1���"~�W!���EMt?��^KS#�Rnv/�^tj��`Ki$�_*`���dC��m㡡a�<OX���P��$�m�������t#�HF��ƴ�����㸝��7O�.�����{����B�����fK�dו���1fDN5(�� � �&��҃�����I���Hfz�LflQIu7A�A5eV���}�Yk���#����eE�{��?g?{�VǶ��3q���*��WY}��7f2��1�\#ߵ5��Ҫ;����q���uV�1��5�\����� ����q^'6�M� �
���ɭ&�FH�4���k����ߎ����8�yށx?�)�4 GBɯ(5����KF�7>3�	�`Z�6��GV��X�jK�Ҝ���N� G�9��b�O�&��k����q3fUq��]��y�ČSdjA�.Ӥ�l�qd����3W�+�K��@������u>���r!��0�:7������q��ll�_C������s�bۖZ�-"7�I�B}����Z��H�>{*r_O��3)�8i	��+>>d�D�%�'<��/���,V�ϯ�q��a4�!�W��><<�����o�&ǧ��7�q�<}�D�Ξ��{"/_���� $!�� fƒIX09 +Dy�p�b�X�ĭ�gc/�J�CNpL�9D!�6U �X��R3u���~8��5��=?z������ϩ\em�h�u��"���M{].��������Lf��i�wq�߇sE�y?.������qF�;�Ny��p�0N���T�
��@����q���4<���fMp/�����ZB�|�7d=!U�9WY�;�U�s��GH�CJjb�8,٥�Z��_ْh��BL����b�'
5V&�X�P�GB�zǽt���:�me�$�8�fA:z�Lջ�9��B�Ij =��
z�I�"5����E��zl��@�hp��w�� �F�D$�kG���c<��8b��	�]��EQ�ē���w����ᆉyݍ1?r:��&��!�b6_3�����d׿��9@���s�OLW�t#��<Yn�Db]��24�ުT�J�,`�f��x�*
��ϵE�A.���X�}�V��W��ykJ̢�KZL�f�!X�@(�}���Ud�PRT�,��VʸVW-��`S4K�a�D�� �wn��І6��}�� �mhC���Y�4����C�	4�ߩ�d&��ߌ*��$W����nU����\��XA�M݆RB*�!;2
?��=)6k5S�ƚ����c�E� ��Lz*@vgR�5���7��P�ڲ�� 3����/���p�!7�|�;�MY�=mM�`�:�Ɛ`CWYG�()���5��I��f�ݺtK���pl-'�.1���~�����S�C<��0l"���h]&BM�Sq�5�V�㻋u�K4��d�V
2��c�&��D����T�"�N~	I��&=
V'���
**��Z��U>;Q��C	����s�Y�Z�8v[�C����y$H na�O������5O4����N�<CBρ&��xb��G��W���{O.���s��=BR��~���Y<c�`^�+���Kgq�ڵ�w���C��R6m�<PNk5����8�1R�^��~^�����oYj�x�7U0��H��q��(���n���M�cB�wh�CڅQy��V��S��g	䣢�� e�Q >5 nke`E��H�E̪�� !ё���� FPY�3���8�3��NJĖ���O�C� ��H�b�HF�xL�s���m�cd�t�n�ҊgT>3������r�a�(]#�c���N*YU�LQ�?ŉ�Ա��Gk�*�w���� 8���o� Ď���(�d�O	6����+���)���@'5o�}
<UԉW���}��r�ؔDx%K�%L�]�H�E�kL�b��1�d	(��d4��͢�Ն���ɣ3�ݗ��e�_?&	A��d� ��+���ޥ�<��6ܛ��/������精^0鸫>�a%�T�*��A� <%�6�$w��!͌=����D}�,�:;����>A4�@�m&�R��u�3w����n�@���4)\�V�/�72b�Ɗ6�)#Д��*���ZI��R�1���&��`%����[��(���H����*̉>(��t��j:�
��Ϣ3��:�+�(�s�OJ8.ܵ���ݐ]%� �%w
�u }�)��(�@��庠?�@&*�W0(��q�>͌}�� �BM�w��%XSD����sR�?�dG_"�O�:8��2��>��'&�ԗwK�Ҕ�Ē�/���6�@�Q�1 ~A���B9��5$�1��O�I|ܣ,�6e�e� s� :���S��o��H���	z�����V��*�] � 6A1N�q"�̺Y`�{�gE�����Uݱ�����:&֚������� �S�=W��䦏B
2�
 !�խ���d�j��b�=�ɫ2}�w�қ-6&/����w"�_�ʕ��*�a�}D���o�K���=����{0�f���9
�k� �2r!ˆ���d���s\FЇ�,�{b�hu)o��2��mhC��W ��mhC�7�^�}G�z���uzH�jH?=={f�w[c�d�|���u�\����}lli�7�`_P�����W�ru %b�4ɮRAi����U�Y��E"�U�avu�-�?
�� ��frx|��tLf�uB�U&<�{g�7ϐ>QMp� ��|>�c����粡Y�,~K^4���)+K�X�պ��\Y�$�\��CX��$�(������$N�
W4�]��à�F&������iDO�vQ@�c�5f �+�=X'K&k3FGQ��3�l����<��m�����Ɍ]�+2 �MF��R���vM"�w9�ә �f�v�]M�M��(����0;���R(X��Ǧ�퀀�DPI��3*�~��_�Xv�����g=�جP��8���g��>8����F%�']Fs ���:�63��v�
�_�����K�x���|�z���.}0����V�Yo*��n:���tq�����[(M�dM�h� ���$S�(���\�&��8�1��!�RI��d����iZ�3��K��g�ű�,��l�%�QO���#���?���CbrQv�Z���?�i>׷o	�����Y���,kJ�dqL���>S���������3�P��,
�`��A5v�}?�H�,�����t�>F��IQr��_%��n�ےI�cNB���T�1���L����}@�:���P��G�uWW��F!{����+K�iD��2�M�q��z���X�Ҍ�&ϐ�[/3`�T��˰�\_ћ
�|����{$rSO�{��R;����`}ܺu*o������kC0�/./�ɣ���W_����K`���XՏy���,�dX/�{��e�E�-�k���g�����t�`T�D���,e�,(զ71��ߓߙ��x�k�c��x�"S�f�i˘�k���)�Ne�<fD��ok�e�Z�(������-�~�sBy��l�������&]\u�c�Ww��Ύ�����$�b�	�D���ở�I�~���HMNH�1�B\�X�	p &� �"ք�[��}A�D�t�	lT6���ݭg =����fɸ��p�4d�D�z\��Ypѿ߉H���dp?�t���AQ��	�`�J�گW<�lR��5� gZ�P����Q/D���~�Dc�^i������E�`#�Z�t��_8�Ѹ?��7�@9��P�����;Y��I`�1c<0��#v�p�#��j�	�:�����s/��b�ؚ�۪gɓ��&l];A����>�����]ݪ���`����������$��2!�'E�y��#Ŀ���I/��x�}��?�w���%������7���Y7���� ����
,ܧ�_<��?���Qtz�4�c��І6��}{� �mhC�оі�� ۰�;O��@%4LN��$lt��q|p,�����D��ɶ܈��LXO�3�s���~�5& 2^��&m!�H�0Wh^�M��a˱A�j�JLT����-�	�ڐC).*���Ae:ֲ�,�z��	H\�YŞq#Y�,��&:�� �M$q�<⦔t$Y���$�,\_�����I'��!L@�A���`� �U���V�Q���y��>��W�.Y޼"���<]�VTG�T�v�#��hT_� ��h@���笲D�Z}
�\ۊ�a|�&��t�~��� �CbI�l���L�	�7�I�敕^)	�tng��	;Z���Yf��q�s��>�Ց�+Y))��U���D�&��@�m�%��S�v��;�qR�5qSp4O�x�>$��5Y'���l�ߓ�޵-=^��$�pp��O��q���:�v@���P^�?=���W.9�6�T��`L���9Ty"��u&�t��a��ɸ��>�gT&�$��j��H��	��B�d��&MҚ	yA�53�	�5��
���zc?	��H���+J��{^�*G��i8'6��N���&_ӏ�ῑ��l�u}����A��U���DMp��^DHơ�ü,4y�$%�q�,�-�B�oR&xy+k�GhZ-�	�bkl,Ċq6aro���QC�z� ��OF�?բ$�
15��X�w�Q���%��d��P��(cb��s�}2z�!���J�p��5$y��s���@f�j�q)���Q�����	��a��������֫�%����6\�J���>�q��V'���'8�,�d���ܻO^������!�Ћ�R<�\��=�G_}%W�W4$��Z��٘�����Ik�tyX��UgrV�D�Z,;�;7���u�$��&�X�.�����J�*��(ǎ�}�7Ž�Tｃ�0����11��l�cz4�2�4V���%�����.�� ��X~��1δ��Hqlc�}�R��w��j��&���{
� ��d�l��&_�ß��!WY��LMH7�㠥�P��}!�^�m�a�g^?|�
��c��i�/�<��Ѧ\�g+02z��%����]hx�B�k���Ddx}��G���m�=I���,є��I�ida�&�Φ�	�ԝL���Q
￳A(�T�3�l�~H-�v,�����8u��\{{l��(7�B����+z����ث�,��^O��\��7*G0��}.!Y�21�������*{�f���9-��65�2!跢󤁄�8��w��{tU�8��aKy�=��T�qp�{	v���sv�+V"&�%*�
�����l�
8��c�5�5�o�B��
T�9�PD)Js0?��B�-��ð��{ߓ�/�D>����i��C�l2%��퀦<��s��/>���WϞ>�0H�n��w����mhCڷ� �І6���o����A�74�[��>�ޒ������U��ɜ����JN�ܕ�gZQn�l~����ݷ�a��ѣG��'�rÇM46uQSmx\Pv����V�4U���*�{SV!bCN��|L� ����d]_]���L��0q��5���'BMg�D�KP�MxTzWV�M��j#��=9-&�4�5fn�.��{�%�)c՚��.A�U��jr�hdZ�KX	�īzk&�ZA��y�Y��W��_I�h��t�jC4�7~�\,�����p��Oh�IV���i�z���S���3o�&sRu���Ǽ�~��4����7I'=�*��X&Ձ�̦�m��~4n&J`e� �&�5I�6��a�"a����I�� @d^+���R+h��e�:&�%�\�A��*�{	�Ώ�q��^��2Y~l�-�׋?j���X@����ҿ������4nU�ݯ�}@\+?�w�gTw �]�^��Ƶ�����T�,۱\l8K	��Y+xR(HP��%���K�	7H�����qJ�L�0���Z=z6��R�nx��<�+H��y
]���7q���D�f�z�`�A�JܓD���"��Q�(�Ҫ��¼J(?�xPbC�	��l��	N\7�L�DD�� $�Dm�h�ǩ?�5���}�t�,�k��/��(A6�Θ]��Z7<.f�/�jC\�RHd��?�F<�Y.g_i�rK�y��_)�2��H�n*Ʃ$��*=��� �Fzu����"�H���ʄ�2q�8�^�d����|�ٔ
�AW�r��B��<����v�i����;���A�)\��C�� �����H��|ִ��{Of�~aN]].��W�׿����8�pɄ-"'b2� �]X� ��J��i��'�z�(niL����Z3�F���C��0����껄��8��ý�J���*��k��h�m��of��13��/`��&��~��u���!&����R�Y
&�w�XY�C��#0�Bj*�;P̎��������)�(�c����}�s˙@m;��$SfIUU_��`�)�T�ƝV	�ת����Vc3�/Ĥ6��F��p�QK0t���<�h2�.����]/	T,�vR�~-x
�5@}� ��8�zh�&)�Y���.�kM�3�(��6tA7 w��<)VQ��I�I5�)$�9��d�(�k= T��dI�s��nMv?���c𮤟��ɤiAHK)�,��ҁ~����ar����͛��{�}���4�J��;" J�xF>T�FvL�N� Pdq��C@6\1�ka�g�
��'� )�o�.�$ΰ �Qԯ�����a
��� �DU�.���Ǆ$�Fe԰�{S	�D���t1�%�	��ɒ�S��� �4�����bU<�7�|C>��cy���e<Uv������s�� ��0���sOiq������}z7��?����ɳ4L�����5Q��І6���[� dhC�І����e�������x���?��{�������������S�= ��Bl�c5�),�S^�M��ߓw�}O��?�?����Y���Ugf||z"y6��r�\Zu'*�$��+4�Әsi�?��<}������տ��RL��@T�0*���1�1R�20�&�ܬ���:���g#�"�ڲ�N�'��)ZH
M�j���ÇryqM�rT�Wnؙ�M�A�Iu�׼vV�v��
n��/Z剤��d8([$5cu����P��\�.����(��U��`T���OU���HNMh�َ���̓DL~f]�8V�#�Ъ���C���$���C�l��P��*���;��@�3��e�Vi!��qD��Kػ�R���Fb�%��B�/�q��&�4��!�D�JMy�^M��^��'o����h�}�H��B�2^��߈+05U����q��v	\�ʙ6c�l��G�T����@�_Ols3{g��	���&� !$�1&��6fB�(��i�y�����@��z�1�`�3"�>7��kSc�X�3�`����O�&Q��k�j�6�XS�w�x�84�	�
#��1��i����@2H�A*i�D4�x4�Qp��g[v���4���u�8��8s �*S�|?���1�(;��f�T�G
�.W��F�a�b�$4���XŲz ���dӄ�^��8�����?)#	~���a|�1j9y�@�?	�;i��)7��#0~'��)��y�k��!�W��p�oʢ�`=��e�J�
�I[��5ޥ�^���S��
���0���|&2��r� >'���d��F�B_³��U:���%��U��-��332õ����E��'��L++���aX�ޕ۷o3�wrr���3��o?��ͯ�a����dbH#�'l8R�cx�`Mq�xeJ!!k5?�V�iL�Vd-� O� �3 ����� E\3bo?����]],���9a� ��j�s�K����8vF	���Y�����1&�c�*ڊ������������c,)3%S-�����Z`�ke����1��Iu�j۪g؋
\��R"	�A8�z��ք>���g��b<���zUh�XRk�|��W*�I�����-�)��Ic����Xٲ�q�ȏorn��F�<�Q�lxwLfS���+J��
�.��+�UbE�:�,��σ�
߭&j	���,��u�����L�;�@��è9?�yQ����nҽ
�iIy�&��9�P�L$UP#`�s�7�Re��Z���K�\^�$�(J!s#U5�Eį�l�b�̵�
��=��,:�$3�K�k5�fB�1�~e�pv��F����fS�o�V΢A���о-������D���T�F�5�Ը}[t��.�&�A�:k&�?I��2�k��1xK*���(N Y�X�x���-b��lóul�7�a}n�0`���ߖ�wo��)���o�B�~ӓ���]�s=@8�ߗw�y/	�F@����<j���_v�O���>��mhCڷ� �І6���m�ý���?�w���7�o���j&e�v�,V�h�ܒ4��|dB:���IԨU����0l�����-��������\&5��1���rL��ji���M�$te\$Q�$(6�M�	��  �a//��!���y>��[�$��x4RpAJ3M�d�Yi�'�r�����|����vɧ�jI]��Ãp�[҆���g�����+K<��> �Ӱ}��YUL9�L�;$��CXu}�bJ3����:H$(�DY# ?^ձ�b7$�e�V��%j`;���k}�~�&�U��3 4Q�c� A_VcU�|O/�ﯵ�	b)c�K�WhR%�������2Q�!��*�c�حI
!q���Ɏ���D%)t0��i:���֤W4YƉ�sځB����{e H��n�`4 QG9�0'�*����9��~(���e�Do�/;��8�s��@s։�����3L�f�.���+ǎ�F��YU�_��Mo0����t�M�x|���Is��.�5�p研�j���mi�����|�.B�)�$`P����&� 5�@>��G'�dz:?�X �S��P���^�$f�(���p$���yS���^$n�����K���H�r��9e� R�i/��������݃��B[��C�H��ZH܎����1�o���4iο�t�w$���N�U73'ߪ�
?_uDٮe��p8V�,Rcu�|=(�����*H�˯{q���i�~�?}Wp.yJ�q������1_�KH��TI�7k3`^��|-,	ȯ��ם���yt��*��H,/�
�Cʭ�U���䤦�M���q��= >n������3y���䷟�_|N1�`Da�;���̠,��(�.�ۧ���q�%̜��.b�&`L�`X�6%ip�T5�q�GTi��[�c�w���46��H�Y��iL&	��t&K�Ec~��xU�)���^�9(P=8\֩�դ1C}�p�0�>�?R�sMk�s.�1��ߎ���� �ܱ�<�z�������Y)��]���F�M�x^����GP0��%M����+�U�3���+0�LAG0%J[�0N� ��-��ex�)g�	z���:J�*�G%�
�����g)��"37��>1j�Ă��L��v��&Ԉ�;�3�5� ���<k���#2�2cō%���(�yk MM����'��B��� ���,�>3�vZ-��ێ��l>�ο���dxЋ�$ w��>*�zs܌;ޒ���u��]��%Iv�)!ˣ�"�z'˗'F���zd�+��"�mPb���1�ܟd]�L跁�}G����� F%ۢ�&N*�gl�J҅~9::�~�C�������*�se8�.�)�����}Y�i�lF�1���]�ܽ{'��w�7���~6 �a�{���І6���[� dhC�І���e���n��ʏ~�cy��7X]��h$d�.ЍN$����$��[՞���/d��@�O'��\�g������Y__uߥIӶ�W�����%X�|�V��3�Uo{��&��ZU�؄�X�rӸ����[T����MR��A��y��Z�K=㺲DR#��5�0H���v>�u�b>"Y�v� ��h���d�r���di�w�"�'@II�4Խ\*���uә��&�s�����XA�J�sԼF��J5��d����H�!�FdK����RCt|Gm	�ƀ4�HZ@C)1fn�6�EźJ �Cp�
��J��5�<���{�}�G�֮^�Ԙ~t�!�B�{T��$R\��hB�6	"��t��b�����*a��wdm~���%��P��6�.�c��$K難��/����X��s0�U٩�qz�%��Ğ_��%�<A�7X��,���^���O\2YR�ݘd�UcfH���3�M����K2: �}���V��n�R4	���4C�6�0GB�l/�ϣ�(��|K4Y��e�d'���t\cƒǬ���,��uģ�F��2�(�A�K�
YT�W摲��\l�4��n�ǚ�i�a,O�)�4&0�s�#��1#NT3>�ԇ���&�%~��d�Ս13�}I�=�s2��D�TMA��Õ��׀!*��)q���%�kKQ�-:��k��[A�Ke.����<�4i��׊�u�uzd��B�@&�.`�-���CL����VkY��]�s�L
�15��"��Z���R�k��W���W����&s�s�����;��;��s�<�\���<~�H���<y�T�./h<>��UD�&�JC'��Y�Bv͓��3H �} �2G���$F��C��k��v<�O�j����R���3k�#v\I�c�3)���/y�`�d*!��
=Z&S�a�TЛ	TV��u�/�����"��� :���H����ud�U1�E�q�.�g�݁� �Vʱ�1_D�9�+�#��Q��rx����*��M��╮B�����J�{�@�{S���p ���,T��.���V}� �Um��]��,�2�}���4V�#0�b�0>V��K� bo�}���׆9\5�E���ZAl����w4�XP�@/O#SrZ�o��cHM��..�)��� f�9�d�(�3�tK�~��$����� Y!�	fA�o� �E�6♩.5��s�K���GcL��cj6�K6��G�3�GbeK4����{Sv��Ir㧃��)��dʸ_H�frY9 �\t��}6���Z���%�-��t��5(��2��T�|�ӉL�3��3��������Ĝ�x��+�T�o��0�n߾#?�я�?��_6a��aܿ|�B^�x��Falp���Z\-�MI���$�������e4S:���������t>�8j�U�2XC�І�-o 2��mhC�gӐ�}﮼���a33b~��tH U��t����تڡa�� X/�����l��p||,���ܽwO�?{*/.^��ե�~ I��4l�c�*����>����l��*��qBC��['�az~�B�<z��PM�
5$xQY�t&�c՗��V���*!)���DZ!��v��T���%3_^^H�YC,H��L$�R�MnE3�ܪbSJ`�m~�W�J��,�����A#
x���DHthZ��@�RE#ރتqU���*�Jg A���h�Y�$2�(�Ω�� 1��h�Uy3�NO=?Jh�l�M�B���m���6�w]1��U�eTu�p��Ȓ�$�{�%lQq+����8�X�4�L�)@�l��z�*�U��B��l��u ��n ���P�ޗ��$;�}qq!�����眥ї����'���	��e��oB�����W:�d���~�~���Ā���36�z��t/,p.><ф�sw����]�MY4g�(e��zӠ�zD �|��9�LxU*��L/U�4���R�7��4'nJ��hKj�iY"�rqeU�����eΈ�ՠ[�˟T��C�з��>�FfJMc�VA�#���R��i�3*�#rVC��,�>��Q�I�r���2�B���-��
20�V-w�GJG9>��J�E�q4�1׋%Q�``�n��XɎ����ђiĐ6�S�yK�*��tX�)0Τg�2v�Q�\}���e��b\U˘�����w��X�$ ��y�}�
}���{�B�+���l�|�HGR��4�Q�xWb��������>��� ꐗ��/I�����3��������|� <}Rc�I�?��@�^-[0{ '�u'Ҹ��� �M����!�n ��(��= �7a��r�Μ�B
r�.�B���!��Qϐ`��� ��Y-�f�kd,�

a�*�^�t�`�� !(R���<w�S:I>e���X�Xv}}�י���{h��=��@�O�t�ץ�\���A�~�D�[RRSߋ�S���{J#���07T���u�$��8V�(��e\i,R�'�`E�.�2Kȁm��S�_���e M����������B3��Mt�����G�U��+�l������:�Gע���d~��4��W�,SoN������B�>��������u�A�� �(�+wL���Q=��!��T�`6��4�����XD����e��� Vu���Lf�q�r�
�p��1�v���ޭMdU��ҙ��S�N�pi��0�*qHŝ��ǔ�^D�l�{�V6�h� �	z��9�<�������������|��3\�Y���R��j�s��Ϥ`��!Qrp��ys�Ȇ�M!Қ�ؐ������j���ݽ'o��}t��J~��_�'��V>��3�Z^��=�����+<��_���_��P��_�W���16�V�h��$���d�us"�C�І6�ou�І6���M;�}�~��	c��|v&�~�9�^���ͦ4E���e��d<���z-g��ȃ/>�I�w�zKnݒ��\&�'ZU{����7��:l�А(��_��m��<�����m��h��\��r�VW3�4V�hl�_�_�����0^��o>G�:���Q�
I�%����3��6P�//.d�Y�B��+~l$�.�����K�aey�����B
"��0�F��%�I
V�u��8����T�u��*���q������x�}��D�&u�(M��ӑꌻ���$$6�(�O,Y�RKL,��7b�Y5�䑁�{�h�i�c���V��H�c�9g2��a��ұ>h�
pg�*�
�dI�P�Qr&;F��R�&c��6�=�l�}C(/Rh��+|S�$�Y�K�@g?�hݾ��Nv�y�7K��{:����o��-�^gf I� -L<���~����;��G������u��oԱX�oH�/�������`AR+�
;�Ȁ����K�D��dӓ	�9�ۨ" ª_Y3#�x��(f>
~6`�40�FM+Y-�U�z��h(��)9�V�05�{�-�'�h� ��H5 ~�	�5d}P�Z_!�r������8<�e冼���2(�vMt��"룉;��c�2)j�Ɣ��'���p��F���p��r�$�W2C�=6�	�I�ߘQ�r^��aڽ�^�����qRkU1���>�A�	�N��m�$��-��O���h����,��pǀ�.���'�̃��f��N���vI��/iʜk"��s���3/9R�y���2nR;���['�r�����=��>�^<?�'Oɯ��|�MH�؇���}C�`(�qBU��t�w\!���?˕9���Wեdm�u
���0ÆY�V&��6ה�[\���F��iN���fk��c������&�����?�F�Ěk~��ʔ%�]mUz�o#�cj@������ x��<.�g�9��AR]�E�°�,^*��R�[V�#�� ��v�P�L��O��x~�x��St�<������L�M�IM	0 �\BQ%�
�k�$�5������U�2�q�+�\�>Y\��g��ļ1�n��EPY��.v:�D���*���V`2�w&`A�b�U�<JƲ�K��]��yR�)7�%ASgA�_���5bO��V�u�;�����9]͎�qH�҈�4��J=��ĵB�=���$0�V��8ٚ�bn۪�d*Ʃ,�Y$��?T�����P	����;�)�o(�����d������_㸉GB�~g��9y8��;��a,��9g�ݻ+��筓#M��¼�R�V?�8uqy-/CLG�ӳgr�����T��B�ڴjv�b�@IF�V�J�~��a^���,����/������h!k$<���i�Y,�y��������e����tC	��_�� iC0�O�7��mhCڷ� �І6���E�f�^e��ӧ���?����_��<{��f������&2��d6j{Ӊ,/_��?������Cb�� ��|��ߗ���f�G��Y��z$���@�#��Y��U�i"�R՟NX�)��o�� *sU׸T�b�$���Ϙ�DE7���MUѐ�L�]�����L�F���Ƴ��M�V�K>`��J��Lr5HW�j5����0�t�kC> �ML6*�^��1I��fչn��Xh��a�K:���#�J;\�IX�PaXEZq���f�&i�f 	��E+���I��&lp��}�Xe�쌄��,�.ȄS"�5h#�`��ZͣZ��/�Io��2ŭ�w
6�	5�g7�ȯ��i��P�	�o>�ߟ��|C�5Yծo4���c^��D�8w$'<��f�}m�>�z�}	��K�є���R�A�.�0����5\�����*8��eh�j���O���������J��ui�!��F����	ګ��M6�C�}�?e'��FZ9��ѯ׹J0!)\o�*��.����:Ď���u�V�s�Ǵ�5���ec��
4L�B��U576�}\i
e�м�c�"h;e��1D+�pN��P�:��1�dABߍ���۪��{a��=@:Cy�["�|Vc��<8�V29��v���/ ���:}����TLS�]�2%�L>�7.H�l �E%q+ڿ�J�<ԥ_�q'9@߅��M�F�鈣����-6��r��; �R5����J�_�0�+�N����$�o?a̟�:���ݧ�旗������z��	��}\S���Z�KjƗ C 7�PbK[1��B"���q2e�2�8+�Y@ �
e덓�D� �$KoT����d0���ʱQ.���$����U��;�o˛o��y���Sy�h0,�?E|g�3S � �ID�8�����r���Dǘ�-�����{ry	�D�U����O�S0 J�$� 4���v$��x?�<�^�`����y���qQ�)���� N���p\2q�VY���%A�H�c<�$Q��>�`�c�ó��Xj*Gfq i��tc0�yd7[�*���I9)�>6��_g ��R�&�F�,��n�}IQf��L�7` -׫0�r2���0I�ؤ���VKH������\�5ظر-G��&a�?3��d-�zNG���*�_�V+�gX���Thڽ>�{܀<f�B�c{h�T&�Ք;�H� 8�����K�2nx�8ZR� H���o|���5m:�Rj
 ���>���~zz� *���;����'k-8�"į3���~%���<��3�����V��8��k��Ju��}�E� X�(>��߅��8	��?�����/�`!��񩜞�����ɽ�weo<��_|!���/�s�y��V<x@����H~��?��r��_mx:��p;� �І6�oy ��mhC�?����>bReE���� �W�W���l�FT��d�j�)6�H��\_���O��tl|Q���w�~O����( �6w.��06�ij��(�(�B�B��J�+ZM�'4DN�yl�������ӟc/|gظ�Zю��h<���y�����/dq�rUH��Ѱ�ɓ3nr�$�2���\����C��6�	I)c�����[V��&���'�;��V*ȯ�U��P���$(�R��lb3Gn(��Dg�Ė`\K����7OW���T�����F�qb>��I����S��V�ׁ�����%e�bK�#ɁdI���L�V��-�aĢP�j%��!!!^�&��GY��P<��P�L\NJ�o����?�q�*�C��Qf�4ف/�&�X�I�JvE�3	w��dL����S}sr��hgv���f�\p�^��2pJd �r[} ēy�8 �Rf��f4O���􁰾�4.I�?�$��x�~(.�e	�xgܭM=8XAH��*g�o�2��e*���b��g��c��-�@���A'�28rM6���pC�l���Q�K�UTʎz��&�"�;U���	���L��
��)Y���2-����X�xY�"7��^̄J�-*�0�=/28nŤ[j��J�I-��\��"��� ���pd���v��e�xE���6����a� H�<I��P5.��y��.���z�{a}���5Ԛ\4�|�e��a<�2K�S4�W 
]L/�p!Kƿ���M�!V�1��c=w|�L���w��\�=;�/^���UX�����H=r(��P"�kO��`����%���0��I�$0p� �����X�\)k2	�|��L���h�����8�/�Ym��>.���u�GdkFb��c0&�М����$��6W �`^�V��`�`P��3
C��أ^?iS�6���w�/w���4+�������*1�y,j���b���X��٨�w��[b��oU���>�;��D,��
���:2J��\�	�5%��������6�f�~ �_v'�	�mqu�?���b,��H�m!�i컮�>V�z����#��> �xr}�K��>*2iِ��a7��i����u2N�x`���+�>*k�n��b���U���*c���S׽{�� )���]���pU�Tv�Uϔ�,gqb�.����Ud�IW������/c�&*(�Y�<�ps�^jj��U��V�Ϊ�J���W���-N�����I�]��D����������˭[�:�̡�Wiw��yF�+(^������O� ~��w����������������?��<={B�,���m��MV�FA��sI����t�������$����y�;��D���������>���7-�O����5��*��ex��D�33{��\�n���mhCڷ� �І6���o������kn���z��!u~����`<c�g�Y���%��^˃�?���}*Ϟ>���6cy��9�JL ����as�w��mEZ�k�i�j��d��$/}$\*�*a���]-���c>ߗ�x$���r6�4�m�K\{��qq~����pc�Z�e6��˩j$�P��`>e��/$��q��9�bEߗgj���q؈N'{��BC�h�9�M!���c����P�"@C�,2�*�� ��x��'[��dnL�O��̼&Ȁ,|Rh�^��6 ����d�5K;�إ�>��!�V�g�����#y�-�Ҁ,E�����b7*[T��P*��#�� |� M:k�HdH�7*�RU[J���N�
���|���$��uMq�V���"����J���_�3��<��9 ($	���ĒHn�q��F�NF�u9�U�+⋮z������>@�K���$ �l_e��xx�y��%����C��vHY*8������2������.��3kW�Mt�)�4:��a��L�5u�A Ҳ&a����ѳ#J(�k+T+�����/<y�8D������ $Pٍ����Jzĩr��1�*�?[q)��Y���,M�K�Ś����2I��+��Բ�bK6'�'e�%���*#���Pe�jl�'qw�y�%�}Z37���a��DǦ��!�v)Qgk�8O��{_mrU��w|]A�9W��Q����l�4i���Q�_�H)����pn�lji��L��(}�Ҝ|6���;r��m9>>a��b�Y ¨.��<y~&�/.�`0#�y~q�A,�Md��H
�I����~�q#���'�0����p�M��b@eq~+�H�/�뺱��3�o�Nڐ� �	s3����j�,�=I�MY,�X�#���Ʉ�����9��:���(��|�cl�.o���\�j5w絉��P-B�= �����B��uq�i�=h�;�}���)�sM��@���Vc�LM<[�l�W���n{�+ɯ���(K��\�j�c	��O��,Q��p����e�R�ʫ��X��E�0n^>��0���(6�'���ބs]-c�)C�A��:_�D[l�F%([���TL&�(�(��k#Y��L�X_'��p�]¾��������c���^ٴL��s̆�/��:h� �dxP?#��2����Z *���9�q��fq'A	���|��)�����1[5��'U����9���
1x���{'�U����ۍ�����#�z�Mǲ�wHV���^�{���a���r�ʄ�1�)7#^e�9alcȫa�@��  ���LO�d�ݾ{"'Ǉ���/�A>����{�Y!eV2V�mX�7B6�J0F���D�<5�<¼=�7���*��l:���z_>�·rtpK6�+y�w�8�m�,���Cy��7y^d�^麕iQP���Wt^�6��mhߺ6  C�І6�o�������_��ʿo!q��谙���a��z�����0VT$>��R�z���7��_���_���m�̌�>$r��fL�М_/d>7��٘@G��$QC�Z�&�z~���6�a��ܬ��M��9=>��)C�"��ǲ6�'w��ۘ�f^�$����l�+Vp>~�X=��l��ӳL\Q�$l0O�;�7¦�K���l֑x��3s��9$�!��$�z�`�*�<�927��-^k�L�Է��fr4J{&�;�s��&0��A��*:��)��N�g2I����v�k!�#�	Za���bZX�Y#�̒��B�"Q��F���7+&������4 {����h�^h�h��l,#$��;��2k)��Hk�� ����z�*z��*�����7r!�OY&��������l���q��M U�QF�d$��o��H��!����f2��C�V)����&�64U��	��5�I��')X1%�~~���l�!� ��1ʈP-p�q�,�q�t�+0�h�mI>O�,���;�¥��{	4H�8���/hߒ��O<��cc������q���VbgV��<���S�d�7���M�p-$�>�	-�c��a��&��+������#�3 �p�B�H�8���0��H�i�(AI.5rO�1Z�~�P!^+K9�4�*檁�|8������n�Ԍy�2�&h7嚀�:i���]@M���S*H�S����4�)U���1��O�d�3X&H�V��[]���xE�����G&L���ٽ�k@H�����N��k���%IW�Y����r�Ґ�Ire/`D�%Y!ܣ��5%�x� DX�����?�5�?�dD���~Kf�rp�Ov����[`<\A3��B��WCR���4-G���1E�V��a}�ڦ`i�2���Q�t�ɧ����^�����s���J���I�6����M���M����J���������L�3�;�gO�_��1;�-��-�Z���'3�������
I騡�1�\�-��NCV�405s�	 ^V�3�lF��c@$�0��l�&�ԚԜƻ�V?.�����P�UQu H&��4\�mm��Pc�wi��	$�*3n��*c����jM��1e���-e&ե&�)�ՔL6��L���3X?U�wWW/���s�I�� �O��QN&!}�ºq�<�/}.���^�ғ�����TFa\�qo17�,����Z�+-�����\k�~2�y|M��f��&G��&���<ܤ\t������S~t��n.�}�� �4g1A��������{$�F��K�'���<3B£b2Q�^Q�g
��0.��'��>߀�-6�gx��s�{�&�F�uT��g�ʐ����8B�G���\��qi@3�^�R�#qx�1���4�Wxi|��/$1Ss7�{@O�׫2�Z���1�;�w�����޹��!�'�`�:�<��2����ϑ���rݛS0��!�(B�>�y�ea�³V�E��?����T^���o��~���/����ycT\�9�� ��1����3FD9ڂ�Ư�����ܦ`>����oR���R{�w0yWp4����������|,�39{����E��Hm乕 2��mh��6  C�І6�o�m`p	��Ř�M��a��ޗ���$=v��2C��_������~F,���CYo�Z-��^����.e �Au��&#CY��}��-��\5����=V kU�oԱ	�L2&��8E�qȄ�䩌 91��sb:�3���$G�1�ON���X, s��/M��|��'��₠4�Ϟ=cR��� l�>�O?�L���qc~Jcٹ\��٬���!�H��j�5bb9Պ�H�� ��RK����F�|_��� L����f֜��yzj���������l΄ZmRBH��l�I��c?�V�3����?���3��Z鬆�����V�y�NC�7*��R%���*M FT#��'6SK��yE�����&�c����ku� ���&r1�v�3��v��@9`@VJmi�1�/y�&�>���
��h
�JH��^���������{��"nx���s���cR'��a�_�y�>o�9g�h2S,dδX� ����I��^�M����q�:���7^��{��$�8JӘ��k�XZU{DN��i2G��t[EU4�I��P�G� $h(�A9�$�ݖf�kI鏐3郄�e�_a��خ�z:�\�S�QȾ`,'yLX��4�H�c��9�p�BJDA��ʅr}��;9>!�	}���	�Z�pn�-!����#�pK!݆� ��*��FM�Y�]�R��	�{p��3��X�s�$�T��¯����w5 ��L���'�!K�&{mL���������F�(�P7!�1u2��������L�b�����˗/	6�7�む�H�W���0��0>�Εa|²���&���;����� eP�*V��F2ޗΣ%Vq#�����+iib���Z�-�{��JW�,�ȊB����$�8'1>c�S�gO��D(er��E1 �#��q[��@bb`��/�)�ta��x������J��<���[��G�/�)�s���@�ժ6�;M"路,�jY��}�%�Qx�{�t̸���(d��x�^/���A
�1��Zl�$#=W��ɪT�S� L�X,�sL.ZV�C���Ś����jD��RJ�H��]�%��v�qksi�[`��Ш�@���Dl�Z�����E���s���(<� �B��
t���%�4�o�cXK&ٔ�Hm�ߓ� � ]��1�2jhex���عu�C��z�	��+�4St&38S�R�0��ULyBJ����XC����V�j�m��$�y�){�|u�t�#c�4� ��Q���%7���p��n�5Ivs%1�N�g �Ɯ�iX�c0�	�v��X��Wϡã#��\��G@�>����{��Ͳ�;���Z�ٰ̫D�\%R�4�\�W��!�0��?�1��
EWrVz�& �����Q}Nh�ؤ��)$��V�s�>���5I6���|��ܐ�K�o��Y+��7�zS����X~�ӟ�[o�M���xԆ�������Ԟ|Z�І6���[� dhC�І��6T�#	�������ɿbb	���=���}�M�ru-�����	H�������3����sVc�y�67�����)��G}$?��Yi��@h��=i$��D�ʲm�Ƹ�n��1���a�8l����7�c�+
�?ؗ�lFF|GBYM&�a�v~~�f�{;?T.�c��Q�Lo�Ͻ�
�7�~_�z�;��_�g��V�Ky�̔�w����[���}GN�f�ˇ����;r��X�>}*_|����e�c�M3�= ��7��yh��" ��c����$倐�F�/Ҥ/�#QPU��������M��D1���ʦS��`�H�MR<�%��Y9���U��[�Y�vWG �Ҫj�j�lK&)�DOM ���b��kց~�&�� �F'2A
��˫���3C+{��0I3�5I��X��sSz���T �u3r1�L�k�{nh� 7�m��;���� ���Z�g��)w�'�`.����\�h�w���4��չ
NH��1Z�چ����M�JN����Bn�m�0q �9~������=�nV�w���(t�x�H٪<�?H�$���<�܎!�s�l���S�V�d��-qx�*��Z�r��5*ߘtn5-�1��u�Qƭ���W�єI��f���Ik�~5Q�CX?�0[�`��Z��Q���\R�� >r���� iˊJA���6�]�8 DV���%8ٿ�^���%�^U8�v���Ė%�7����ΥL�`
~Z��$��f�y��;�!�˦&��Sk�8�	)�Y!1b`� �
�sqY��-@H�[a- (��F�4�'''<>�i���gնX�z�2��*�n/Լ��A��Lj��Z��%�d�L����*u�%� 9��R�\�K2wa�M}�w$�k����PvI�#�?�5J���t2"�Q�c�4mxmJ	��Ґ\�a]�s/,mM�멲g�Q��Å�ږ5��(0�u�n��c�2�d��N����/��1�i�*a7��d���D�z�TYǴ����/��Υ�\q��`��49[�`G�	u`Td�eP ��xe�����[0���
l��J7n��tϖ,MgLȢKm=Q�!��t�GY��z$��uw��s���y�@��|��wo�/�{W,X�qr^	y�RV5潂� �X埬w߁kf�~��vJV��1��d�F�җ�>&|��c������(,�Ն�>���&��;3t!.���FYO3��G*�ıjׂc$&u����L�%@�4��*��x�BјW�a��d����f�9�Ֆ��5��!摒�c��-Y��Y.<�,�}J��	�{٨���rʘE���-<�ZH�edRG`��sZ�������s<�����pK�.�PϞ�\}C/����	@��Q���x�O���m��/����Ξȳ�Oe6���eÂ�?�P����ܹ}����e�r��I�3���nxn~_^����ŵ�Wk��EԶ���.�W� �6��mh��6  C�І6�o��|��3;,�R>��s�{��&O�J����} _=��|�����
�}���ջ"lT���HcÓE�|����O~��(l� с�G�uCv ��* �Z�0�ɉyLT*^�^*I�8	/$��!6��%f�o$^��)�6l�F&+Tps9j\��A�2����ᆿ{���ȏ~�Grqq!��������� +He��������7��iz6�%�َJ��Y���4��qݳ�/��� AҠ��iBB���g�[���6���������4�
����F�ML`����!�t�`�[HG���j�%�t��o5������Ɗ����27p,�&L 3���L�����h,!Q�YݼR%�I�q��U ��@��0���F\\o;&��@:@ ;��tD���e���i�Wfr�U�n�NcQ@<!���Ӯ
�6�ﯡ Fҁ}�l9�*S�S��ܿMe�6���v&��Ng���*���A��9�]>�Ǻ9H���}�z���5}
�>$�*J��ט3;)��c�x�O�߼Up{S���s3�6QY*����F}v��_�k���Ն&Ϩl�4�1�p� � ~@��ـ�I)TtÃ'��$ ��HR�&[f�E�d.�l�	�/�6�DO�jl�Y�njL�+e�� ����h����)T��j���;b���Pl��Au��47/��j���L��>Ɖ�H����D��lۜ+�<��GR�8C�I�QN�x.T��;�	�m�K�Xt�zR��!vO�.�z�A��k���^��:�6 M��&A��@.�ј�ց�lΙ��ίR�6��2C�z+�:��^���0�uQQ� 3Oh ������"�l0�K�يZ��%�gaL)c��됊I��Ӗ�R����X���}�!՘�C� zR����ۊ�fa2~Q)�# �K�V ���u�/���H�)%��e%��xJV���p>�M��̈	AZʁ��<��@V��%�{�34��`ִ��9A����\���.��d������U09%�G� $!0�%��S����^����@gŹ'I�z��A��d�V�c>r���;[��i���Q�:���]��X	X;6�J����L~��
�Ox����&�3���m.9�&v���ѢK�� � ݅{E�Hx����I�_w�Hz�:��������zM�-���`�B��Q�)�;\��6� @�	�.<�a΂!�eyW��@��!;��Uvb�R�G���m7ێ�Ա$Q����>�\(�m �k�y����K	NR˙g4��r�M�����u�ļ�n���xׁ��v ��}:�S���r�����b��s��E���	jX��96�_�W�80�@7��Xw�\��&<+Q?J$Ĕ���|�]�*<c����syq.O)��/�����֗��V2���/�Ex	��Ϫ{�@q��J���C9�w_%A1��f�X�͸f��<eL�R�n�/G'Grx���&ˮB?y~��wz|�/´�sz+C�І6�ou ��mhC�7�Jj(S��ٓ��ɓ'�CY�<���}y��w���TΞ��=G�(4՗4ᤁ�zC�$�Q�v��)7C���0�hl�/"3�
�N�! Pa�K$Jau8�a>�sC�D(�����t�VTruq)�́|KEO�q��Iϰa�|�W��A�:�H\Q�c�~��ܾ�|���?�O�r|z"�.~*//^r3rz��Kx�<��\��T�ٌ�UH��@ww��ߛ��7�{�^E~EyM8�����	,V�{��~&&����Gg��6L�QO:�c��wT��U�b�7i�{6$��Lݫ>���@��2!���h\ �k�L�*�K`ԝO	�cP�W�T�_�Xn��U-MWU�X�qW%�� �ƑLɰ�s�4��cK`c�$4����d����Ƅ%��cb�(:٪W��9sēA��s���=~zb�?O�^R���X8�~��ܐ'��&�@�>[�xOd�V+�飲er���oH�5L�!	���Y�o�~H�da�B��  w
�;�'@�$�4������:o�4�V��Q�����E�s�����	�b!y���>vX�H�!�_������:)��(q�2����9��{h �rNЅ	}BP���X�R6 N���Y�z�4��YW*{�����?�8��#$�c)V�s1ً�q˸�(&�t�=&���c��p��1�1��ɕڤ[)#*M�i��F���SR	:�^P�L�~�GU7��Iq�<�5�&!׃į�+��4�����
�b��	���O{�=@ϣ�#�̙xЪz�.�W2���ky��*�U��F�m�����x������y) Ӧ#�s �Xk�&*���j��iD�}�j���"����C����)ML#�8�x� L��\�L&٘��1����"a�b�oU��q��_Ab��V+��=��Kߣ՚ǜ����H�{�ȧWO�`[�8�`z ���g��~#.���ؼK��qT�cRO�Օ�YD@�q*κ��9���O��Ze�܌|4λ����z���@:�H��X^c��I��{A2�_w��(�Q(�F��sý������b���[r������
�9�����q*E\�1pp�(b���x� �D�X;YD`� b �_c�懱g1�O%:M9�j���S�1�s���/wE���w�MO���x�;Iv�ܿ��(���U�h���0FR�7p�%���(�i�m Hn������3��R3٦_��a��m�GGG�c��C�*c��b8b>�/�m�Ճ,I��&~ů$uƈ*{�h�]�s�ށ��`���� �Y
�30)�"��Bn�q��Y�X������a���Ϡ���b����9������.��u��#���� ����/��6��b���&<l�=�J����nסjٟ�OoO����M�ܶ���u���G_���3�u�8��\���+���d<נ��}O2�0��xn��'2=�q6�B��8��x)��H�����՟�w��#�І6��}�� �mhC�о��|��aY�[������NN�oQ*b�`&Ƿ���Sy�E���*-�M*�a!���%*Fᛁ�T�X��
�G�7�ʾ|�����.���������Z��Aj���q�Fko6�[�'��b�8�����V� #QY%j�#A)����kj<=����^�_���Mܜ�ͪ�O>�L�����)?��������&�> ����������r���b#�G�2��d� �)��Al����BQ+�ݵ��T�:�as9$���ql?<��� �~3H}��ْ,�u%�}��sμ�fխ� �(� �)3u���O�G��I�'���5�6�Y7	
��`"� Y@���ys���G��9qA�3h@����C����s���^k� ����zYN��<Ѷ�)���G!�V�	T�z�	�)-�zR�	�E�X�_��n��'5�9���\ ��$j+��OZ["�K\b���H!�����j��k&I��iM�}��$��~�2��,I��Kd�b��B���/�䥫<��+�=�������$����!Vú{ᥱv��QI�+��ģ1���23��J�J�x.3��J]���VL�<8��;�#�ycɭ����5�L�������K��s����Y
}�+�hC�=�Ł�m2&�;�%P��`x����ѡd]����sU6��
C"���A��u�i���I��5a`2/ \�z�A2S� -T�L���ǹ0��X��!�$D��HV�ǛuE)��*����4B��1/Z�_�~�8�L���Xr0L�M�
�R~n���5�vc�l���(
�U��������:}+�I�d_܍�x�t\�o�����22��Hu�8]&�5��76��1��(��s��2H!��1F���-��iί���0%+�{I_&#]z��y/^}��Xl/��<{��LC !u�I��)ǌo�$ B�ƿ�
��Y����������Fo"aw�a�3П���Fl��@�z�r��~� C���!|j�tIِ�	f�'æ����5}�)����e�EC?tH�$�z�d<ֆ�(Y�q��{�V�b��T�%�� A��)U�^͍m�:������y?��^__�xX�����5c/��� � [nZI*�<ñv�< �c">�3����c1��-�����K]K�o\";ۘ�5Ào�]�V�|��7�.���"��$ݾ�����g2յE] ����M��i�ћRT&�5�/��n&'����d`�w((���m���v�Q��gQ�p����� �b�W�F�8�X�Sν|�ǂ�X��;��3 ��Y[�!<���� 7 üje��ߖoe+m�z������0w�.x�wIb����\����e�8��m��/�a�l�z�B�v�4Ҽ��ۚ�k��8q�;��0��K|�?�k����DNZ�}���(M�)zY�q��¼�4���~z����]\;I���o�(9F����R�[1��/�1�&��<� ##�^9�M�� Ȱ�8Z��ql)��с�|dO�D�s���Ͻc���X�;��46�e�c�w����S�A���0�qIiL�g�CxV���2�y�������_IW�c�?{!?���o~�w?%��{��N~��hӄ�^�j��m�����}۷}۷}��6f���f�����#��O&���ߤ����s	��F�Gc�ȕ�!��
O��L��8؟�rttH�@7���W����?��|��2��1y �ߍn�P�	3l3\f��4.!8H�2�c�X	r���	�2��\�uW�Z��
�Ќ�#'����]� �X&�MJ�fёR~���~�⅌t�x���|����>��W����gRl*9=<�$����8P:���(�C�J`�	��Nǒ�lr^qFԬG��6z��9A�&PZ�H+Y��Nr��n�?`V��=�z�����0R�Ue�����ك^�A��	�p����=�{�D�[�a' ����w*S%]�3����6&!T�`�U�!�a)�F�w&+H� 0sռH��z]�v�@��]%)Q�5���$_<���	8�]�S����7���ˆ�-H���@	_��z�@���Bb����������g�O=������rZ�����\��\G���
�����vIK�g��YiIc�/��jerP^*��Śf�^3|��$:9�4��qR��q1w1�!9WTV]nJ<5�V1)���<���߁1���8�������<�k�˲�Ը�� �P���H*���(�_ A�a����%�\����ڱ��p
�P�6a�XQ}ǊA⮨�B�4�1�#�a
��NB	�nR�"��^��0��K�'���X�)��E:z��-Y1�U���GI�靖�֎@K��)��J k��@b�c�Hh�t������$��v@J��TN�G�Ӹ���4��+�n_���p2!���l�j���֧��e��y:7��� ������������TkJb�VMHp���F	*z��Ar�� ��xҘ���RS���
	#ğ�`�#|&s�z�:�0v��A�1��%z E��Y�Tdǒ�um�[�7�ossL�%���I��=Vl#��X��P4��5LD�+�������6g0�0�p�����$T=�{�vI��������y���D&����C���ϵ�������#��c�9�F�xA�N'p�}�YXb�1>�]`���S�2|,��}�������*�/%��qp} ��1A�~�m�	=�m`�����ra�]�Og�2��B�-�������R�	�bҧ���%�����0���&ȣc0X�E�d�,�%��	����lm"U�۱z�QF��1�����^������?�;��U��K1@#�2Y�y��_'�3�=��h��D=�e�B+Z�I,[��GIR�����_b}�{��������]�g��0���(�A�$ʪ�E���~_�6I8�1��،�+��"N���?���Ue�I|F;2X���x�4�deD�b�|q�q�G�֤c����yn�c�����Ф��ɫQ�*)�N��a�aR D���#�u�홍��c���E#G�\KБ����Z-%f�C�0�$ʜm,��b�oEXʕ>���?�5X��yo�y�?�,}�t��ͦ2׽�b>�>�D���,7�������C����X���?��,��7ߪ�<������0�۾�۾��ox� ��o��o��ko���1Y��W_~.�/�e>��W^�/��-��E3CłU��<������֫�|����諯%~��G}$?���W���ϹY���Zw]@�i�M
�R�K�VE:�(�b	۠MP�xq�JŲ���1[&��<L��w��Z1dYl���ek�t ��[\�\7p�zI�]l(�{�=��w����!��7O?��J_�	�h�2ho斌�  7�f�!�������и��6�Qز?��8`H(򕓔�p�A�5`�Z�$�O���� ��͵�m�a��L��.|�lGCo��X�86�J�5��Ш�m�(e��Z��_���	���Þ��b�7�x�(���#Te�jZ��U�H�����H�4a�e-��ѣ�UF0�*VW���!� ��&�h�d�����ǘ2m��s�ֿIB�H�{�̕��B��}=v5���y��Wv���&l|�?��6Q���[�0|����L!��H׹\�-��+��=�}�Hߗ��)����*��ЀU����ss�-��u]
�M��ڪ}g�v�ʍWK��4�G\�sK�!)u|rFɭ�t�D7�.b�P?�C���|P�Γ±dp��߬2�D���|ԑ$��X��X�֞k��@z�q	����uV��+��=���A�:�!B0d⩬�){�I�1�EF%WT��V���Vy�D�_PhI��6���p$��b�2��9����ɻ`&�.�I`Ud�`������T�t��P+��8'K'�遆��I�r<�d�H7F�UǮ�u�ҋJV�G��a�|Ø������80���c`D`�f���F��� qK $�м�d�t|A^l�I�2䢐|�Z�,킬X��zH@� @�F�vc@��Ч��阔XD���^栎�b�1�]K�2VY<��C���V�q����FF`,��[ϧ�%+��Z���8t�+���q	����jk �.B5:
"0�ԁ]1M��4n�&\�U�d�z��'��y��+���gfp,f6^7�[�6A�8m�丘g_a�X� �.��㔱:��3v�m�>����S��D�1�|��5��iYz�Jc�Pv𙁯Dc�g�j��u�5���T���7)����_�ǟ~*O�=��;�a7 �P�e�����c�m�މyB�X������,���$���I�u�x�[*2�pL H��y�����Ve��d� �&[f�_O�O�� E���
�t�_9b+�z�Nucٸ5�>k�j�1�c����3^+��ҷ�|��PvM,�5.Gn����g�3
��2�cE Ǯ�{Q���C�fl�����1�\9��?��|�W���9���ah�_�3 �qo�_�q ������+�����>w�ɸ��n_��b6�x}},=/��07/+��a��x�6C���0N�ÃX7����>�#��'2��Y�s�b9�zRW1�˖�C�'0s�@T���gO���������>=���R�`X?y��Ϗ�s�c�t�v����3�ǟ�Bf�%A��"k�& �[��]�O����d�r�ξ�۾�۾�F�= �o��o��o�ކ"�\�Z6͊��H�<y�H��?�'��0!�T77H�,F#��ml� �����X�d�e����>���뿤�O~�w�~��t�Q�fD�Єr 	�m�@�q��w�DFc�$Yi������Mj�|��1�$W��p� �D X�����ME�t$�>�Z7�9�I��v.�ɀ�T�G�Iќ����ũ��+?�ɏ�?��� _}�+�`���r}s��D��ri�ec��m�����4Hh$n��}I�����hDG/�>����Y��"
�ۄɔ�I'�ECrԥ׮��~m G��)��@��`��_���ε��5��1��@_}I���wG�/�> �NOO	2��24�{$����1X[[�&�' &$# �E���;HBI�=&��9G����X;.!�D��ɥ2��߁���:��A��5���8��Ċ�G$�����.��6��D�'�v%��9�O��Wٞ�73G����_�.o~�_듍��A�P�V=���׽�1���c�����Br	IT��Ο&+�#߳�Q�� ���0���d��HXt6�s�ޖ�	��9�LèG)�g H�-Ws�V���XǍޗ�Z��z��x�t e��%��z�;����f56jy�D�X��J?�3�=�\p>�^�y5��r"���.�� ��ŘD��:���IB	�s"���,�ȃlV�[�p<��h�CF $�x\�O����Fj=��>z�1�����1�2΁4N%��� �5�1���.tN͖ _���5�.*�������?9�*&q> W�B�����V��X/�Z��}Ș�a:H��	�� .כ5%������4�9�+�A�:��x�A�d0@ 
�8f�iO:���c�;��^z�cAo�����"�Ybq�M��Ք�D70Ɏ�CB�qve�G#|�ƀ�l�)E�N����O:���!�8FJz�@.�@��l�f��T_?��p �٠dZ߿���H��:^�0NhƎ��1�S֪�ɤ+	��ځ���	i�cH���h��lʍ~~G��~ lmt�pM��P���%�ipO!��>Y��`kD&�$�F��y����@%k(���
�5xl�M{9;9d\(�<}�ّ���L��(���#�a�C�%j�齫�% �~ǭiM�����.(@?���>�{9��hL9���ܙbw�	�P�:�c르5Z�)��,p,82�B3��̧3�Ǜo<�W^�?��C��?�3��}��G�v�'��L��z���M(�	����X�����,�Ū`�󀲿>�~
T����x4���m���m�d�F�lw�Ó����ј kg�a��;�~��e2F���䜜QzbR�Un�PA�J�0b�t>e�9fKW�q����Bj�N��<�"�cA��46�q�=ְMaς`y�-V���˅�v�b|Ṍ`Cb~jf&Qf
>",4�$`�2Z���3Α�HԶ�O,;@��� ١�X?VB�P�+�� y|V��� B%���cv��e�se�kb���>|$G:�n^�>۳���Xg0>�pn5�GX ���Jc;� 	k�` ?�����=��yz����X�̘ϹX�7�dr;�b�J��w��P���j
ɦ�������T^y���]��e4��s��y�`~OSy��<~��>����7�t���������w��\]=�F�ב5a�'��
�}۷}۷}��m{ d��m��m�~�m+��a��6�����������J���,tӉ�6��rMiʺP�&���I�L�=}*?���q��˯��յ8�'�%��;	��,�&��}���g�p���`N��[B�	�,' �Ĺl��8�q����`Kr���eI��8>c��ծ%H�/$��Vu"!�\dr�`"�'����\����oy��+Y�7�@:d"� 0C` i���EE���
"V}�Z���D:PO�(�j�����Wa�]8�@��%�+�A�v�%38'Cı|�?	��u��E��b@k�˝����.��7����7�\r}���Y揞q,����)�R|ep�>���|�{��&����z�����^�ᨴ�
6a6��Iת�Y�^m�� f=%p����ӎ��|��3?(e�z`횝�д~ �:o�*floc��Ua�{cr�9W��uH�x}|����~VҺ����0}~�����8_\��I�]I-�Z��`�g����? 2�ݒ��ex4��j���T�_떉���<�7��+D�<��1��e�YJ�s0"�Q�� ��rծ B��$k p�M,�9Q�s
�܈�U�� s�$��RC�9Bɴ2���:'֋ad?��H��0p�5��0���$�ge`�!��8�i�o���SIq���S3^7+jSA�~�8>�b�$��`���l�� ��	D�MnJr`�l�����ډ�n qt�|���E�H6�#7ix�}��8�d�,�`ܻBe�~f�XŴ��	���c�Dx6Q��Z�@%3f1<��̃,�X�t&G�i�N�y����/E�If�b����:����	��`��AB�~ i4�����i9֕55�s���0u�3jc�	�����/�4}x�� NV��rzS����&UTر(�� o�����Hߋ���4��d��1	3��[[�:�p"�W��\F} }�Sw���ޣ!��J:�@�rf�/G;Ҁ��kZ��~j4&�j�Ƭ�^�'p�ql`Y�����r����k�=b�R:a!g�#��8�W.���:�-���1�[����E��008l�k��]ߜĕ�7����@���}��F�^�����>�VV��Lm(�"��_�m:
@��;�ǔ�|��7�Z���y������ڼ@,^<�3�GqG�k ��,�<�%p��,|����:��R�_ǳ��@���Qm&��>?m�V1VW�K�W������j�o�Ȏ��ceD��ǃ��$�5���T��y���\/H�{�DX��B<�ohG��/�='�c��մ�	`�m%埌?��z��#2�/0�2@�n7�l���-`$;�W� �W� ��y��}J26��^P�@c��><A�+,@�:O�l�2&&�y��Yט*Q+-���{��d@q�x&� ���9g2} њA@��`���#x��)�<l�3�8F���_}U��� ������ٙ�11�N�+�1=h<�W����\6�5�3F���zy���G g�?��ʪ��i��j�^|�|�� ٷ}۷}�-h{ d��m��m�~�v�������A����l&�ЌkQ}��\��|Z���
�B3�
����$���8��ؠ���I� C�Ê1`�%��w���x���KI�8�J�릖�݊�H\@ڄ�N�P��vZ)$0� o����� 	�����:��+��<�n ���'VЇ%�c��4�}���r��!�?������}N�����I�Z�gT�G
;ST��2cV �J�c	�j�ҘH�|@�|~(��� c�>�8E���wfX^Y�7�F�.)�3$p��x���5�D�|Q��F���	�T�W
ӔǹRbd�2�%�%�����m�	D����i��Ԭ,A&�!��@e( ���B��J���D0�0K>�#$M���P��Ǥ
CHT�q�&�J��`��n��V&� B�����n=<,����2D��{�����<��������w�"�������>y��욣{O�u�jxK`BJ��<�dVyݵ�
��д�=�A�9<�����{$(�z����#���]�+����]���G���JSed�t��O��T��UT��B�,��W�������WHLaL�ږ���n̅8�ھ�v�z�JR�{)�$�T7��I@�$z$D�Ӂ^���s3����L�wQ���7a�nf߇�>�q��1����<��R�`"lX5����_�u�`��dQ4��<B!�0[�΁�%s�)�2rfȹUzofd_D����s�g����'2_@�j�����q �! ���Al��{�@⧒���U�`@6�I�Z\�I��~�hd^�by�n�"9���t��YТ�\�Z*�5�`�
��ז���`)�Ѳ�X7�%8c��2�?:�3@����Pɾ/���Ѣ\����Ș=�v&���)e���[���c�ڷ]=��fʤiB���� ΪT2��\?�1;$���d� C�`�+���%A��!�y��t���z���:D�z����u7�I�_K'0�,&NK�L�=�
��'�nRl��n1��+y�B�Qg��?f�<X>H��#��Tb�T�AҴ�2 t q	��ɘ�E�p3��L���t��v�2 db����wޛ���i��/()���ou�ق�ޏ 6�oـ0����u��hk���⋥�Gc2Q��������<�����_nn��W�����Gq1>B>ւ��q���e�Pj�]G�R��a䘭ng�Dp	s��$i`]����	���!�����$u����>O�h�C[�#�z"��H��A� )sWȁs�8�/�O�6����Iy�8E�1�D9�гg;Ĩ�<�i:��<��X�|�i|�u~���'�������VA��WsN��G��/�U;�i���[�X%�+�y|���A6"��ll���t���b��31�8p>�c����N�dl�H��L�1X0�B�=8��rJ�؉X#dgh��1����!��蜯�����.`0V�l�%�� ���uyyI	��|�rt|*+}�����5۳C��9O�jX��8>�Ek�����"(������y�g���k/�^�����|&��o��o���� Ⱦ�۾�۾��hLR�Ɍ�!���3Z{�I@��'%h��k�-�K���]'�3��X�����M��<J�Y�>Đ̀�4�S����$˃����m�r�le��I�d��r����U���I_x�89X���3&������e2wC�l�����N�{�$a����c��?�y��住>����O���#}�BVn㍍�i�'up����DaL�Й�W�7����?x�������hd͗ê�j��dO:܄���\�n�MHp���Sm�l�їH��%c��l4���Mʑ��/V(Bn�]% �	$�!������%с%B,y�0qB�W���#�Q�qc���z��5�B!5v�X�d���B3��_M�%�����'-p d�I���Ǵ`5�K�y�*�{$���b��%S$rl)"��k�R��U�V5�+v$��V�������5�}��R�I�X��O���X� �gv��bs�]c��dE�<���Nv��$`� E��7hA4�!/C�m�
��b��� *^���o�A:Hf�\�n(��B6,5SV��CҮ6��%&f���+Pe]���KqӠ��J���,����t��z=��pm�#4�ח��	���~��s<e Q��i#P�$]W����\_�K��:u�M7����	���c/���)����Y�o�����,�D���ӑ�i�n@�	L�	��z]��<�s��TAHa�0Ȧـ�1]m��G�%�-3�<[H�s����pȾ�dK�����H]��r/��=�9���)��ZH���	��y���p`,I��V�>�5?��̕��W����z�K
&_dl�:����1�KS,ב���nz� |A�1����׬�NC!�18�ba`s�X|�Ж)��#r�7���LC�c�>�7�Pf�%��]G0�@��9el")��ҫ�d����p���w73yR`ԉ��rpؗ��!��V�m �g�@]��&�����^W��D�䳯�4���lV��qyrv,'��1��냕�����X�"=� �Z�($`)	�:0�=��Uܘ�Zvum����m���K[f�Ŗ�����]Bx�3�|��g��4�K ��&����!������ Z���b�l=����+�����@^}��\ܿ�o~��{�O���d9�����qs}-�׷:W �1�����6[��l��b�Y�I%���=[5�ge�k)1����& m&��&۴e���P	}?��O��f4�g��� 6�hI0��g�$�g���Ka,���l����,�bU��� ��]柁���� 
bv��=C�㩶���A�}`�h�_W4F�$�뽏�y��'�I����� `�~����h�=�ڜW�_�\gh��"���%�S�r@�	�����T�`�s˫��V`il�Yѐ�K���`� k�^k����B�㪒��2�"���(r��c@Zp��g�����{��c>{�u��u�L�'ڟ�<���g+JD��56�3�~(�G�`����z�`��s�$v�d8�IwvC�YUl�������������?�u��۾�۾��oE� ��o��o��/�MFC&�~��5h��	����EMy�	1-��0�#n@󥼸����c�xe��+iڛ�!F�r$L���\���?�k!�����ɱ\�����17��yEP" ����$�wu�6����n�����f��9�U�7f���u��M`RФǵ q�����'''�؃�O;�MO��o~K���ߕw�}��<��?����JC��H�`.�.|�̲�ӄF��|)�|-�n��x=b��*%�1h���y��N:������;`J�|=jo�]Y��(&�P3yPAB�l��-V���)<�����T��ѿt�y!q		��#V�Ɣ�B����cPNx�f���/]��&rրZ9MnT�S���]R�$�
�
z�Y�dE.�:�H
��؁5��'b`t�gHB��ٖ9Q���n�E�.�1��J�U.�/^�K��ğ7�51�����˾��a��`����e�xI*���0B|��K-;L/I���d�_H��ܬ)����<x�5�w�· HDuT�������x�<{�XV�;�ήe���^l>$�i�3�璴I�J��g҈L z�ڂ�K�c|1A�صҹ�l$��B�� ~qB��ʤ�c'(2�y�'�P�t+2�a!UT1� і��lKF#�����Dil}��F�+�T+�1�w]	S�:����ϻ�[#	��x+�@c�i�p�(�Z�������	��(}o9VNյh8@1����J��MN�vzg ���C\Wl,�^3�����?��-���� Ki�2P"��]�����Z���v*+���Ȏ����L��&�E�d\����\�%�����7I5�$Zg�5�=�lSO�Y�uB�e��T5�
���/4�or똬e��쭝w��!�w�C}�(��MF"����/�;�7]]��?��<�)���.N����:�!�j|�-�r�ҵ��}Y�HM�G*ȗ�����:����k������/���tN�O���Xerԓ��� %����}�.u\t'��c���އK9>��1�%��ِ�l�di��*2Y-���bC�����Ae���/@�6�ƭ��+J踸���1jM��֠h���<$t߂�u�=���~�1�%���1�*Xs=w�>|6�"vXu�yDn�E,3پZ������S�21!������Wz?o��O֔p�e-f��/��W�ٯЛI���C��I�x@ǟ?	y!���߅�=���]#d�,!�U'1|�*��un����JXկ�v��!z��b\��������|�u,<�xy)4�c��]��`�P����ڱt�Y������80w!E
�E6��v;/��z�tp��Cb�-�pk�P�׉y\y��]����r�\�{�?8�KQۇ��~y�C�T/�Zn�?�	RP�S��j�I	�9<��-�3Zm�onY��d"�C�"L�J(�W9�6 �8޽�JL�y�K��w���X��W��cPU[�9��u�Yi��6�m�F�]� �'��'��:
�F�ł@X�`���xM��:�%�%&7��Y6|^V�8�kW�Q�a���� ��#z���j��v�����}۷}۷}��h{ d��m��m��E����n�S���% RV�f���%�a4L����h%�s n0���I���@��.��`Z:��H�?����{�������c9??��'g�� ǖ@��@�#Y�&��8�R	�(����H�mu�����|`��%�-��jV��=���$��= �pz���$D���ߧ����OK���Xɵ�t����g���W�KD0��W&�Ӛ�[F��u�iȀ��T1+@��}�`K韪�cCD��3��ם�����ޘ�JD��L^
}�X2]��?� ������C��VA�9!�jT��H��RK��)�*M�c���Ǒ�Ǡ��Q���p76�%��������{Ml�K��U)#��8����p��ol��%J;�M���;����L�c�[����d+���[p�K�x`��xx0�WX�N����5�k��ᓋ�U�~>�s��IP��wv�}[�[��`k�z=�s�g@�����18y��I�(���R:gr~:��΋�d6Me�MARk�� '[�<�tRz+��+���:6�P� *�뒘U�Ww��|}�y�Jw$���t���IJ��j�ыf����t��b�J�2��4���,�f���7[/����&L�E�Tx���X�r�\7�Dfd����\F��+�Z �`=��� �s�\IV�5V��M��QI����T�.ǆYb���D�z�؁��@���׃�t�S�%���P��R�/�_
�C�0P����29<�k��b]˳���x1�媒���Ư�z)��g2�w��s]W��R����F�H�{�H�ߗ�˛Hn�\�,	�狜�8���0���̽�j5����Nt�0q�턲�{����ܿH��d@ ���������L�<�Z�X�A^��}����}���:�$��l�����f2���y��w���P��@��P�z���7����:�4ށ!�Z˳'�dz������k29>�
�7+Y�<��ށ�ry�_ǔuQ�z~#/���nn����H�q%���%�i�&���� 5���9<�$[�	 `�9��\��X?sq���	�n�!�$�B�u;�1�
�G?`���E�O�m�Y�~�M���>�N3���;�kv=?<��N�� Y����k��A��?+�[ �����w8��֤l����O5��X!�O�rxp(��_��}�{��񗲘��ӯ�p�Ww�\3���� � 1d�?>v<��dB�ym@.���ʅ��� Y8�����V`?E��8l�q�G�C�1R8O����`h��k�X�0 7����;� ��K�u@)E� x��M�ͼ���&�_ظ"���e�(J��L�WU�AFM�k�����ڑ���y`�<ר}��y�]�= «���ُѯZ��ʘ݂Ax-��dz]���w]��(b��e�"���T�Z?���W����}>�w��7��g�#%@�_��k���<z��1u�@( X�3>���(���'�?�Ս>����9�y����ٝ<��(A��s}��#���/�@�|qϿ�23�:�q\ӆ `���k,O	6���P{'�c��[X���_�������o��o����� Ⱦ�۾�۾��ii̍?6����������NJH��F��?Iٔ�������F/�|�@�E.��.�i��wO7<�C�����
���H7w�v_Ϧ���c9;>���J?��QG�^�ߙ�L0�*�f[y�N׼"h���)Y5�ez{�c��O�M>�������ْFڐ�
�4�r�{b�ҩ�Uӫ�R7��|�ߐ���ߗ_��s������j���N�KYy�4�e�1����� �apw:�궎���dil%� e�J=�'����D � ���܈Wl�Ʉ����k:�z���S���y�zn,Ԕ�@�1+�C0yRV���F��W�XA�>6�X��#�Q6�$�a�\G�-��Hu<z}�G�K.t��$��:"�+k�"��.�e#Y�i}>|2�'C����eix�O�������x�m��/vY���������y׀�˾��f�"Z�/CE ��Z�r��KzF�7H����c�Lm[���!lh�{��ҁ?8Kf��{{-H�DQ� �+eC���I"$��~�&A)��PG�2���H�e�Z�K�Z[�*탑������վk���\���N�/Q V��C��\�E��2��)Mu4�h�la7`l��P����x�jL�D8*c����񚙳���"c�T%rrܧdH>�qY�1��$z�\��=�SB��`.֛J����������5�2-/�%[������C�|M�.�S�Lh���ԥ�qrP�� �%����B����ӾԾ^,^HU��S)�+K��{��y����$��#���<��X�yf2Q�I"���r��D^}e$��ΡHv �r*O?�X�յ��D��Q�u��������j��r)��J����{O�z�OCI�";ݱ|��K��5V�ҵ&쏠j�[�����׎LF�� �7��H
���뻩��z����y�~_�;d�m���Jnu���	Ա�Uz?��l�/�����_o˽���t%��VXߖW��iL�������rzq A�A�dK�u�����;�+oݓz~-�)�m)R 0Z��G����J���~��R�<�)��z=����ݗ���'�Rh���@^��kZnm�8b@D(�]+P� ������&t�)M:/=�c��B�8�P�0�x	>�H���>n�J���F��X�9��ҙ]{��n���=��kȮ�W�Y�{��z:�����
v��B>��c�5����+�gg�>K�����<��y��	�쐆�v�E$���:����z�Zi�,Mg��	pE'��q�E�u$�t�w�m`� Q�zI��W@<��ֱ;ǐ�`r-K�$C$��1%�2SQ@94[�0].<.�@d�=@zL���=_p�8�1l@�*��|z"�"2��.��<]"�.���~x�7G7���?�y�D��m��Y��#���+�1�~bN� <�	�3$ۯ5�����PI&.F�Nk�����K�w�ܼY�_!	��[oʫ�=�u���t��s��ݔ`�ykU�����Y�+Ƙ���ۄ�HO��Y�F':�!��$[�����~�_�ًk]Gdt@���(�<|49�xvN��L�Ҫ_ R����v�0[-��:���_���g���{��0�Rٷ}۷}۷ߊ�@�m��m������(�A["��>�W𥛹謞e���l��\7L��C����3f��NR�C݄�p_����#��$>���[n�?��K����bC6B%�x���(���n2�0�aX��[�����H&���B�c��A2 �=>=�o}�[�`~��'��������Շ�n�������\fwsIө��T��n�.)SQ~��
�&ҍL�Xod����MRQ�	 �!��f�f �RA`&�S���A�(Wk홸�A���N�26�4���8Hb1����	mJf��%EB�K��G��sjF�)�g{4.!A�� ���2�92 ��^�-r~ �\�9�o̐&0Тvf�I'4? j5t���Q�L�S�i�H��2X����x�}�/�//��]�x�8��i���XFRn��;b��NR���i�l_��V���n��ڿu^�\���='�右۷��sڑ|�% H2x
�������?�A��R���~�k����Dw���e��k��`�q�$�uA��_�w��}b̬��3���u�2���ϙH�u':�J�Y�K1���pByJݡ?�.�Z���4̳5>�_�y.t��_+�
���X��H���|y~$��)t<��������1���W���DC��G����ok{���O��X�~���f3�m��"wk㇩��_ț�=�{'���������e��,^��Կ������2�}$WO?�l9��`��ٗ�gz\�^XP\��o���=��j)7�C)�C�L����qW��Z���,o�IP��H�asa�Zę%.��G��;��KL�h�1N㨞��ǒB�k�K�=��0ױ�¿"d�}�8�:L�	�5+�_<���k��9�Ld���j���`�\K��"�;3ѻ�:�4���J�M���r�Tx0?��ޛ���8��7����ǨW  ��IDATy��3�<����qs0J�xr,��.�ۣ`��m!拢CD�Ke1����J��r��Xx��Ƀ�D��&����6:�6�����j��>13��Wy8�	��X��l�\��^kOo�l!��#��}%����H:�X�wu�UH@�{D�y��5xFp&�
����������%�.e8�)}��u�5	�CE��ω�??�1rO���� ���R�z�6���D_�߃���X�[� (�~I1� L�&�� ���E�rP��J�]��g����������M>�{@{���t1��H��!X� %��`ƘwG͊~��um��Ï�����{2��e|| ������9�n#L�a}z|"#�3({�%���3 J�.*| &!%�g/+/�d~8?�U0�F�ը���5���I�*�|���!�f����B�������e;�zX�b�Gy�a��M�����{v��=}��Kk���2�ɘב���ݳ����S[��x�'͖I�g!��F��Z��n�l�R웨%�:�l��l9��!�	V�IX��9	i�\�R'2ٮ�v~4QH6��t��8����<��X�3:��s�ϯ)h�+ӵ-�/Ȁ'����:����l6�gZ��t{��~�(��p=0E}��ߑY� +�����/Ϟ=��1 ����t�$l_y�Q�.��	,BxU��I024ɻ�>���g�現���G7�_������ɷ��ٷ}۷}۷ߊ�@�m��m���_Dk�.+��n��q�o6�`bEh��K�� ��ķ���陜��ʉ~a�y��z�d���_�7�zC^y����2Q�?��n��U�fYPZ&�M���Pz�.e  ���U��^��O���r�!5l�2��x4���{:|��n��+�g����}R�#$y�b�8�GФ�Q-3�)M3� Fۺ�}������Jz��h����*��A<Ĥ���rzx�d���ؠ�.|��<JƬ�����$$^&�\���t���'� ���tf�`�4N���yu�� L6+ �����8L����<P՚S�ߒz>N��o<ZҫB����  �:2f��S^�����T$6��4���$�S�y��m�/H�a�L�Ck���yM�H(@'�7Pw����C�	���	 �:!i_7[�&��f���F�әl\�8��穁{
� ����z��o��/���qw]2γwBO�i�8��Xa� ����u�<X;ɶ�KRQH�al{O�3����:�$�7��� ��� �U������B�l������k͆q���'���$�K>��t>w����6��k��ܙXK��������0��C��T�~�J_3%�5AVZ�(�L0�p�`;�
���J�ӧ:^_H�|"�2�X��ɫ`�\�ۗ��k��Oɡ��o��PN2}�D>��}i�Q���'����k��,���D�.B���	�P?���sI�F�{�]y�w��異Z��c���䣏)!uy6�����wy�7����tu,��Ʀ��%٬��T�q���$������0���=IG�#Ó�ʙ�z��T��T�/tll*�ge��rz����J�w�x�J�b%��s9�A
+%e�;�
~>K��V��5��$Ԫ���������[y�\�a$x:�8�!d��J�Օ�dKɆ��']6ß���L�B�������t-/^�,gK5��q����n��?���˻��ܽ���j�xst,r����Ih�>���~�B�:|:�"a60N|]]=���;���f�g�HA2,f�/�7��Hpo6k��r�ۗ�|!�����sCc�,�<���o�i����|ip����P��Ѡ�iQ&���>�5:H�ł0���]���=W�f��g�k9t	)���(�2׹��k�Ef�Fח�Ռ��]������YdkJNt�c%��N����4歏+^����e M���1l�ܭ���T�gZ��tL��q'_r���U]q�|�}��/����#v��[׍=` �� xFD�aRY�"q��q��	�b�,�Dd)dl`��3@�w5d<+]�7HT��f�������D��t}��鹼��;��+��O�����١�}��8�-��O6� ���J��ƀ~]2k��X�i{@'܁|��'/5.n�V|I;�[zW�ʭ�s*��Uds�3r�r��`�}���[?*>��0;%�Ș(��Q\2N�L�9�p����q��&���yV��M/���7=fX<P�s��I]/�d!�9ɒ�����{`%tred���|HS:yQZ��&�W9���ޘG|e�य���(q�O��ɲ�e�OX?��� ���d�� ��И�J#�%��<Iοr�����gg:�ul��P�8�^a�c̢@ϰ��1�cA��!�k������1H{dr h ���&�=�a���wMj�Xww7��~ �ÑL�3Ɩ�f&�Jc��Z�_?�k�1��5�,�0�$�$2\�c ��s�}q-�~����G?�|��_&ϟ>�޻8~��wO~���_�����������ɾ�۾�۾�F�= �o��o��o���hݎ��A D�2�%��������\�>����G�J��1����~"�D	=��އ���CR)�O��6M��Ć���3$3=[�$�,q��&(Xi��v��9�.�� 4�Z�,ր�;<<f��6l�k�p�L����0�P}��L6�Vr���Ar���dMz�X7w]Y�u��=0?�
�;]�R|N��ЮTJ:Q��J�'B�>Umf��=Be/�GJg&��"�sKT�S��$�K�u��*�?������UMVu[mٚ�Nb!���M�i� #��K o%��D��b�G	�\�Mn�c�G�JR7uL#Rx�T0�kb3
%�$6�,o�LY'��D6�LڇVM�~_;��nڣ�06�H6.6�7��L"xv����I4i��Pf�9������K��V!{�V��%7<�&�'mu�O��3�t�xE�}�l�n��X��I>���_�iⓙ�ي���de� �x��v4�����@���m�
`���'/= ���c��g�K�ދ`��BF
��q���������{��#���5���
�0�{�9֓��"*e=-u<�dz}%�N��{o�;�.�����S�JW�P�λ���qO^}�B���~ ����0��H?�N�\W����y\I?��x$��O-������>ޤ2��y.�^<�luOO]c��ը�KoDR�A�� bzo$QP�ӫ���[y���2��f"�	
��9�$i� 1YR�l�\0Y�	t|�C�1-7�� 	#��[H�Z�r�/���啓{��	� �k��%�=c�!��Dde���o����&*pI�6	0���"�r9��rt�Q��H�Oezk��P��u�Ax��X&�&rt�c#�d�C�l�jx�7�ί�����\��ft����)@�n���z�y	I�D��\nn�:p��1[E���\�t�8)ǃq5�K�݄�0��넹���L���W���\�o�RA:�ŵ|��:f�rz����=Y�zR�:QQ�&ݥ.�| 	`�iJBEdS���T���o���������z!�k\�P:�{&����S�lt=�oW9`��ՠ��d��W+1�b�V/h��2��)yѮy\��{�0jc��ۈm}���gtxϠ�U�{y$��7�~�u��[����9T��{��1q�� �PR�ݖ�f@�l��҂ �M��� ����J?~,O�=�3}&Br����ا�L����4�\z�t��c�I\s�>%#s'3%��Ս7I7�"̧Y3`�Et��2G��L�kLX��`��m,.s ��لcm�/�y����2����1�%���I� ��5;䚀�Q�5��\�z����k?�9��>��g]�䕿� V<k���g׃��d�g��(�w*���vh$�ew����H%���ʿ�o�L\��;^��z,iYO]�F��M�/�*
?j������>�OӁ����	�5���E;��c��^��H� z�S�O����_�狟1��FR]����3������4�.�����fe� �yAfI�����X^�2U�_>�W��9�9��o������O&_|��\}�Df��
u��z'��:^6ڷ}۷}۷�ȶ@�m��m����ڪ��m��?�������(aB���D�?��xd����rV�;X�T�N���r�I���jE+��g٦l:�q�
	���C)�(�&~}�z8t���\e&��E ,x6�\�nrGܔ�6eL2���ɍ���. W�z���@'�L�B�Ǆf~D�3uf�h0\�C�4�����\��xG����Dvެ�E7��N����Y���J״�W͟I�����|:���L�� 5"0O��nZ�	责ծ�ͤ�L� �����=������[$�q?,����3m��L*�a}�a����sq<H|�3�i ���b%�^����0��0�c�d�X���,�d�PxYVɤ3 �O����da,����}��'-0^���cxؕEi\Ҋ2\^��I���!~�����Va��=(�M}s�%���O��zy�\�qv�B��8n��o|b�'�-��עZ�8��s��ec&��I�y ��)��'b�.0���d�I������1tg�,A���M �~�g"�`n��zw�1v�x`� H5]|w������8�J��8��,�zv%��\�T��Z.//5�=$יzn}�	�	�A�@��f]��� D*��0��S�2��0��sx��4@��a�Կ�_�T_��O���r��d��Y͟K�-��X��y�I0�:\���Z}�N�/�^�\�r<�K�f��YJ���f=�k���q:���}��M.Ya���B��Y%���K��Q%��{v���fy�sV���D����ɵ���B�$)���z*Y���Ny��0�3=��sѾ-e<�$�>��+����fӅM�� �N� =�yp}ϔ�ɺh���>�cܼ�~�+@n�uJ?�(�Iz��jDɭ�X�G "��V��*���Po�z����0_�Lb���U.��+���$2b��8��������rY��� ws�߯t�_�םTt�v!�I�D�`�c�cS���|�+�@���x�=�/(�.Q���@�f�c����:<8��ᅎ���8G]Rq���Nd0���>�x�ԳǺ4rn^Z}����`�n���"�p��k�$A�Z'-F$�z]Te�@�1|�n}��Ʌ�3<���&xG`
bB��՘�� ��D����S� e���4nB�	p�F�e�t�|�����g�Ʌ�ӓ{f8����&� ���/3�+xֿ��s0K)�m���� �����C1�ʋ� z�s�ί9f�^�I��H���׏�Z�� q @D�}�"����(l�U� �W��?����#��� ����+���,��|�i�Y�^�b�`������0�0�4g#�Y�K������ ;,۰i٘%+@䟴�.�!#��v� /�U;���L�JK�C��'i�&��s��ND~��WdC� f�����d����;��Ǹ��U�<.u��\Ⴍ�Q�\�y�I�>�%J{,���U�����z�X�3x����mR������K�)�s>G�*XU�~}�w���?���y���Y�GH�%�L��ŕ������˿���}���j �/\t���$Wϯz���;�v�>'�o��o��[���~��m��m�~ml�}O&rt~"�����o�+'''���x|�$fr��X��T����]�&���#a�6q||�����	IH� 098��e��*��tl�;���y9`C^����*{���#��4�KY@�h�1ɟȌ��ț�F��W�ã�d�$k/e_�č?t�M�k�z8�� EP	��H!;��E�@�Ъ9��.4kK����I�+ͺ!K�UzzN��4�M�����u{m2&�s}yC�In���:!E�	�3կ���MG;��lU���F�f�6����i9`i )�d6���ha�Y2B��B�Zн���϶0/��r] 9P�,�\;&s��h.]�T���v@uo'1&	j��0��v�~86�ļ5|�
"k]����@/���<����,����ɞ�aZ�Eˈbr Ư�D���d���X;Y.�����O�->A��6p4����X�@�-���U�\
���@��0���3�I!��W�_�:��b�p�����$�1!;9!$�|����]^΋��Hb�B���HȠ"s��K�\��\e��[:��{�ҍ���}-���/g������2>��8I%_���=���u��z�������pD$-3�����dB��L��ձMfFv�Z�_&�g"ihr'��eu�X�M,�ٕ�����s5H���A�d�b.2�����Lnb9�}M�x:|��\��V֋��i  ���z29:԰t@�L��"��@|�S|�H�HO�|���W/dQ\�{7�O��Xc=W�����|�a��*����ф\@0&zQ�q-��R�n*�����D.���$x
�%����Qj� ����O�2<� �*�:c�����s�	=��Lnn�r�� �,�ODǺ~�����Pǀ^r��K��1�����x@�⋯n��s=z���Rv����E*�
�O��F?[(B�����R�����}�T���C�͹|��15z�u�g�K�	3�ObW0%��Td�=Zb����QK��ۘ�! �#�C�I�BI!&�H�te��h��t�`���H�fz�����O�����\#<���������P�s}$�k/��t�Y��`��t�T�*��
,��{�������燏��/�����v�6�B��]JQ�[�t.aBP�N��/t\��x�;P�CF�
��[�D jL�+{r��q� #r
�]�[������S0 D�γt�aTWO���v��e�x)'Om�#�>q@�أ���q�`��p
^�{�g����f�Nz�O�>��qRؖ��v}"��9���uc�BM&˕�e�"{��RHiȮ�#x�g��? "
�} T�ao�c���'�%��2D�8'���3�%d����Պ��%==o[[��� Y�9<�dS��!W�U�_��� #UTS��x�?'�9����gA:�2`у�c]�z,t �5 X=`����S��u-���	^n�>3BF��7ߕ���"o��=��ril��1�BS��3��,���/���aw�h���DA�W�l��&�q��e��m��m�~�� ٷ}۷}۷_k�z��ג�rɪ�@��N��W_�pC#o�0y�*��v+��L�c�����5e�:T����V����ƴ�kV	Z�'���FҎIz��LRt|�$b��o��T�	V�W�������N��k��=�BR���H�~�m��/~��%4%�$V)S���w�Y@��K� @ A9�,�Z���3�_ ��D��P����#��L��	 �=7����A�I�ڤ1:N�	�DȜt<��9W�8sTl<Y�p��I���^���4�+f�,�^g��m��yJ0�Ȱ����u/�%6���l˕#�<�w�1�p#��K2'����JIK���������~���R=t7U�:U����K�N1"����́K�=�2a\��8��͎��}��Ru!�ѕ�r&�H����ױ����ɫ�l��S�"H��aN���O�Jqi�$Th����� ��C�KNl�1�y���{1�$�q-��y86N$��$�|���'�\�.�My}��Kc����e�w8�7�a��|}�Ͽǳ6� q4�I�o������@��l��>�%9��"�#JSD�ħn 6훹{��Oz�ݡ�do�hw];�L��x� Z�f��JrTS��W��k%��JS-Sc��8�<5���8:_�����u�]��D����#�:@r:�T���:4�_��@�;DRJD� ����J�cJ���i��ԠL?b�5iJr���(�Nc�#�H�٬ dF2�K�L�iW�ͽ���	k9�f<|{��Q<�YTr��=�����:�c��DMW6:o ������S����2ZI������\]#�\�����Jz�J�S��d�=��V�.s��kxf�"�G�29�X
��ĵ�Z:�i����T2�����j�"�����������Ƽ�F���U�t�</%��%�����U*z
r}�&��[8F��Urt��q$f�c�$�'�M��B���k���Kc���꺗�}K*N�s"Ǔ���v[k<1�	� �X��8y$�����Vo���>����2>�����C�㧉L����Mi��$����d �L�c�4�Dʳ�mɱv"� ����q�$w�.Ժ� `ٔ��uFz��ޓ���c#e`���7�!$�B2���� bn"n�y��1h����:Đ��Z*�����Q�-�ͳ�<k��%�K�K�3�|�(�u��V��L�ֆF�U˴ݹ��� 2;h�5vi�=$�#�Q�5�G���]% �"��a�S����Hi�o��";�Ƥ;�(�|���p��j̘�%��pL��b4��E]���޸�=�d�ݔ����J-�oȃy?�?�6����@3{�,��lrY!�N�&�D�f����H��;��[�B'c�K��̸��}�x�*EX��<�04� ؁$&ye�����J2Oml�yů��Nn,qǀ����|D���� {�X�"�>+� ��n�q��gA/�g�Ralrgx�G�.�X�v�xf��c�M`�`����>�9����,i�Bh���S�IK��X'8��Z��a����h\��`0�t^�Oyڃ�@���@��P��gߗ�����>�H&GS�G�b&k f���?�����_~J�>P�z_;`��]�����g�w����睦	��C;�C;�C�#m ��������M�J�V=��0�l�����xBS��c�FV�����n�Vٖ+���
l��:T�/d:>⦈��e� �T���S&&pn���%(����B4�v�NV��j���G�Vb��~:l���O\ubU�4B�a������W_��w�ޱ2�Kq������-��{~w+q��Ma�2x-�	p����3I����&��-�1��_`�o�kq�}ay �̎n���D̑�}&������I�mc�Hb,��U�w\�]]�L��
L�<��\AC��ƿ��vП�
���0V)m,�Ak�ּi��Ҵ��3�������
�"�nͤABfO�j� ������~�r�������%^|Bͪ�����ܕ״�'|�� �m�����j�nf������O �>����>����5�����K]x������-��Wj�_�~��>�٥�	�yM��3W|�7@��"U�3���׮��d�w ���AU������/�=Lz�p�����=���$�S�j��v\69�9u`���X�K"�\��F(�u��V�W��x 9dW4��==N��T��d*�j��ױ��#����QY\��3��]Ǫ�S=�UL�&MY�j�H����XW�XV�S��g29�X�р�x}-��Wz����a�[�;�MA��Ƽe=���D�P�S�2�/�v����TƧ��!�(���$�wrs��)��q��	N�7z�Ap9Dr��d)�:�뫕�y5��k�����D���Lҳg4z��j{#���(��ɵ�0��z�~@�t!��0�D2���>��BNK�=�jm0�t~u�����R�z���Yf@�,�+�D2�����)���8>�K:)�]^����k� � ��j\G��B>k�HjV�Y�k]2��!1O@� KVv�#2=:�Q��G[�d٬����$3�N��aB���H_!�O���΀��Br��L�� P�'d BR}�� y��:F��*�B��N%�O���:��S�k=�-��!�#�͈�P6��潹�<�s����g=]��ĝ����:�:���<c���tk����L�<K�B{��ǯ�L`Ϋ6~z�t>x��Kztm�5�#x}������Tí*���&lk���>��+�p�V�#��k@���`�Ɇ�S�E
�D���}�& 4�x&⸌<c��8lAfc����C���00��tn_x��q�9��(���ýܳC���KW��k�1"�Ԡ���5�ڕg}t�zb����˔�X{z�ƀ��Hÿ�3Li�ҥ�j������'&�x�l�i�޴�c�a؍�=`��"�oe �����ɹc|x~�e��ދ;\�� V\�c��-�¤E�s��p�=�O�spǭ���d�S�Um@��Y������*n�v�~���+��1��>���I��u�7����1�Lz���gq���Gg�ѷ�#��(���@�sHM.6��¿1~�����V6��T���_|$>{.}]��Ⱦ�||��� K>�P�4���������O� �C;�C;�C�����@n&�p2r_�|��Knʐ�����e<���ݍ���O���Q'[�\�yD��p0f%�b�dr���&}�O�)�Q�t�p�L0(.�ۛ��tJ�s&oe�)��i��M���	4_Q���2��#P3�?0����^�HL��]�#�xM���~��ǆa:�������; ��ib����f3Y-V;
��IxC�wq׈ߕN��<4B�D��	&$�aeR�d�ĭ�G�$��ˁ�W3
M?>t�)$ќ�f�3H�8����q3B������! �z��>�윒HXvyn8�
��ܒJ�w��q�`d�f�ި�-7[�� $�ۓ�H�����1�7Λ�*�d+ik����=Y����B�˩x������%��l��vM;�|Bo?��op�1��GMn~!!�ݶǦ4������7m���iy)-�h���'��?g�������W�l�����3�߫T��-~\�����ׅM�kb�O]Bu�r;m���/�'��f���PN�Iy/ T�z@� �:�uv�
n&׺���H`º*7�E����Hz�3`z�d���q�� ��2FPa��+�c�! ��X^e��X�[�ǀ�^0�'�QX��i<:�my$�� ��|�M(������j�m :�G��)W�t�$�?�9ԗ�\k�Yp.&d��H���S"�䲼���|C�cYDr�?h܍Oͼ�&�RPQ��|t-��V�o/e��(��|8`����f#o_�d�:��m�ɊZR�p�ئ�g�^9�����!��I�$��>��X��L�+��x#˫k�f:_�ܚ|-��̡\_o��\\;�Y��G�H<�3���ߌ�б&<��rz}��� 0�T2�c@:k<��+������q5�E���	9�l0��hI��oIWw$c��K=�wz�*2v�N�����%�7N���_O���3�8�6`:؁!�A<��� o��3�:�"������55�� �\����bW`솰��ysTdz�dk������>fQJ1,������P��0vS�0�sвI<h�u�w��Z��ۨ�ދ��;�� �6��h�{�Ή,U�C�^�/�x�K��tM�
z��d�5\�+�I�*>?�z��������?��d���tS*�7�g0��6Y�`�DI���[�aQA���؂?��_���ߙ�YI@��}LE�2ߐ�J�̯i��>��fE��f!��"c��Tl�-��� ��Z����|T���M�d�ٳ�%�'�jwx֏�� ?rn�d�ti���� >{^2j�NX��˙5�L$�MT�=�k�%�2��G������c���Ȳ���<d��0�$������d�>�P�xm�cJ�`0��X�,E#��H�n��_����>+ʞ�/Z�j��+r �a�{����Jڹ�y�.�
u�����7�����9>;7�N�tϜ��5�g�>x�1���Z�?y*<}&��P����y�J޾�*£�����z�èn����_����?�ȡڡڡ�Ѷ rh�vh�vh��N  ��6���e��N>��o�����nZN����g/������՛��[�/���;d23q��MܣG���'��1�A7{��geXG7�HD�����{R;��Ӊ2�mW��f�ך����'�` �֘�t����eu���ڬ(}�*�a�/���|��|��5sQ��H6˼M�`��j@s���uQ��]U[m�8u���QJLYKHq��VM%(+4�1�Ye�?V���ͬ���.yL�Wa��NX�W0)G�A���(�6��	f����ȱȞpI   %���7�Dã�MT�B^�v@�����	$�A��ZU��`������U�S�
ˬ2#Ĩ��- 	Q�5L�!Yׄ5A2c��o����"i�=4�(lA�l�|r�=@0/��*���VSJ���Oȯכ֟c�ű�����	P���H]�y�$�gx�*PBxƊO��󀂈��Fz|�;C�}�7�7R7 �X!H���]��ICg<{���z�Irms���d��L^~����=��30�;�A�c�����ޗu�k���409��Y5v�*�;�����2HN9��l)�ёt��yuerv������V���d�I	���D6�T�$$.ل΢	�a풖����\���6����}f�B	Y�h��y��?�k�Q2�:��k����`�hlz+�NE ����XV�D./.�͍�b����x"Y/
��{5�6�S�#ō��[I����):!X%+	V"�Y(�^oȚ ��?EE������>:��u���NY�~}�s}!e�!�$[��SR�/Q�ʶ���&��|�D��� 3%\fu:���wW+yw���;]�����5������Ӈo�2veq���N_����딐�wr2��~��P	ij#�c��y���Wr}��d�f�QB�a���٫;)����|�ggz��2�^%i7��͌�f����c�a�Gc^JU٥��v7�����AI��̩}U;�8�¯����
u�'}��$�	N	e �e��=`��ķ+J=�a������Mz�8%�l�o0< ꓫ�d��y//��c �M�g�����}����M m!^�e=sĳ���*���!N��p���`��#�������& 
��0������d��3�HgO�9SͲ��4	2 � ���C�=�A�   M�3<"ct�n�8
�d���05�_p�}��X�t@����]C���V�N�)2�s�E 5�c����+�+	;��D4�' 4Jw	H�������߼Hj�ф�t2dA��04��%��`�7��4@l��cHfҭ��9'�u@F�&�˨����3{v��N�5פU)���}�Z�#�W�؁{��}St�mJ{���A��L�%4}+���y�PliB��#;�0+=�6̔`�a9�s�BA�+:`�	�\��N��{>�s�*~��v��ac:H��1� ��w��]��?��$:����1�c�d<��12=��&$t���>d��P��@������跟��M���L�PFeY�L�����폲 �C;�C;�C��5�i�LG�9B.���~=�߯^����o�n>����/��/�|)�W�L"	H�Ұ���Ul��0x�?}��'���ȋ/���Z~��_ɒ�*#m���b�u�h:��i߄ܒ&w5�$��{3nB��Ix@��K6F�<

@�E_���dv{�M����2v�����S�U���X.�9�uS�i8�J����3�j~��{1�\Y�	���%䗛�L�c�M#�ɱA���K��<!�ă�?�]ߴ�ѶH��z��c�br��k�䱙m��+I�*��p��a�n`5fd������3���`�9�9��Ip���I|P�������磺�M@{Rl,���R�ӕ"�z�m�֯����e�1s����0$�m�Z𕗕��6��MRz;�Ł�� A[�X���v�d�y���M�Y��i���|�%��G�e�$U0��hBR��>���K�{y(���	"��D������ M
jg��h��<X���,�d��-!ظ$�Bj�S11�d�P�k`Ȯ/��@MQnY�Z7q+�c׷�윗���:�=�i/M�s�gX%qG���k|�}��&�咖% E���V�����$����9ޭ�;:g�d��e~���yÄ�n���qmI��ti^�O'2V-��S2vAHz$�
�ˊu,uٖ���*�U���u%�y%:3!�T�B�/jl��S�����"w2�%��L��s���Y-�h_�i�a�=����T��"����)���+Ж"��;��x�}��p�c!��䌂D�]���3������?���)~y�i\�+<]I�XI�)LC��Y��tBK�Y�(��!_h,\f��U.��B6L'z�'�炥�L�]3J^�������\�&I�v�!�ɓ�<:��-5ơyek�E��D��#��.��E�}�$��c}���|ND�O"9>��3S��Ӄx����\>�RD�,6	�`��sr�8���E"w�cj��*�С�=���:�h�1Yl���,X;:��BV�;��_��;`  �,�z�����!N��ڿY����t��]@�_�b��:g��������(
��ܟg>�yp�K�a��<�<�&�>^�y� �c��>.�Nn��0jx&H��y�	�iV��L�Hf�V����Ho2V!�Z"�d�e�c���P���t2z(��q��A�8ԉ�蚭_1���� 8�
�\&׍8�������=���ky����_�\�cױK0�r�_!�5��>�U̹�u64땮������숅X�oC��R�B/�]�PV��ۂ>y�}?��/��C�J��q|�/ݺʅD�����=�����?>�k�f� ��}c�X��ܚ�����Cc99Ae  4�.
:��AqcA���dzd�*��b�Կmܳa� *���q<C^p�^��a��彼:�?�P��w-r�����s���THw�04�/����T-��o��T�>�p �
���|j`
��Ɓ5xV^ܯ$;�2N���w���1��g]W��(��{����i���[���
���^?��д��&��5���������S��΃�B��/m���t��9� �}��.w���$ �x$�q~��$ʪ�'���yh�vh�vh�� �ڡڡڿ����+�u����V("�D���7���x2�۫;�C�8�]���_����̑�����?���kyt��ӷ�^���N�nD��m�i%|u'6b�<y�]��m�t#��^Qm%�����>=��b97�T%"�бt��]Y/��嫯䋯����B��%Y���u�`:�������I���7 _�c"���tz��[��pT��ļ�/�,s�]�b�d$����gC2�ƨ^���L��D�P��fC:�����ZK
w�Lh����6?6�Ec@�'E�DC@�݆:�h^:�i�V��>�+��|�z��EY���Mk���n�4������Q;i,���"���ʆR[f�Ɋ���PE��3i+��X���Iz��!].)��*�M��x՞�~ղ7���;Ϝ0 a�\@ۗ�����c��O<�G�B�բ������O���,����޴|�$}�����&0�����;�V�������gn����Zln��8Fi8����c��>Ccg�쓠&e�f��3[l^���jռ�P�|���z��>&t��ER�n�ծi��k0Q!�$:G�!��V����0��F�H�s�%Sd�2q\ )d�4]V�QO�����b���k�)�Φ�;�B����1L7���}%�s^V��*��Od<=�x:$8�� �K��E������* �!*��[�ѳJ.�.EØ�q��H�=���`�D%��0�J��I�����R�	A$0����Qx�|��+�?��{cJ�%��IHA�jy{'?����8��0�^w�}��R�xι �EMJ)�ׯ3��"�3=�v鑞�x�tK�K�1`y���+ �"{�\�!�ϱF霈0/*z|��C�N,�_�^��M.���啞k_hR?�]3����<�@��Ô";�vI��(Lh�"�;��	���zU�pБ�S��C��>��/d|��G����5��Tք�*�� 8�!7�q�;�c}c���b@��Íd:?�&��.��=���%����l~1+۴���餡���l����V�g-�����Z���2�V����Z���=�|l��h���>�e�r���7>ߗ�ۗ��~I����I�Z�9�q	w/����tY���S���Z�亸.V#jW��rw��[�8�X�%2�"Ɠ�+>W|��߶�·�)Zi30%�ϓ��G�2���I��g#�6�Q�gR<h<$u	���@���kS�"�����
����̔وP½u,���U�q�~����P�8�'��v&��/T��Ӵ�FL��{�iLf��yĘ>v,x�`CVK���kN��ā�;Cy<�Dt@Cv�I�z��� �g����({-��č?�&y)�O� 6<��R�&�P��jI
`���`���c'BB��c�\��c�9��i,`�w �1c9�gS�:��)���Y+�`��ج[	9��G6Q�ז�݊�x]n\�F���nv�§�'���;��,h�	x���y�F��g�±����z%��RwWF� ���ꚝ|�;Oy�C;�C;�?�v�vh�vh��m��Td��d��)�*��Ⱦ��T��S9>��d:���N#\������H� 1puu%�߾a����_�Kh^9��U B�f�o����i{�&6����
Rof�]�/D�$|�?���d����D�<�uF�n��]�]�zw)_��Z~���/�K)���|�YՍ`������{�t#V��G�)A���t�cY^\�|��^��C&�q�QMy�y��.�ؼ#����!�
nM��$�"&z�-S�of6��ch����2��L{� �����&#"˂�R9ֈ_���Tov�J���2��^���q��29ªc����Y䖐, K���yo��*��0��M��PA��'���>��MU:6�X\�)������������=�/�V��@/������C�,}$:��C����$�=8F�Ʊ���U�y�����h�����N��'?|�5��7��;������2��i�ڱ$v�4�Z0"�x��b`E��g�-E� �����3F�m,�c�?��A-�{��~�<t PH�q�ߕ�7=�'�2�Rv=�	��J�����x�����yH��cG33�-h���=�^��4	���.��d累�L��j�˛w�|����[?^�z�a�1u,�~"��Z�,�ZFÍ�+�ȵި�	���>b|AX�v&r}aXɣgC&G��|]��_fs���]�4v�2!�꽥wI����@�=�4���J$��d<��鹎ݭ���_�V/1��i�t܌�XS�9dP�#8a�N��<g�<-����?���8��G�B�X���\4��]v�dz�`6�?ɃD�C�"�Y'�U�FewQv��e��,��e-⭐r��=y��I�@���jdi8=�J�'�w�浞;��T�ҷ/�L'	���'˻����<|2��a_F��?\o��MC`U�\�5����0��aM��&���67���o�L��\�@�����09����L=Fb~ ���*�uy1��4��X�5��RG��?����!����H�~\���T��^��ǟ��	��Ǡ�^Ю�9���p�I��X n-�=�>[#H���:��87���S.�#�����z#����%ו�q���q ��q��Eإ.%��ZLF��Z�ۯ��/��B�?}"�=�率���#��g�6�{�CFXD���[�_C�5���B�U8��&4󭀒}oJ�_��yl��G.���a��_`}�<�P��S�O�栟Z��@J8�I��9��~�ܭ{�d�y���>s�HǺQz�G �?���`E2�m}����IKy9M�G�Y\�7&�F��!;=[G����o���[��ϦQP�@ou��W�_Q%6I���}��Cj�ˊ���d'��r����)e^C���X��V�(�3���5�ME@'-y	:�3��� ^U�~1�$����{��5���Q�%��8	��<����b���咯�,��b&��麰��O��X��{������4��]cE♮��&Ǫ�2ܳ�z%��׺������`v���~�`�8�����e��9�C;�C;�?�v @������M @_�Ĝ?z$��>��?�X���n865i�kI����0@5��d�����Rno����!���L>��s���-WousTs�?�I @����0>�cR��UL�j>/���f��7zH���rHo�WL<�f�A��xw�N~�_��w����L:]K��
�.�]�I/5υ�6������c�z~������[�$o)ÐI��|d2t�E.�H0��U<�#4�O�@�@��<��ľ���p�����6�$�θ�&��N��kP�5�M/�prG�jz�0+g���Y8���Lg�������L>;�U"фq�4J�8p~��:b�
J�4!o�Dv$4rV�k�M�� B�	�+pz�qh^ @6�xζ��t�X��N��׮"z�M�&��=�c{��i/㥢��x>��H�'M�lZᤲ<#�30���4�<�k�b�)z�B�,�p��޻��V�?���?O���=��r'c���s�l_�ƒ�I�����(�c~y֊�_�'����Dj��ʙG��/F��!�u��1+��2�2�[�d<���<�=K;����/��,���J|1zPCr�9aG:�4�x�yAӢ1_!2�?����|[3��BkۇAm&�ǠV{���2�x'�ٕ�׵<}�ى���N�sN�$�Y���|�6��~t)��}�.�{<��b&W�����ײ�+�a,O�h����������	��-|9���T��X/������zL(�|�Dd�]6�T �!��G��l�1 ����A�������17�!+��\_f��*wwNB��ؐ��G�N#9=Me<t�w�E	�IB�v�G����_ˈI���������=�T�aS��k��2�DǛ�&�u<�R9�s��c1o�=
S�c$��3���e�a���KD/훼'(�oJ�1�ܺ�$��߰rIЈ�'�)C
߸��M׳Ъ�x�鏃��u��c�[�1A�`'�ԍ�y�8��Q��2��!�Ĩ��@�u�ښ��H�{��Z1O��e�s���̼9�o�7*��Cn��'�^�ǎ�-���7�?�k����{z��-�
�.���ð��=�g2�����A�*�f�_|<O����I����}����u!���͋����ӧd�<~�X��S�D���q��B ��x��T�V�_�u� a�@O����,�cE]���@�`���Ӄw�?ٱ0ܒ�� ;4D����0q:���eP�@m��&d��Q�<6`s�����+iOQ����"� 0�cޘ|���	Y�����l��:{�|��}�a�Ccǲc��{���u]���j����웘�տ��D^k�8����rǱ!&����ʳWQ\����{y3��5_:Nƭ�&���=� ��8���xb^$`��3�H�������N׊�zE00h�]|Kx_���D��V�:���,�@Y�-�\h�;�o���;�����gr��!��~O��r���{�_�O�D��5�]���|ų��W_�y_r�OG���m5���������h� 9�C;�C;��N��o��?�H��/�R�����p<���U�6d@��C���
?V~���X�NO�ŋoQ��w������dv{��������vI`T��I�`?�Q�%RjK�09���oT��]]]�x8�k/�]�}��%�.��akq'�..d���Ō�5NQ��MM^LR=h�H7�Q���0��.|'(��}q��A�7o^S�z�${������/2@$��=~hI\$n��P9���
|���bF$C��	��='L�jxV�"��K.��D8H���t�����>	��@�ڌC��@;��86���w����nrQi�Ĭ���;5�a��L>W�+�ȃDF�c�F�b�b3�v�'�%�J�R &���0��|�O��f"�zC��V:	��S�z�(�ޫ_]ܴ��0��w>�u�������J����{�*J���ױp�>Y��>���>������P?7<+ƃA� �>��!�J���I��$��g�M��F��/��H<�wcx��X�.��fc&� )[��S}�Y�N@N��Pes��oz_�m���+*�ɞ��~�zm�����=�ʸ>� � �K�A�ot$��YE�У�wYC��B��cJ!F���^�(�98I( Kq�lL���#)�#��הtzx�c3� 
B$�`Z���Vn�~-o~�k���R�Oj9�I��8�Ө��{"�~W�J�q$O?�Q�l�ӿ��ݭ����t��Ͽ��~�s���H�Oi�]):���d���fSi�J��N��4����$}&����+=xA��&�%rr�H:�o���5�Gdo`.����#��0I�ƻG��H� &kpU��wKy�����M�Q��h"r~���%��1˶�?pȶM�֐u��q��[����|�۲B�){rqm@�`���DǢTm��}��Þ\���ז�N:K�+~d��4���,����Fno��+=���X�4�-�!����<."zS�d�"�A��U�d��O�g���1Cc���^�< I�Ȗ2j �(���~��#"T�c�E��AV����������w�Rz^���%Ϡ@�|�v��ǡ}�<����΃a?F�u�ܱ���	L�ﴟ��i�Z�+�=XU��ˀY�U�5q�@���d�rw��I��� ��?����N�L'���39?{(ӣc��]9�1C���Ud���$���
�Dv S�笶?�'{�>�=�tf�Z �·�}��xň��r���!Iv��^x��
K�ǲ ���ހwH}ekqH�>�D-�"����V�1W;������!�s�i�Z����?�0��Y�?���Ub똍q߯�^)6�����@;��9 { ��\�_/J���K ��N�+�!䭼�-�~�@�>Y@x��-��FcƼ�":�u�1|>���l�F��\ϣl(޼�Zc�\޾}�ϴ&g��A&mi !�OMGߣ�"M���"@6���[Y�/�2�_|�\�����;��xO jtc�R��#J�B^���Ɉ��H�I�H���{���
��(@8>>"S���H��F�iW���grh�vh�vh� �ڡڡڿ����8yp�P��#������Xe�Y笪��&Qf�܃z�]�A���)�� -�.����?>���7.)T�	��������G�:�%2�A��%iJԬ^����.�0��*��cT�Qʩ¦��>��W�fH^x�i$>p^�w���������ӏ~$��?�H޾�`�'�Q!��3��!�b��gc�� �`|���Y@V�0��Y�|zI��sH��Ќ�k/�a�AHҵJi��eUڊD0l�6t;jj���jLh���� 	B�Pm��A��Ee'd�@�$?t�!3�eH\��Id�WQ{ǎ\B�4�Cg��W�%}r�'�<؁$:�;O�$�J��Z#�F�R��>y@���o4$�i���Nǽx�����q��$~�R��3�ص�ش2�Z<��ke���;���'�%d"�@�s̓6���7��}��_/�m:��r����T��o��y�l�t�I/�@�9�'IMJδķK�d�$&��萁���d+��䛥L�c�#�{��t*�})$rL'�ْ�A9"�Kǹ܊���C�����ɚ�:��8�M֨q(^��'��Me����I�+q�җ���W���>�L��Z���s����d�=?Kd }��J��~m��F���^��I�n	8��7s������+�� D]�ͧ���_\�FD�?yx��8�{�]J^ne>���� @��&���J�#�/zn�,אJ���^�|��P&#H�T�F���λ,L�*�S�O�ε^���2�E��&�	�%� ^�jy�.��k0���/H���r��<B�~&k��P1t'<��*��=�赻��y�P�K��!��Q$#�؋�l�Fǔޛuq=��XN'��*W�ኵ��>�k;2]i|������l�'yx6�s�Yi9���L�^V��p�c�{*�AO�M&���jWH7eH��N��>-AŤ. $i{�y��;4���@�]��M-i��13�2g��X��<�tNh��1��Y�1Hh�[�)��^l�@�>��ux?����X9˱�]�
�gx�����e���՘i:$)7�z��<�-+��t�om��C�c��I�$��+��ݞ�Q|���Ľ�ο�_�}�<������ϟ˳�O�vv!�W׬���E�����b�H�^�9��hBr+�[�m�m�Q�� ������&�~F����v����rz%%D�����5���evw�c<�$�=��+5v���̔��r@�3��&��d@1�G'�����2����&t������ܱN;�yowL_�����'����LVe��u����!��1	���`��\���q�� �)�x������H��\󵯿�J���;NOO�(>��r���!���a^�g1<g��K�Q�-;��Ƽ\Ү�Dc�����
D4*__��?����,�q�b ]{��|�Ͼ'���F>��c�yJ�?=:/w�B�Wx�����=>��F��<89���c���S��%�����O�������t� 9�C;�C;�?h�����ؕ���u�r*Ϟ<���L��j	$��*d�L��(C��'Aj`�m�h2���YM���'��?r{�u2	�Y,�d�*ĠMl�����=At� ��4a�s ���*�X�fUm�
���qG��S}/�])�4|���d��� 
ILl��dE��@޾}-���������g?��,tS
9 CH"�Dz�ݐ-��*#���M01 |,��	��%��A3M��p-H&��C$��൰�5 �����<E[B�K0��DJ�//=���t�]�ӘT�67��g���C�I>/d`��+F5�r[�1Q ����`M���+�N��4ڑ�i�м�]R�'�k��+)-��!�H��;:d�f��~d)u��4�#�O"x�(_��A���,9�����@�y`��q	�oʻ��{q����h��%���z]���i���*���@N�)��l���k7����>����Ŝ���21sN��)�^8��Iиs�	���}��z91Kr6�_	���1i8��c�!::�Ʈ�I;R�<��F�ڡ���[�G�Q^m�>����7d����X��x`�*�oJ�X&�1@����J		�2M�����{��)�H��c)�Ah�lk!� Cl~wA�k�'�;	rRO�D^�%2рP.�����<'[����#�gzl����0���t��2_��/~��&���\�}�g�E��a"O�4]�b����=,�4�_��,U$=��#_�5=F:5|8D���H�=k��TXQD�SP{�k=�ʼ3���,�[��ͯ�u^$7S��U&�W�̖"k�a"!Seo�IE���`���#��Z�z#n�z�2i���9�J�[��s��z�Oq�VRo+��J�\��u&��L����<8׃f��wR��S6��Lt����gs����rc'#���3��P|���D�%�u�Q���%|(!��- �7�5#�����_��
�5�����I�;
�g���a&����� R����x	@H�m��z�P��eC��j���8�|o]�:�?�(�_�n�b�g�D�}����7^�>��Mσj��x�/��zI��g�Q.σ� +�4Ě
)7���$��86���t�!��p'�eRX��Ӕ�#�ޜh�Ȇ +�CL�S)6���o�7��J�?y(g'ǌYXW���ήu�"^��J�������`�� �#Q@�M�z̆�l�P?'��0��Ń]�>xE<ߐ����h�*"���b��K�RFww���`�>��	09טY�5YU��P�W_���J>��:�F�	�"+*�I��"[G�LУ���mY�x�ӛ��5��!�/|F/�L�� ��5�lj�����V{����gQ[�Q��>�W�O����Qfƕ�f퉭��K �:n�7`��g�B�g��}�>@�d��u�GkJ�-W+I5��yT�k=�V�n�x/=I?���A:�C���S�X���Q�1��P���̞����N�{��:Q �ۅ��/�9	��z�5�����_��������çO#lL4W��Ձ[`���u�ۙ��2����4��$cQ<;c����?��i�������D� 9�C;�C;�?x۬+1��ɽn�O��ȆF��)�lu�t���-�������4�Db8�(k
T�1!��A/��t"���w��������F�./hP��8@ ��z�p�w~����Y��]�D7aMP��@�<�%[�BxK�X������ن�xc�h~c3�Սg<�4��x��IM|u�n�F�����Ϧa�n@��sy���?���O~��ҾA�(6�1HDC��ؘsmT��f��m�"7��_����PZZ��	�=����¹T���$&���D���7ۮ���"��iE����jR@7���)#V:0IH��.��GL��R_���$�FfEkGb�)�D�uI�JB$�����I�j��LB�}�-}H��L�z���4�?E(�&�
�5���<�d8���#a�o�3d��U�wM�!Y�+�q]��;(��cN'��hL�ѧ�#M�0!��;0"t/4�����>��3�< �y�Y"��<�ě�⻯��>h�I哉��lv	�����D`h,�X�g����#���}	0�?�[v�>�5�ŵ���<�2&X�����	K���v�聩k�/��I9S��@)u�� :2&��E��c�����2G�DW���&�#g�k�K��:�T��m`�%2����3kp�Fr_�!m�B�dr$���rɔ\��+2	�:'�W��G9;I��
Y-JY�*Y�U2[�&"'��߄�$`��<H��ӕ_���b)�7��T��B�;���� $�3�E]������MӓE�����{H�=� IGW�a���z^g��X�N�-��F�{��5B"j��rt֗px.�j?�o%���,��H�:mon+��C&2��^E��,�8ZJ�d�7�����Y���üNH� ���]��ٓ�l�N�7���B;���@�b��g?�a_�1�����S��^�:�FcL&���4N�rw��h�H��{���\�t��d����Y8\S
V[z"I��P>%��7���ױUP���F�ʆl�0�>G�BbL.�9H����:��bc.J<���W 	�L�{��n��.y��!�����a���@LBB8�^bL-T�{O#2>]L�s�5vE�~D>>��ڃ�����)���}��C�h�`��2�%�B"s��/M�ݢ�oϪ�玵q �au����H��|H�u������G2����8��qxrBp��_|&����N����W��l�h<��	*�Ky��B>�^��X���q�3�P��S
�K�qkLQc�V�_V�bj�,:��i���#c-T���W���=Ä�PVs"��:C1��@�>�����,��pK���瓤�1�� tk���*��qO ;�i�%:�c��'�Ny�}��}�,���{K�8�c�4��/����&7�󯟈��}� ��Hy��fy^[�l�	� ^[�`�6l�ze�`[���)��TRV�����I>���gA}��]�Qb�ǎ��@��58.�O�L�QrՃ}�ϡ}�����	s^x�Y5S��� O��r��/�����y��#�L����\,�9 �nwt`��\N�ؾ������	����2ٯC;�C;�C��k ��������͉�R7�C��v����R�i�M�����/��O��k5�<�	b�� &ţG�t�����H7�]y��1��^B�� 1��,���r����LF�K�2����N�;bE4��A�[7~�d�]Uw�/5���z+A���qBM��;���j[K�JIRh[CJ)�pS��1�^����_W����E�M!�AJ����������ꗿ�l�r���Q���x��m�$26�X?c`&� ��RC� 	3O�k �1�W&۫���3a&d _�D>��#js�A���;�Bc%d�,�ȕ��%���:6�H�u� }
@�����%�n�M�@X��b�����/���H2E�Ȩ(d���;$��z���]6LF$�R�9o(-O,���R��Du�
��xH�l��ј9���%܊-�7�#:.A���Y`�M|7q�VƲ��,>Ø%�^D��<h�^�(�����}��Y�W#�dn I���OAe�|�68�1�#���A_���:�z���Ҫ���p`/`<%�P��� �h��1�{��7��J�1O���H�Ҡ��#Y��XիU	gk��1ɺ\����;a�$��0��D�
�CjݮI^��g��oRi0�v���^"����/VK&�pN)�H�v�'�3�%�x 	z�P֥bl�%n6z�P6Ն���4kG��=��z�Nފ���� �g��$4v���p��T]�lo%[�h���U��vOΟ�%�g2^䲜�w�"ÉȃG���cΔ���7O�����K=����d"q�X�3*�K�W�c/����&�s.=��"O�e<Z�ҿ�1g���f.oR����?�ht.���F���z�}��B��د�{Y��y����0��[�ZD2��d��s�ZX3��.t6�r�!�>�X/�H�\��եCN���c>/���q4U�#��pXݛd֫�"w�&K��~t��^���T�G R���{Wzo6#}O(s���A.W��<z.2y�Hf��z���٥��;y���dQZgS��@�b`-��h_f�Ab����B�vWʺ'�~I�DGu��u�fRE9�E��|� �'J ����c�H�_�0�8S���י��Xv�4��Z��w|�x���-���]�X4(����^�ҡ�wʑ������4c����Q\'����$����g��v�?��� �ŒU�"nAV1ֹ�d+�/�����K{��#�k*}H��f�zE0�RL8״�c!Q�Y��R=��H��aױ*2:p�-,�O?c�������~����r�g��hB�,�0�nf��w��+���j�ヾ����L�y�<��HW����Ky��N&�s���2�{��g�n<�5�����,�TlP��;�	յ-���:��WCa�s� U(x���5�%Q�<,v~l����l���I5��wj�(��y(%ȑr�c.��X6K?%��u��ױ>����N"�c������4&�	���Cɤ����&w��q�"�LU5ԑ�lm��޷��{I>m�U�+��̾��Z���e�1k�T�jʹ&T�`�N�����;�k	���z��^c_��D�D���f����[>EA�co�s<��L���`{w�"�$��$Ԓ�c��7�m/�NaHr>}�V�3 ��/�4Xb�3���wr{5�5�'2_��Q�����Y��$��:2��d�?����17u.�\�5unuY������g�r�i�_)%��[<�k�_,ڽH,C9�C;�C;�?�v @������VE�[c����n�
�6Xe8�o^}%?��O�?���no%��%gb��l�p2���nĎN����/��@bR�|�%6M��W�
�r����K9�1��Z,���t�6�͞�8=�����gu&����M'\,bV���R�R�+�n��ʀv6>C��&.�k^��Ve���%���r~/?������G�F7�H\ ��V�Ws3^�摕�`Bk\2��:z}Wz]f�>�d:3��mЯ����2��!o>5���0�u}��B��=W$���MP�2٦���^�l��q��Hd���'aZR��`��T���;��q�jW� �ޓX���&(������x�ً%dP=I�P�g� � 2-��4 ��"��+1Nk��&NZ�U�2�M'����W-���`/eI����;q6@�r�
_��}?Pq���h�L� $4�*K� �W�;���j�e�lϲ���ƛ�{ d_3���{)3_-����{?������ٞ�/��Y��|���)\r���o������&�bI�ڠ���������e� �yy:Ĉ�@ʭ�*��E�9p��Q[Nf�F8��c2\`E	q]3�m|!���Jm���!|�s��ve�xB4�q2�B�L'�L�i�s�^�g:�&r2}��/Eؓ�G3rx3`,A~�?�k<�l��C�p%������>�񙬗Y�%��z�P�������k�EF�HE�;�)�*��c��a�M�v���$鑌���]��dm� S�4FV`� �[�� ��P��	��3���&guy�V�OV]Y��#D���6��~��cG!Y�Ꮰŉ�/ �2*���,�萻[f��"��/����cg����H�OF��/d�A*K�����*��}1���&ȵ�nn(�����h��?���Ӈ���cJQ�Cp�*J����՛r;�d6�i��X�爄��X󍙞7�*��5fЎ�҄	�nղ@0��*�����t>A1����� � �P����g��z]m�.S
Iڦo�'K�w��4���Y. �XC �8~���a�>�p��A�u�m�_��|l�1�|��6�x/��ܭ��ic2�2�	�86�tN���X-��!��5�I����ZPHAK�����ys��\�?�@��s̈́y�{-3Y��u�Fz~H#!B#^��p4I�����o�bUo��嵎�[�R���?:���\v�u+��3I ��q�T�2�B�� �]�PB�n ����YlW;/�&;I'�̷��Z�|@��賛��.���1X���ɶ�V&%V؁D�B'=X���`��9rU	��"B��"	��_�S��y��Y�09�w�e4��O��h�u�I+���1�:���t�x ���7Y �؈Z.F�M��l��.<����@�:���{Wٺ-\0?�m���Y�K`�w������-PW��B�%
b���iE�4���N@�Q�.N�̛h���Ll��&s�cNmu�ո9U0y�@��
�8����mQq�@���n� ^� j��3�iS���ј6��ȸ���~.�߽���r��a+���4dX��Xɡڡڡ��� rh�vh�vh�6[�������!�Ҷ����:���~�{�ٿ�D^~�{馑,�Rn�j���q �m&7�nȎO���|��ߗ	b��eD��nC��b���!qu}� ��n�f<���c�ԧ�V�cS�Ѩ�C� ��}�l��	&vRn�=�rK01g�R#�(�s�?;i�2躤.�d2a"~vw+��� ���Wy��+�#�|B� �H<A��wi7q��&M�:�Pv�{ؘ������e4HeSl	<@:J, )�����1���gѾj3 ��p,�FLR�
�ke$�qF`rTNc�L&�c']���ZX��@�����vf��{���Ed�Yպ2t� 7�'TA	�,7�v�I�V ��dP���7a90��BU%:������;��vt(�7�+Eel	H~7I� �S�	�2����&u``0����~���⨈x�P�I�$��`�� ��$���II����pᓁ���Z�l��֏d��U����IG��f�IdX�y�L�M������|���`�O8X���^&,j�1���!�A��!��A��$�'IO��>�S@�r�� �a�ߝ�.��������}����B��0��D��ʐ�c�/�;Jb�>xPf�J�K��a�.X"U�����!��-�I����jI���C?G&�#��W��ul�K7�4f��2��Z����h����%|C 1u.��| ���f2�n$|!A�KRo�@�"B��#��k���dvk�[��[�H|SҴ:��ɂ����=4����f�b
��#�S��z���F^��d�D�9�3���[}�@�
GyG�e+o�.�Ҟ9�.��g����Ɓ� �`
�d_E��r�W�����Hߧ��?C�E���D�$��L䷿���_�02�=SWWK�gK�����Iw<04%���s)�\ѵ�e��x��L��M��D����{��*7: �g���r�G�$�U�hA< ,U�Y�o0"�Dn �8u�T�xO'��LZ�H Myd%�N�M�F-���>عЯk�X��Y;����ܟW>6y �r2�dQ�uX�g,J��|�0[ 4�c4Lr�8{Cv	��0���}`Hz���9��!s���$=Z��J�X ��#@m1�k�F�3H�}��C>g��G29~'�����8��I�1`ܛ��󊸹���՝�.$H����z���Η�q_��L�����s�1 ظ����q������0���N��1
Hla� �(�M��-&�<��غ��^�<c�>@����I4�W�0:~����(J��Ohx0d��U$}��VL�AVi�gz�ffNI̎1A�/�X*$�5�ƚ��%�{RX`�?%B��y��9�1Y;�9���i���:���=�(�Y�v����3i����1c��p�^i�P��'�}�`�fd�v��/�v�H�}*�?�	��PL ^��<w���6c/an��K�h� ܣ F��2�-�b����h^}��̮nm=�ҥn���Ї�� m��׫,�W�^ɯ�SY,:.���� @�C�]-����W����@>|��������d��(J�Sk_�t��&N�vh�vh��G� ȡڡڡ�� Q`��� � �"�]7�tS$׺9z������B��P:+׺y+f$���6���������d#Py9I����	��Yt\����z%�RMK&䰙J�>O�����������'y�}zIjzǡ� i�U��ru�q�YT&�S�9�I$+��W@�?�2`�	 ��|����ﬔ�t�%�~�&lr�kV	7�d74L,���~�� ���^�d��zɤ��tzLl}�������f*��*�}���`_��v�VzN�����3z�
�.����vL �<AJn�}�����%��Н�k��<K����"�� ���?;F���a�b����6�K� IW2��d~�ǎX
N���̀m���1�g����cEdW�\���~�x`��i��0��X�ڤ���hA$����x�q��H8ژ�Z�H�\�=ȁ>�c<C?c�������m�3-��*gZzO�^����ݪV{q�VW�$��|y?�}�N�2ܟ�7AF?���w�$��^�/����]��V���]��n�$L���C�*��Ƀ�Q=�c�:6_pl�9�i���6�N���dՒ��`��ȼ*���% d�0���u�o���1��0tF�z�~���fR�kǴBQ�ƞޙ�	%�$,es��R�6����Ha_��X�w`������<X���#	Ƨ������,%�^���ْl�u%��sD�w�{���h�$�2��%�QzR��}�^d2=Ⱥ�L�HM�d,j���1�8g�^k���Rz/�ʼ�'���}��֒b� p�)S��Ur�_w��Y�$z��{�-ev-��%���҂@��f�K0,7M}$���+��,�������M�K��F�zM�&��|6�ʗ_L��9t�4$P���P(�I$��_rg�K�fǬ����AT�=�C:��2��3��P�^f��8�"�9쪒/��e"�S!���x�R)�	�}0����4n�5f��-��Bƶ�OM������=� ?,��L��ϯ����1���6�:� �cKঠ�0�#&�����d젎��%�z�?Hh�I�Qт�tH���w|���Blg����@�L�qp��S8��	-���V#{Ǝz�o���C�����c�l��d�|�j\r���6V�1�-�[���;��>� Ĵ��� ��7�O\H��r��:����B>L�rv�@>��2��(ͅ�X.�� {�����g�k�\�s��`�������Q�/�9���~@�9�H^�D�N�_�<j���`��L)}F�3��0�X�!9���©���c�t��o�݉�[�5 �&���5�.��X�``b�8cp��j?z��L��y������7|��r����#!��}�2_��!�6F :\���فX/�W �~����� q��s��Q�`��գ��K��~Tkq���O�nK�c
�O����x,�թ'���:�L��7��g�E:����9l�'���2�>Z��p�AO���L��OP`Uhk��1vְ��h��=��ua`&�����>W0�Rzd�|�ZcĚ� b"�E�ؒ(2��c]���W_}%��,��[}�Vϻ��}�A1�:�nMi�gϞ��~.���ϴ���s��2_��؎�؎���c;�c;�c��73�h��o�(���L�t�p�;�,�k�HBU�3���<���1o��n�ܤ�� 8��}��I�ۄv�ײ^md9�H��[�]�&�aV��vNc�7hxQ`.�$c�6�B���qo@ �qH�v{}�tO�:���9Eί ե�4��g��?��K��O*o^���dz?�
���&65���`iG�����+C�߉Lo�H���`ʍ
�<��*�QN�hT���'� ��9�  �1$#��ߨ��=��!��5�Y�Mm"UT��2��B�$V�;�Q�I.!	���Ч�	j�JM\l%fډ�P��i�^��A (���i���t�a܍�0�I�24&i��A���`C����'��t@���Hx�$:�}�1#�0xG����Y�;3
Gý��������m�:� ]c��K�őU��}lr1i�Nq����s�c�0ٚ�;���L(��܁�4� �OPz���!C�����ⓐ�SHD�%Pqo�AT*WNBL<Hf�o�D�!�{;cuAR�ޖ�z�g&he�����x�Vb�K�E���>1�gZ��U�d����x���Z�Ӿ����K�st�5	,Ļ 1�%v�U��ܡ�'�`1P�y��~۽	Z�i��D�h
�f`��K�[�d��;�*&췛H���?` ���f6���Ņ=_�����D�'����EB @#�J����ድ��C�
�NO�ﲙ�}���2H��ch+�^Ho�P��?�_���.+V|oPU|��՛J�=V_���'#��Gt�l��m#}�Jn�� �6`g3�rr�c�S��h��n]L͘�eUv�$��*٬!	��r��]o5��>�x�}BC��0�ֱ��U��� �õ����+ٮ#9k�x I"�ǲ�7/>��m#�'���1#f��z��BV�ȣ'�����|%�mJ�2x`%񀱊Rh��^�o#�|�!U)A
Ȏ�����x��`�5&HϪ�r���T<+��'(w��{Pҏsr�' ��60).[���xΎ�q(���S�В�����it�cI��L4(��wd�<�� ��\G���	 �##�>o��Ds��b`�+=�� �Z����:`,�R7�f�P\�7�WS��&��u���D&�r�03ƙ��,��֛7o�_(�=�/?�T^<{&k�ww3Y��L�u(ٮ��
�U.�M!�ш� ��\�ϵ�o��˓wV:��
� ��d��X8P�a�B����J� ��X@Q������)=������(�9��u@#�����{b3\7�K����\�(ہ�y��fb�tJ����k�Cs{�������Иf���S��uQ����*r�<س��2~�����[�
�=0�M�$����W����1�r�𢹹��V��d0��O�b֞X'�A�iG�����Jf�d{a�9��������Ru3(� ������xI�߱.��9]LgVd��D�^�1�/���7X���\��Ҋ0���9`l�}{��蟐OE<����b])�y�t������Ypܞ���xO�<�7Ww�gݤ/�vl�vl���ю ȱ۱۱�N��>�͙%Su�V���B����t��R�[g
����K��ƺ�.�@�P&̜!̼���K|:��(a��i ��VV���"Y.Vrvz�s@�f�e��Ƕ���+���
���U�b;����(��>�B{���a�&u��Ø�����Ѣ���_����_�����O�G	]�L𦠶�U�
M N��瀂n+��sOJ>�=�記�@ptY�Ko�B(�P�F&�Q��b����KD�<�i��pHQ�.��.�n89>o�ǲ�]�,2�1�\e1��I�d �D�� "��#C�hM�=�`�_i[�9		�oJ0Ď��n�����v�����X��@�%����>s���_�)'��6"���?|���*���f��6�?�K�̆�7G^��<м�=��gL��g����G c��s�87�a�׻@��]�a��^J�_��͢����!����;IK�����Z�^�z�;��z='7��w$G���Ƞe��k����F��{؄��=#�3_�5��,���{�V���>����9�����[��d�4i��L"�1<��C7�>�1�R7IXS��>5�)��fbRo:v�P�]�V�`�]�f��#�8�3��E���{0G.m��΄kC$�aO�z'��V��y]��d$� �4]=��3��d:n�2�w I�^��SN�#��4�F޾�\�׹^Dc�n���I� �_2�9��
���D 5��.Dr�x��+�T��:��}F��j��5�#ԉ���$N���2J�P�.e$�6���0,��xm��d҇)���G=�����l`x�j\D�����H>,6,z�9L�7:�&Z��N��/dz����K�h,�㉤a��&c��H}f�I$��䡼��ȋ�w2�U�&����R�2yF@K�\}~HƁ�����| H� 6 ��[���]���Rd/�y�%�k7.Y����B�c��>��5D�����	-�,�MI��ō6�� e�(��/�U�cH��V�>��a\g[_=Ӌ���KEU���1�'�W�r�" �x)!%5W�ʙ������w�3�.ؔ:O��
�.�9c�B�I5�G]z����������|������\_i�RJ�-0? �C�
��V�HP��杖	�_��٬#�^3��P�!0��9lF����K+���K�QS��@
�0�6�c�B�?5�o� ����D��@	Zq���W+�l�4��Y����gۘ4�:�"�
�@  E���c�	���l!��Ӑ1 G	 2Z��Cf��Q�ɥC��F<�TZū�*�٥x�+c�$(�L�I�}&(n���g� �[#vL�3�sn���>&4�ԕ���u�-%K��@&㱌}99����%H_!}��"��t4p�c�Y�1�+_� 6Gv}��K[�\^^��}���G�}$o^�$��%�d��q{�,���'���zq�D`�P��f�J�ɝn[c���;�	%eL k*ۮY����l�728ȱ۱۱���# rl�vl�vl�3Z�HPcG�bh<�f�|(?��;n�߾y��iy���u���90��<|������uP�&$y��Dr��39u�Qٿ+snʝx��3�NGr~2�����dyиj҈� e��v��#c��lU��V�a�օ�@Z�A2�H��h�dq�^������~+��o!��G�]�%����喇Ma� ��;qw�����	H���m�	�TV��Mf��_0�$�F��,�4�����R�Y�gt�V�Jn�k�@�! �9(~G�1�Ӡ䒕W�O3Y/�>�!��9��.4���Έ���;�8��|u<���&"#��:�E���i��
\�R^5H�ڱ���" ����a���x3=0��ϱ�9�{�C�q�R�&��Ü\L8�MlB� r���lL"%j�7��0��/ �*qƣ�HLZ&�L	�!���=h�z���L�[Um��B�\A��4��aW?�PZ���.�H�T'M�%��,�@��`�<�����5����g��dry��-^��1]z$����X�MY��_�����7��N�X߫� �SQ���H0Zr�K�5^P��3V�8n�3�uA`Z�=+z�N�����S�4�1���!�J3�^�A�υI2>"$�{��$@���$����1����uН�чd.,��RC��	��/�BVRgK	�렟7�{�J�� �E�NI������ͽ���V�%s#�ߔ�wJ� ,��6Hq�%Ծ��1 ��d���"�Xc!|�����u�D������lNw�����VR�E�1 ư����L���CN���Տ���L6ԠJ�0���g �Q�Ū�}���R����B�ǩx���ä�p?��<z�''g]��B��J���q:��Dc~\��#N�z3yUY�<F�@u�F�s����@�K���b�tޡ.���] ��a�q�;*�3��ִ|!�4��d~����I���ge�[DW ��Gsl&(��0W����C�X+��`Hdv40��]l��w�C��S| ns\��z�^"��|θ��8y��Nz�q�*{��� �eܠB�ƺC/#/�w�R#�C�A-����H�"��x8��6`��/�IҴ��2`%f<�����C�]L93ψcL���
�_����w�O��.������!PX? ��&�$B{���|����WCOk��B�)�1\���A8��P��:�m�w� <1nՁ[T,�0&a�D�rA�1��>f�y����՜�����WH��ݕn��F\FB� ��H���_���z,�{fB���dw%cw�B����?Gl�$��~�����	�#rl�V�30�/�LB��+ϵ�yE#, ��[�󍢠Ajw��L�M�dVy�0�hDƩ��ޤ���W!��=�5�~U��ϛ-��{x��sNOOe��:tRa=:8��ƣ!=4NO������vC'e����k�s.�R.�L��^vn�a-����֟�^��^�2���������~��>�ڪpE!�{�R��AI}�(��7�!��DV�)�G;��U�(����O�[���|��c��c;�c;�c��iG �؎�؎��~��{HH���M�
�U���pO7����w��=�<��/���&�H@������97e�a���o~K7;�ᆯ�m���b�N�%gU�ڐQWݟe[��MF`4��p�{QU��:9���xLb38�u�G4"G��7>GC��*�JVf"�[�=�wFL�a���uh2	ڎ^��l&?��?���������L�o4�aw��ʛ1��;0i�2L6A��� 7��E/�$�wAy�X�k�#�L�]�L�{�ojzgTA%]e�H|Ŕ8pՊ�H�wF��>�]~Nq(���"�U�I@�V;���C��2ULP+�~�m,�Zޮ����P���7<e"�-�1�sb2��$!��F�،�%�PFSr-0�n$����2�W�O���7gO]r��x{��zLԡ��㌂��>\&;4��]$(CK��v?-YXҷ#w�K�d/i�*~=(y80�<k�3)<�3#�o]�'�{<��%f��z��a�W^"^�
�Pv˟�OzFȡ�9������)�Kx=��)�xLJE]J����K���L�~���³��Y�:��^�E��$2�I���bҶ*�{���F<�V6���2�����n���K�5���8�o�+}��Em���eA����;�����Kڟ��ԝ��r��W�J9M2�����SJ�t�������etƓʀ�<s�똌ۮײ]�e:���.�G���C�a4�&��Y ��'� ��K�K��oV�X�l����|��Q?�AjjL��x�p��rG+J��Ѱ�=i��9��QO.g��{7��Oq��(`�̧� �7��m��� $��U�Tu��k+�S�7f�\��V�ZZb�?�<$�Ʒ�#��S�@^q+�eAI �g�J?}(����M��o�7F��'��������`����CD�}�_S�<[�zV�}�l/@�$�1�l}G���<�X��X����>����W3�������y���@��-}"�c.�y�2xx��j7o���a]�����C���/m,Db��g0�8UH)�����;]~/q��v>:��@��Ƙ+��k:<���x��u^�k|Bq�3��ml���0���b>��q'ύ�g1��ސ�1T��w2U��QTP���,y@��um @�^Q`f�4�����L���z�lg�����q$�'��w�#����'���g����&2_h����<#����e���\�u.-	��P��I`Ay)�\�@{��0�G@��,4E/9ߑ��,(�~��{�Ҥ�0�#���A�Rǃv�dk TE�K� v���ԄĤǙ�T�M�^��~k�  ����8�@0YH�����I;���3L���,Ȏ=�X;`=�Ԙ�k�RdR��  d� �I�rq"ƚ�1��џ�:��u���w���E{�c�p��$w>C(�b'W�9T��."\�؂%��1Z��;&
��\z���L<��n/��Fc��Ņ�e;&�	@��uFA�4��1e��)�%.m�9��!��?��������Ԁ^h�UA����&��F�;�-��3��'O�ȷ��=����:��2���xF%��21a�B��|����O�#}߷�%-�f3]˱۱۱��# rl�vl�vl��V��#[r�
}����k���cb�酬0�ο�r���\_ת4u�Cql��8pՖKnĆñ<~��	�������������+da $H]Ҟ��r'3����e���J$�_�|.��Ԥ���r*�Q�2�*�&+�M%L�� ,@��rrYHr THS `�^���$�1	O H����_ɯ>���Տ��<���u�
=��z��5���o%���S�0��h���f(�����}��M"JI���S'P�HF*
�����+Y�ll>��������F42-턛�Z:zNÁ��t�[3	��{M��l�i8oV�d�xYʛ4&/T��Ҳ�ױuU�`��N��7��0�HR�|�%�b�'��}^��;�_Z�	��\����ɘ|���� Q�_`i 4���t�;&���(�gӣ�,ci ��{d�ĔH�Y}`	'�>��SN��'��|h�.��'!A�c��aY���`
0�A�rҚ�>bri{��{n������ATa�Bb�>�h}��{<x����x�V^z@�WD�y�*/yqX����sq������c��=�Ʉ�כ�Ϟq��Vk,4rrr"�]F�����L���������S*���\�>�I_.�j�4qa�$��#���ᲑNX0�-�od �
wn���@?J�Ğ�sOX�]�J�~GS�`BV��V��s�7sʉ��d�Ϩz5��ٽ�澑L�e��Q�7J���A%'�DF'�\�٬s�/��;��ճ�dM�M.����@���+	v]�7z��l֋���)c�h�ʥ�� ]k����
��II��I���eO:��,�NT���Q<ni�j�ș�MPݮ����@RSe��S#�2}�@޾���"��ܘ�t,����Qdx�'P�ðn��A�r��"���!HО�  �����q*�IM��"ϴ/�:g���_�'����b�85Ծ��E�J��S���"=~�"C�"�"�<�XUu��b���7�rr����'��tNz2Č��G}�|p.�͝4:otя�\F�|b�7Qi�Xd�P��\;F�C�ܘ��D58<�(��� F��j��v�G���+/���j����f\�}!��1�m����w���(B����p����sV?\u�%pW�Ǽ%q���Ƹg�y s��t`�ް|/9ȱ���\�@��A@�r�q���?v���=���;�(p̗U�7[ǹ-�����0������?D��d�Y2^��5��`GKjJ i�1!e?-��5B�$�/:ߣp����H��� |��'r?���s^Dά�$����ݫ��۷��|ｧ�A�����N\�W��t�i�'N�/�Z�
�_����7�O�oab=w>iٯ R��XT{?ie$�h4�]Χ���ڤ�P�q����y��H��#���Fc8�d2�>�#h�sF�@O��z����a>��DȢ��)Ȓ�Y�XÄy��G�Iө��;���d��D	����("�0����5n	�!�lk�."��U��-�s��5c�dZ-V��dx|<3���a ̖��#]C?8��>֜��ɱBJ� �}��菣�@�K�<u�31VG��Nty��Њ
�\�vؿ�ǡs�D�� ���jd6������ɏ�c��_���+]W�@��}Ě	����h����r�y�;0o�&��� o�/6�>c���a�\�����O��B�8�џ�����P癇���k�
y�����rl�vl�vl8��۱۱�o�y��`n���b1�rC1�Tß���p2d5Yb�W�rZZR��b,��n�߾~#���W��_�&i*�Mf������<�)n%#��Ͼ������܌�f�$�2��	v��ߙBj�0r/�e�*�|� �ۘn�Q���~����\�_��'���������,^��]0
$+/Sd�E��ljG�sE�c5DQ�*Hߊ�M��B�=$� ��j��.�֔�X�
��I���ȹ.ץ�w��\ۦ4P	_l�|����� �C�E��J]"�=HD1�P�Đ73�Y;�)4�,L�uQ[�̟����Yii�#�߀������W���w�Z!�!��*���F�ޟ�|#'?&�8&�E�Ȯ�����s�t0p����4gzn썜 �#��i�
��b|�M�������wi�I�Oz��@����s�20����!&w���;��B# s`��>w��84/n�`yx��z�w��;_�Z�F{��<�,Q�l��V���B9����.�������pv~ ԅߛ�{`ȼ_콈>��+��}`;�J�&[&�# ��L��L$��F���i�%�<)h����{!��8DNp�BJ�t��LN��i2��?���t,�ߘ12b�&�rr���ړ��\���l)�r���h��g��12��I����L�T��	�R�x]�
��]	��+
K*5%�����rr���tz�Ɓ�U�i���8��	�\���IC�=�q,V��5$�Ɠ�ex2a%���ƛ����B�ۘ��y������>�(1����s�So,ncN�b��d6�Y��?��)HoUC����0Ϗ��"�4z���!���@_�)�\�3��'r�%��e7ZJ��>Ĳ��$�������"2�< ��ۼ'o�fz/�c�x֩�2�x$zc���Nv:�*�'�?�^w��"�~Ǭ�e� �kxZRB@�(��K㘌�8����u7҉F�k��x`1�g ���cH�$-[���\� A�m�uX;�X` �l�����p�z�!��{�t�zss��@�!��T6�ot���]�;��;�C�ڱ'��6V���}<����2fTC&�p�h4�붛c��������ı0]ls�4���y�Q�B
��p]��b�����Ԙ�И��y=!����'��̹θ�A -� iƣ���[2h�7��"��̇�Y�Q�*�y��䊣��d:�ʳg�Q�:X��_�X�f�ǓHk(��37���=�^���^56�W ��:��_�$���˷�:��`.�a�B1���D�Q�~������}3�F�
���:hߟ�ֻ��X��Z٪���B�O����,a~���"�+�݄��r���r�WyE�/9`>���s����꟬�ퟹ���Db?@������1���3�U�[S�L&��(Ĩ���<ac�y�?�g��#qE}'����t�{9���(��?�����Z^�|E�X�SX��#H��2Ɔ�[I�qt}}��%���Nn�����_˓���1�9\��k��X4�ޓG���#^X#�=�&���~M�<?��ڡ��[K�۱۱��o; �vl�vl��[k�ȳ�l�;�C�^��`<��+99ˠ��'*�.�&�ɖ@W@3fՍS]r�4�
�����_�B���E~��_��n��	D��3�_T���x=�5��W������Col�,�ǽ���n�����M�Df���W4�L����q���q��c�G������O�?��<��K��/)�w�ܼ������9�� )XH0򚅾��Gc�Q��ύ&d8��G2	l�i�*�b/M�=�G��=,L��l;I�Lf����1f���܎wUAy1\#X%`ol�K~ ��6Y$K w i01� �#d��+E!'A������7f��̛c��j���*�2�X�	��Hf����3�G(#S�5 �cot��i����f�H�Y��~y�&����X%�nKЅƼLj[Ră&ЬO��߄v���'�QIl����О	���G��,ٹjh|O $��zǇ#�lh����O*z��T��C�Έ[i�,+��PZ��'�}^��,�\��'6}	@�����1W��"!m�ɽN��D�)}d`έ�>�_�9����9UM�"'�K
�/R&x���g�d���8�j�ppʼA<ص���t�f�&b����҉v�������W!�}��i?A.�|yK��d+@��KvF��R����~��x��ٕU�]h��^Ų\*d���� �$���%���[�k�k�;i�+�0�4�/��| �!ez߳���X�i.�!�S��H�L0*��m$�H6�d�Z0�;9���0�(����U72A<�f2��?_�r��Zd�3Y�*enq=C�>��Enn�<�r%=���`�4$��|�T��lPu�f�lZi�7�p(�t�g����{2Z�>��b��_-�����[_-ry�v!����?�{��`H>�I�1�s6��嗔� 1�Fr҇��� ���y%S=��"K�̉^7�[���w��z�=��R߽�f���I,��Dv�[�u.���=6��0dH5BB,��Ԭ�Q���h��RWHN�4w���3t�d �-�S�/�����Bc|/x*�q΍� �9H�e������A h;��C* ��j�e��}/�Wu�r���.���9W0�X!%�Yh���b���`�HD��8&>�Wv�Hc�5�v��Ɔ�=�u�X%�i��dz��[�T�ߴt��3�"&�i�l�0A��i����g�*|��y�gS0�Nu�%Ӹ��f���N�`+� �� ����3c�^ *
�c��"�<!d�����d��Џ�O�*g,L釂���cyu&&P pLD���_8��_;�d����T�,��	�3|`�Bțѐ����5��Y�C��1br��F�|��C�D��m��a#�5��2i�0�侁%��Sc���ŃŮc�`|yhc��b,�ɱh���J ����/.1�t�g��;E�����UIƕƷL�7��R\����U�mPce0��
�����an����u0�!���31�8 �jK�d2�՛����[��O~"��������_Q�,�WDV,���1[rI�D����^����� N������C��P����F�1��(������� i�C�@ju3�5�_�������s1]ɱ۱۱�~�# rl�vl�vl�3	k�:��|��'&!��O&gm�$pB�����`���T�Q��,d���������_ʯ?����&���A��;!�ʼx�ٜA"��/��z���p$��O��׍Z-˕��"��p��m(�*�'�9�f	�.*�uS�ןN\]��ۻk�~%��?�_�������ם��]��'�Hnj�`��8�$i�!PQ�����k��&N�
�!c��L�Ԕ����E"}����m��.3&�gҥ���PA�!��!�]b��k��\HR'����S�ϥ�X&���Zr�br�bb+`u}Ih*�9�%���hk�>�l�E�`B�2��J�wA�Wl	z-�3�
U\W��T5�6�L'V��*ղ�=�w�s$�M��a���RP���Z+n�$��23V\˞Y�z]8� ��n�
��,��4�-1㥤B�v##�u�?xx���:���0hZ��38<�"q��O�J����A�
6���L>+�3⫪��uP����M���	C���O�(�������g�xf���A:������8��'��g��2i0<34��-��={���x��]�� (�և ���j�J���(�qnO����x%�n+Ѝ ǅ10*�w�Pp��%o0�& [$�a� ��F��7�P��� I/�"���0�r����+N�'��7�ٺ��R��0��x!��to���"!�/1�Z6�R���_����@>��Ƽ���3=���t#�D�[�f搖�� Ѭבͭ�9p��a�1(b��*�R���FN��*YϦ���=b>WoV��e%�16hޭǥl�9���)Q���J� R��Idz��٬"��!�-L:��T�'"O��}�耎�Tnn*�~�1�@�+����k��R�g����tNu�������u}"�EE�*��� �H�z8��o����)������7���9���{{*�陜t�������"S%���z�� �쏈r_iXY��� @��W H�#���.e{��{[�=��X��l�^B6���L��N"�����>@Pk뿨�Ǹ�i�����No�b�����P�{Mv����W�6Fp�r~=>�zp���y`sHR��e2��wƪ�nx,���fY��g`��69.\k��v[����:�Րd.�sc���e�g������@� $�����Pe�d[�x�ѱt�8��7�-��H��JV�w>���u3&�	�R<�k�!��`�m^,�g���J�?�K�"׎�����.O5���\dH�8�S���,l���
l���$@����l�1�he��,1�+�c� ,���$��r�é��+K�����@\��\���P�ӳ� ���f���3)�7`��\{8��H�����9�v}/tc�i� �����IQ����`EGv��c�������݁.<�3���	�Ȉ�s���ԍƇB㵮3�"�H�`�%�}E+`V���	  � r�m�N��a�f���.��� ���S���3y���7�M(`��@�����F|. ���[��յ�����ٕ����������ji��E���띎�Z���s�����r�\۱۱��}; �vl�vl��[k���t��䆈��#V��7+�~�J./�J�6�e2Q�b�x�4ȃ��FC5�b���r��O��Hf�w��2k$�n�6�����B����n�=�2���d<�Q��!-��χ'��4�֍�F?8�V��$G��Xu�6�m9����/壏>��?���hj��=J,y��<��X-x����� `����2qk���:�ޱI���̣ʓ	"l��$H,�8Ҷ�H�;/$J� wFߐOA���b��UQ"�EU�2@U���U!�`���.!Q&�M��s$hV��ߡ1���T9�B��_���Q!�v$�� �iJV�5�ɼ�4{V}T��{aн.d��"�̋�	�XbIź��w{� �����3�{K��p>�,����ƽ�%i�vx0#�<P��[�uCy
�G���ɬ�jM����ȨJ�X���Da�/ :U��|���U@n�oDL�wG�͊��k�׹����B��x�����V���8�R]�>Yi^%k�b����c7����֟��X����"-�dIM;��s��(΅��;��r�kL��ҕ�|��)+Y7��>HD�"���� ͆>qh�M�����v��R���X�\�uVxN�mEM �,�fzV�H�g��y��զ���œ'��ɟH�?��Y&��R��'��.K鏯X9���ޭ���e��,a��J�Œ-#��U�����D�p���ă�H��I���F����j���Q��]�s!�I�>�ٲ��}f������kY�$ԫ������T��U��j�C�=:U��<CRz~�3�:26��}����Z^<�ɴ��ͳ��~=ƣ"O�̎�v�XEr�6��/s��&c�F�룺������䥾��@w+�{�n��'��ۑE�'�d��2���\�}��'� ���nԓ��ys?��v��{'zb���б,݇y2|�J�K��U>���f)�xX�t��'�]�8bB���I���nN��"������ �V��RRrɒ؍�Lƪ)�6�Li�t���a��1�hG-��e� �]��K+��<�ǔ�q�����}67X�rʍ�q��
�}ZД��j�8� :9ˤ�+`O���N:��h �W��(k �a�g��;�*�� )��e,�y}�%��}1菥>X�Y��z۲�`0.I���i�i��^o@���L�	q��k���fj���JF�ƚ~=�� b�C��w��*:n�(tIp��xR�&G*�(]��`�<���=c���QN4�.��W���{\���"�z�v�ɬ5vNH�� ��X�� R\�p�	�a���#2��m2P#v��ι��;i������4#��="cv�揄�K��rzc9V���# r�KQ�v�zGA�$�����]go_����-�4V�����婜����Ʉ�B�\��{�Y��Y���1�efb>�����װ?�����_|�c<3&hڥ�]��T�����8&�b�fÚ���ޘѻ5�����|��oɷ��m�|uikx��v�L��2fO�N����,�z_��T�mv{#?����������'?��O���?�c;�c;�c��oG �؎�؎��~gZ�IА�0�Mٛ�����grvzA���6����*�0Z.���&�c��Z������W�_��ݝ�xoK&��4u�C��4#N0�#}"!]q��$+��,t�F��"�f	�^�LzE q����������֍�x|�ʴ�%q�6�B�?�Z>��3��6��-{�����
Y�3ɲ+�O&'Tj�I\n,C��#��Izl g��E� ��{8�0&�dr�=Eń+�ɡ�]��B�%I]r؀ J9?�$�Zp�22��k��H�Dw�$�b�W0C��x/�"�E!���]E ��&;�%�}� $���F����v�l3]Wi6x92:p���$���B(f��/@�KW}�j�*CaΉd@��b%e�3e"&m�6�dz�B��
&a��q��eU�`�y������ �TP6��"&W(s�5�����Z�|i>�}{s��*QwLd�L�z�@�ԿK�����n����H|�<Aw�k_��礮���^���L�Ȓ����7��@�O,zt@�ă#� �/�7b�c�ӒqA{N�ijϧt��*�0���˾�퐽rx�s�3���gOc��Vv�VI�g[��KvL�W5t�����g�ۚ��z|T�g��x���� �L���>��2�鬔ׯf���I����:Kһ>�SČhA~�4��l�|P�t|ϥX�:fr��h��e�e)(}���.���� �iG����D�;���d[K�q����DS���ٍ�n��Wh��+Y߿��8�sؤ2E�v���S��'�/a,ޓnZQj�0b��0dG�x>�ʛ׹�V�}E���%��<|�~�M��S��^��ן��^	嵺����xd�\�n=���������F���&�H��������ZZyF��a�#y��8�d��=ϖRo��� 6��/�w���JKf��la�k�
$l%�8 �36L���S�����B��^��5,ea?#y|��#�=
->���#s�I�U���b��<H�۶,4�B$ܙ��u]̭�q��	�z+�X�Jo�L�j���fn���*�8��?�9���?/�H9�[D�q-�Y��|�g�����M%%�}�<Ӄ?�0�c����bC��s�d�{c2�����>	Sl0���.�x���F���b �7�]������2Ҹs2���x"�<�;�|�al��D;�=�Ŀx���p�����o�Ս����`����PIF��U=S�s�K+J{	����K�9��q1�
JƓqW�k����[�V�����'vs=b�k�Eb'�e�3&� �ghx��='Y&�gvl;�5!=� =�9+@?(��s"K�c�r�q1���9y�������4��X�^=�T��@
ˁ!xIv~앲�[���~
_�_ӹ�����p����?���u���zF�.��+0��Y�&��" {s}-Ͽ~!W�o�w����V'�5�o�������唷���1ؽv��?x6_|�̦X/?��ѿ:�>X�Xg���L���mm~X�3nB�Uϭ�޾yE����Oe���c;�c;�c��jG �؎�؎��~k�(�%��m��뎥�lTp/VKn���d���,�K`��yq��Œ��F���ܔ-V�f��Oh��\�@����n�*`UH���n�HI�1�9����-c�9����d2��P��2,]����sy���_�<���lֶYD�?�M�r>��UF�J��0�eWd��v$�"2`Nmu1�E�zz��Gb�ܚ�$Bd�������I�8�*Qh�74�\��n�0?\T��S&VYUXA��n�}�<�;Z�ЃjC�!�@C�ZH{x�m�����|3 �f�Uˇ�}=
2D"ʮ44/'Ҹ�wWn��K���g���u�eG�����Bcf ��$�N'���'��_m6��i�yvy����S��wd��lW�U�d0�>�*�÷`�z��T>�ov��YEt�echث�[�ɑ��jT�Wҁ�zb�1�n_�ЄI�U!�l�}�FהpҾ���I{46���Cv����䉓`���^B�{So�w6�IO�А��c�s`��H�qƮ���By}v{MD��uw;��E�3�iLϾ�[I1�m0���>��|�[Pџ�?����0S���*�Y���4�,�~!q�^˒VD[��d��'�6�b;��I�L�+=߁>��*�ʱʪ2�s��x���QcQ]�iT3��<b���_�I	(�AW�1q&/^��tXC 
����$�5�r��#�si�$�AI��nniA> �EWn�ry�|!�UE�I4�"�~��̦��O;���V�Κ���&kZ�z_'ˠg����i .Ez�NǑ��5N�����B|�t�����eDfIO�a���| ٫���V�aA�m�8�e.o�dr{k�)�����(�qR��Y*'�=����#އ�B�( ���蓧����4[��%�t*��1��^�B��B
}��D�0u䞊f󰁁��#}�8�k9?J�4�x�q|�\毧r���`�ǋ�E4k��{	0�9ZO`�w��!���D��B�i�=�矜]Hs�j��ؤ����<�}2���(�ga�0FT�^��������{�T������0~غ�h�d�9Vbƪ��c��g�A�'r`�1��L��Q\����E��_qIo����B���C�cp,��^"�`O�����%��:}>��$�E�}&B6��If��a��܍M�
`RX��Z�Zc�|�f!�	���=��L��NW���Vƪ�1,���H�T ɦ]��Z�����e��{�⥎ۑ��s�#q^��9F�Ñ�(QJ� ����ϸ�s��n4{0�r�{�-X�غ�l����_�`BL������ݭ�U�bo@v@�򟝖�ù`Eh�X�Evd���癉<'�K��7���/�P���d��i�߄���<�ť��fD��!0k��ںj�K��Z�X�+D	+������Zff�g���|�3�[V+o�q�{w���=�w`�c<� 	 �1������k���ժ�^5@떍��l�s����Yݐ��<��s3�<; ׆`0_���� ?�r��0c���@��$�pK�/���r{s%��=�w�7���K�?k��|$�����vl�vl��{Ў ȱ۱۱��4�^v�)� �\���BZ��d�J�HJ����W�]cëfVed, �CI$� {`U{'L�a�8��p?'h-��2��]=�k��=�l"��D�>���@٘���۝d��F�3݀v&���G"Y��S��srv���O�*$����1X��^w������M;cUj��V���TR#�U���Dи�(��*�YWPW�d 6��9�~��~?@��d`�CsTl�M"D��AB �$�_�����U�y~��	�ܲD�Yj>G4;~e���&OAϐƊ����k=ƶ {�k$�(�R�5�P�fP�OT����a�{q�D��_�H~���ϗ���3����X�����_o�Z�z�bBb���x#q$|�|��Ɯ�"�X.v%e��+K�a���wy���)����@�>7�����> ����#gz~H6!� ���x$O�>��O�gEo__�]�������X	�r�	f>!�A���ơ��փ>��$�dh�(�ښ�.���i��x�����{�|����f��Y*�@�g�1I'��\�=�r�_:p��~$�(u��b|2v.`�,	0��ڳ�t�z���0��ձ�Xf�w��K�=�����ca�_�G"�酭G+���)��B�wM&@���$G:C=F�$l`����D\R��v�_z}}�1bO7#�5���:�i6c�����cU@1�I^�=��?_P��	����C'��2<&��V����۹|���	��"�C�8J��˵�Ηz��v)��TNOz��[�w�`)�ya��e���{����TDãG��x�Q*�=�5 �H�˕�h����1�y��LN#9;��|�sF̒���I��R95��
��\fS!�/`|���$�a%�I;HΚ?�RT�t���sz,��h�ޠKV.q�����T�W2�������X�ڇ����Jb�T"����w|�2d�"c�B�qv�P��W�a'Bg���S;�E�9�EP=4�r��`��d��A�,0V
���7|����;�8�M�s��mxࡱD����:�ݴQH[��|�����ڬ���K�جw�$������c�!V A���:۸���FԼ:V�|Ř��`���&���a� e�(�8�����P�����@;~���=z�������]���crQC�����;η�!qWl)t�`k����V����T�ɗ���bDaD��^9QaRO�s{^.�����Oot���Q������C�j<����_!�F�����U��N{ѣG�����ΣC�O�//.0�����X?�s�-�疺1���q�ޛ�Y��0��}���v���Kc^�)��u�\,��?]il�����)�!�����y���5k��p�00�L '�&�Z�1����r��	jc� ����r�ՆlAin��������w�δ�٫_�,E7	���[�M��#m����� ��	��9��V�3�C�����{&��}�WL�A%[G�P$晄��H��SX���c��{�4�q�@�8�7���,�a4�1�/\��1�vS[�U&O��G(c\V/�v{}#�1�˧��D�w�1	P���p���]���i#���d�c�ұp?�c�Z_����\�ݿ������۱۱�F; �vl�vl��[kIr*�����\��CYf9��hȍ�7Y�"�铧�{pª�/����	�"���C3:1s���D^mKY,7^����t.}}O@7lJf�bU6�����+��!o�c�oF���X�{���1��I]�d�Y�|��������z�Ro(��sÆo�X��v��þn���ndwSD�m��M�)]U���̠J�d�a�V���RVL�3���$餉n3c^�]<D�B�90#h$N ,�(81�İߕ���������G;�@.Հ`�d�V�f����#������4�ޥ�q��1�w[V�ɫm��bC�����*sq:�����m��R��J�o����y������U�44��I>�����"���_�����t;=&�*V�/e:��z����t"��H��޲I�ͬKy����fw��쏺L��c9���B� B��@�b����`r�^�$�n�!ƹ �V2w��e0�-�R�� I�#��M���W����$Tox*��اRwr�ץ��G)�|�F��l��q-�����rc��Ar���{���7���P�߱?��1 D �#��ۚ��%Ґѱ�]�����6`��jW~�%2���,��gw�b�24��{0^���$I�&z>zT�V%�����@��ttD�߁�['�p��9�K�B�/����J�ma2e!||ַ�?H�21�2<�3_�bz��~G?t���Ґ|].	��7�+�G2Z��Ə���G�7���<���R�@�y��5g�'�7���N.E������'��_�b��,W�:��G�@Ӹ�M)U�����b�^�If �U���^D��Qw+_?&Ϟ�ұ:�I�?�^��
鯜�,��J�녍s�]=ި`2��YJ���Wӕ\�ڥ�)��ZߧӇ<}��G�ʌ=Q;�
7 1�)"y{���+*�P�
Ǽrq�ʹ~�Ǩʷ�I�82s�����]�&��q�����ϵ������5v��_�͋��%,���@�J�� dc�<�%ܣ��1� ����m=�J�ՙ��:2��������t��W�y`%�ED���8#`tf댾'!�����`F�|em5�'�@�@�L�w�6Lp>�_� ��H��h(؂؅8����M����� 䱎�����`07e���쵺�0������؋�����s�
�c�d�'<��99>H���8��Ƽ3v����jWs.ƺs����T6LB�#u�Zh�j�ч���(��0�9�{I�n���r��1�q��������xE�'��Kt���� ��5$���J�k�O��;,�X�朗'ry�Eѥ	$��w)��k��P�&�_��p f_^��|Q�
��M���1sw�Y��&2��� H���tbDy��ރ��9� �)M�5vP���~�ezO�-!:H.�|�R����NNNx?X���/�K�G��� �s��a�t�;�v��� X�MD �e���v�
�V�5�H�j���>�R�w ����	�:��ׄ@��Ctn���L��V�8�ɰq�8`�Bp�� 2ĊnXt �;3<w>_b�}kɽ$�c���Ș&��:������?)���4�d�D�@f`Iel4 cI��.A��2�9e�R��;�!tl����{����Ț�[���������,I��,#�W��"֨�}�ky����_��@��(nM�� �`��R�4�  W�c��	,��c;�c;�c��iG �؎�؎��~k-e�oH颸ʰ3a5^[�t>��}fR��A%�ȠI|����,9*��:4��$ 5��t���=��i
���O\���Mm�͏�8G�z&+@��ڕ΅�J�&�,#�ؤ��9"
i$i���~{'�Ef2Y��%6�ig�jGl�q�#�X#	 `u����G_����ըH�on�{������m��IޝI�7�TGb��Fc�Ԭ)c��D2	�ʑ%��9H�AK&�HL3��;��N�F7���V����#)�͜Ԉ���94�2)Y�j��ɯҪ�z0�NS]�Al	q2V��AdΛ�!��@I�0��Xu	zas�{c��?\�b��M ႊ�]%�*�����~Cz����CvW�zrv&����z+�wox^}���n�G��r��W�^�,��n�����V^,^�6�$�P�ғ�(�z�P�w.�_ȣ��Z�������-_ۥ^�������ן|)_��Hң��*[0!9��o��l��ۛ���$��|�d�V��V��Dr���t�#�����r2��!���h����x܁�Y�}6�0����z�,� �[�o��T�� �c�
� ��8o$�2z�X6��,8\�摃���P�Y����䣎�� Q���Z�ul�`+�ÿֱl�6�{�:I���c� c�%�5�/w�cT6�$��U�IWj�`�K��OT3�����#� ����QL�J���&�2��?��x0��Ld����A�qU�h�И�\�u%�������ʷ��7N�z��o%[�"�O�����<���^8��|.�J�ӹ��fz��{�����W9M�-�窜c(4���Tz\Kb]<�Ƀ�=I�9��jZ�۷��x����pV`e�.���t��˝����SI�6:o�Yd�9Ct�7V\<�sLr�C����Z��
A%�a�sPl�K�b�V����k�LjH��LD"��	K�7ٝt�SI`�N�r��N�YO �	�0x���_ɍ��� W+���~�)d�46Rcmk��r����\N�ip�H=W��o���=6����Vm�ײ�,����+9d����B�IEό84���5�] ��Ҙ�`��|�vdc���gǸ_�4������ L0f �sb�_�2 h@�����9f�����Y=pa�Iġ7P��1=��U�m[	$�1E���Gq�j�
��F�_l�R��?���{K����$���@���c!�f�G��`�a�������ɀ~	P���g��	vdf�;}=bp��F�������QJ��d,O���5J�N$�5�F��.7f�f�s�^���&��x.x �=c�B�~1������|b�� ��6�y�s_,	�bN
L��2W�?$���v�����)���f-����p��5���[�4gi�n���VCI-�gz=Y�I/'���<H���%"����B/�//=~g�}�0	̼�ȧE���:E���iu%���1/�� �ȃ">��տ��9����F�o���#G3��s�2 �m	^#�䪸��^��d@���<d1����d��獁h!?�<�|J�%x/֩u ����"d��l��7Cv7ba�~ @� �;g��s3�U�: S���tE���������_�79�c;�c;���v@��؎�؎�w�]�Mu3��z�(˾��R�:֟��1声Q� F�a����0Ѱ�_��Z7G)�@��0Z~I	�䕵7p�����!:�U�7��|���V$�c�6[V�è�
x+�`�����@����y���6�΄���F7~����u֍ɔ�Ӫ��*�7�A��;���Z�13��KL!D�u�6	} /����0-�s�d�ytX�o,9��$,�dBb,�]���|L��q���q��d���ba�/ӥ�{'�����P=��ŵW.	�Ę�����R�Ğ�'��Դ�Eb	�M��6�h6������{*��JB���}Ȋ��&�C�Lv��IAp�����
���C��~~�X�.I�;�1t��P��er2��H�轟�/e>_���B޼��a��d��>B����O(a�KM^�׍e5���������H���k��w�ŋ�z�k�ǔ����ln���y���D�t ���/�~�	���D�����Q��D�;2T��C�r/�r(U�'�.�i�N\�˃#��7��"����N�� d&H`�����M�~&���G�y�YE8%WP]
�����Z�q�r�f�X�Z�1 ���̊���7[�e���f�UY�nOw�@\ HIPT�B!�#��o���_�͔�؈�۞~w�WVfe�9�\+�@9�v`���=�vV6��5�c,hoo��B�J�w��r
�q���=I���]� ���J�1ӯL���?�R1K]��iJ+��\�!�6�299̛:4K[`ٳ��A�}3��g�>�^�~.�}%N)�Q�ݽ��||�V>~�H��`#����n�}K������C!� .��#m�W.!c>&v��E.�&���V���T. e5D���r�cSF	�&�$�d0���J��Vb}��D�	�V:�oZ���ͯE���g,���߳i$�Y$���>��2��'�4���s���C���Q���[��cz`7�L�{���Z��׵$�Pjm���Ϥ,y�����od��{�����SHx���4� ")�Z7�����X8�����Ƕs��9n�5)��$�U���W�D�g�^�u�~,e�m��?��/$�L�>[T~�Zo,@p�%�ؘ�� �h	t=h�lWK�{Wʫg�d=���O�0���V�_�
 �������ր!�/f6μ�����5�0�ƺ�|��k��-��#��8��Xl�4��R:o"�q0�9;�$��� �Z��E�>�>�MR����
��(ܵ�5�s~q֓^��o���8'�	 R��A����0Ր4Дd�b�3���������k ��X�k��k �u�`\���� ���3�1ї!�V  Eq���{XH��M欍e_.e��S&�|�2S:1�)1�p�HI�qk�C$y�~���y=ރ1?�H�v�sm��=J�Q��a�^(H�k�W��,)�x�̈́v��I$��X��O��sd`����B�Y�5:`�����`�q2�1�fq�5�ޱ��_İ�!-�Y?t~^�A���w/J��I6m�]5v��8�}RQ`|�f�HGɬ�w}*꣏��@��s4:a���;��=U��v
��s3�D��w�H^��^u�8�h����� �O��.���،�	�ݗ�@Tui2����[��ca`��vc2�lsH���މ�T�~齃*z��<?'�/4K���\��\��\~�� 9�s9�s9����P�j��	�������/~ ��ׯ�7���d�Ng�\�f�3�>D�1I�5�S��s<��`<efZ��K��q��~��}'|�����"z���s�Gl�{�s�� Џ��'A8����Nk�}u�~z��V7��Cο#POc����G�B ��f4:��]���$6uM}L%,�,A ?��6�q"�7�<4P ����@ٖD0[�����m<6�h����]��jHl��ӈ.�E��� ��H��i�g�������fnra_��%.'�_`*�gh|��h�ͯ1�~P���E�i/�i���� �՝��^6�R��;uKy�@��@}4��$d�׀�x����K�zv+I���o��h��<�/��Oe6���r+[�ۯ��(�1��j�E��N3��&�����	t����fM/�?<!�/mO��3��Q�o�g�A����|+���8�я?#ۡ�G��6R���LyO�'�K<SÃG/��"�6 � �M��Ru�>��������.����4.+�3KN��O�"�\�*�k�I%6ּI2
�c���c����ݹ�_H�����Dc�8a������������]_�Y��q3�"d���	�j�hCfs�[
W`Q���sLW�Ch��${�,�(0skJ��Y@)�۳����Ρ��;��>c$ۧ\&=���"�>�l �'it^��K�����e.7/'�B���ӿ"[��X��쌙vݗχ2��D ��
� 21&���^o&���%�e0����[	ʝ>$cb)��}8��7�{ov$� RQB]z4m6�	~$iM_�:����|�P��� ̌�$�¨�u�&���J硞�Jɾ���R>³@�2�=�t��w2�
�<uؕF7Z/�ڎP���#��"�y`d�+��ż��c-�w�/�������3��X�k��}qH�K�c� ^}5�t�HVK��m%sm����`<,r��H����t<i�%;�G��H��qp�~R�3�*���b�}��[�sY��L��gHpDfңC-�jB:w��S���	Ϝ��S��7'`@�ߘa��������@�	zG���!���ӱ��Sm7q^pI
�9?��>K Ht�~pǹ��E E;��kS���6��d�"����l90(�ձ�����c~��d����Js���ۂ9Um +p���c�E��l.�LLʥ���s���r��B5��z�5���� ���f<�p�s�vܪ>�)�>���c���ǹ��=0��w������\Q20 ܙ��Z��  �Ȥ_�9���#�н�GF�2H����9EV���Ǉ���Q���{>oBӷ��]1��������{?hr�^J�6v�����q���o�`�Si��e�ĐI8��+�c����@cG�6����k����q~�W�=�!�H��]d/P�F��"�D���P—c����Ԥ_���Z~��|.%ic�D&)k�cL\��w�����	m����\ړ�$�O��}�YMv/�2m|����*�DI�d��OhB�g��7�}" �x`��m����������r.�r.�r.�����˹�˹��?���&I�<����������7�|C)����5��j20�l�L&#y��\\^[�R�f�F@� ��$�1Ӵ�ZyЍ������o�0�Ђ`@c�= Ä뙗�˻s�eFiu�{ւul��6�t�oǽ#�2R�w��6{�s\o62_Υ���_$�7�ޝ �vgA\�1B�_l�P:��Θ�ߓe�c'hY�ބ�0@�4���g�6� z�h�b�h0�&9��P����`A'fʛA�u���k �����]� �5��Z�40��B@6I+�f��h���+�����|���;��3�!�#��|z?���'K��˵<ܽ�w$e^�?b�	�D�k4�v0��'袷�s��|b�%���0 s��h�lݢl%�O�m��ه�lk���R>|��������,��/���}��"��l�`>�pr���?����w����h��6�y�.�r�2z��~�y����j�u��a˧�TT��]�����|&ː�;���hZ~�,< �A	���W�����{Ƈ2�3/��c<�ğό�����W9e��>������\���A��P�{N�I/�����h�	qղ���LY�{n����y<=�G�2^��I�'�ȸE4�]-͑��}>(g ���T�L&��6�y��p��N������{��e0�E4d���Ǎ�WZK Ez��[��~|�s��/ �J��ܽ-��ޘ�zFYcaH6h8� �D\��_��"Ϯ"���FPj�����׌��|��[���>�`�c���=�v�6��M!o����or�xv���e$�I-:��>0W��/X`ՆF-��`��_:��Wڏ"��(�K}��Ф�Ň������;�o&S�?�x�S��~���P霽z�� ��v"�l+Ŷ�G�p�@�X�S��.od�ׇ�
AV����f]ǆ��N��h[ջ��õ\>�z��r��z��M'��d��6�R揵<>�<.��L
I����^c'��Ij���#:(�@�6J]�!�b}�u���<�� ���Q�r�i6�;�V��g  ��1Y/u�ׅ�[��4�N�g(vR�CmD���$�K9�,������ ?9r�e��ryGˢ�����E���T_k�5v�B����< k��|"��?dTe��4�j����D]��0�-@�j̡�e�#�O-op�E�s�tzAp)�w��(9����>L��6qh�`�L	�蛶��ٓ�̘�x� �v�9�5I�Y]���a�GA�1�V�?��ɵ��=-�:l � ,M.���R�={F�0�^0wa� JIw���?YZ��It��d&�|��B}�o�_ X[�}|�ͷr�᝾7mɰ���(v�{���<7P��̂%���`�U�)�&�_�. �����33�L�P�@�0!m�{6$��e�s7hq90-��$+�ԟ�1N9�y���XM�c&�߄�u��>�.R; �)Z}r�O�o�+�}�fÎ�e�'^#eG3���1��ޅo�d��$xhұxBg�m������x�ØL�
iB�F������}��'��5X��I���ox'�9���c�k�LB8F�ȹ�������s9�s9�s��.g �\��\��\~ВF�-��Ųtyq-�7��'?�������<��F��߾f���_0�PT�a����H?�B�����Y_2x�LPÐ�o���R
����_h�c7��(��p�Gx�/M�<�S ��}$7|�t#���0K�G-������8�@����hb���o���dWZcS�kPz��tӚp��ex �`��^��x�S;Y��m��=D�Y��ixj GώڤG��&&h��9���7� <� ���	5�i�j�  P��	冨���C���I���17���Dԁ;�bh��s]��	0����Q#�� ��"��XD	�?��^>���GS�LGdE�}�'����#y�� �n-Q��J�׀���f%�ѐ}�F�9��٭w��H>~x�u^�f[Y�����wY-w��򛯿���9��B`���u_ɻ����������濒��я+�d1�@Ze��Ӕ��ﴽ�θ20i|�����!�AANx���z�L�{�����K�� �Oh���m^/M��=x����M��O�����N������OO��C�t�����U�Q�8���`d�$9�.��y�˝>>�Ǻ��o�3�?����o����!oW�;� ��0�̭���r�8�":_�;A]`��l��!�h��:/�g��X�f�B��Z�{#P�	 J�En�Gr}���+x�b�꩔�"O���g�X"�4�̨�� �y���p/w���X�w�I��9m���7H|`$�v�h�E���3o/�W����%@GHc�m��ߔ�'��R���X��|8)%���Ը��zEpl�.e�V�a0:�DqM髙�c��B	Ý��e.�pM}��O8	^J0�:E}�A�`�X�m�F�t��u�>l�o'�qf��~�����s���dwo��n��O¡L^>#�F�7��wҋ�z~�b�k���H*�aľ�������"n������6ӹN��>`v=�)0��@�Y�G��!��WdJ�YF�|��X�3��@�D[���TZ�6� @�' �����{*�����9��`�0��8'�]E�]�	/���ȪrL�� ���F��mر���v���P�I2N����E�DG�"�5�`^"�Z����v�%���[�����1�8Wx�nM3�ω�`
��[�0G�������Ɋ]N��ǼT�&_ �̱@��~D.��t2�
������?i�ٚ؜ ~|��g�k_+h.�3ɲ6��ļ��<� ��Krf�=u�F�*pD>j@y>[�D��i?�;���( �Q3a���^�Aߞ8
\�a�g:]/t�-P
�@?	���μ� �>���~ F�%��nc��U�c^�=b�\�kCr�DC�������8����t�V5%��Ԙˡc\tڪ��cDI"�ȑ=�u�:�����u䈠������# ��D���ڽ�^z�D�#g����'��vi�_�qvF��8�=��Uoӽg[RR�= |\p�Ce ������<�Y9V/��	�u��J�Է�\��\��\~�� 9�s9�s9��4b��ˋ���!_~�3������@�|���������n�)(��\�wn�����5�̘��JP�?`�<s5u�:�sB��BJ� i􉦱�z�7؍mdC9��X�T"����/�g�;�M^�FL?O��X�,���L��N��a$/BFb�8�<�c~�w �|����m�ϱ��k!��P�d�6�J��ʀ��t�� r:�vh]�����G��w��@�ò���|0"rF����1h� D��v��x��� �'�w��QO����#��kZq������BÔWp��7�'t���Y吂����'72�]Qn� ��H���b�,��Y=Ѹ^�������^�ry9�@����A���7rqy#����G�CZf��:/�� Y��}���������A>�}'����BƓ=n��P����=��i)P�*���:�TM^����[i��fS�\`z�Jӱp8M��=��QQȲD�dKp*a�4�96����ZJ�E�(\VsD��A�� ���!*V��ٲ�b���wD����&�]dn��('$A���d�yd�}��ǩ,ש����bt �N�"7��C5}x����x���-˛�������@c�e�3��l���z��g�X�Tۢ����m��}B=���z���]4r�R�	�*(6����aN�r'�v+��N6k��2e/$�����˘�E�"����L�Y��\<�˔�Vz2?&��$��g9}�U�O�]Ꝏ֒m���ھ��Ӷ�p g?�1� w���Y�|�L�ml�/�g E�ڎE�׏d�X���R�+��v.)~�&W_�^V�+�����(\rT۵�>��e����5X#��� O��N��:��"�ojyx4�.�0�r+��'�ހiu���1Ri[&ږ7�L2�3�Z
��@�#��K;����]._}�HB��+���s���fQʟ�կd��K	�C��ԛw��5�Y$X=�kiRy\�r�>��ܥd=Z�h�'@yҀ�*� HX�'��D��x�7�;�\�urf�Y*t�R��S�������z#�V	-�y�u>�ƌ��W��}�N�i�L�0 ��!�drX 8�IT�Ҳ�����/�GYL���ƌ��X_���������˂��z��1�<��q2���t��ɧ�������A�Q燔��RS�����L��p(�b�U$L ��d�����d�(��y�k"��yZ ���F;�>(���vp��'��%�#z�D��Pׇ���ŋ2 �b(�|���~�VV�D:���3�ٖGOɰ�{����1� ����`d̡��4�#�0&��x��e�14��<e�T���i�l԰;�3�q]@{�ypr���שj��E*҆������T������(G�rN%�IZ�A��裱G�N4�9'�y*�d��ߵ@�@	1�/�!!�L	R'7I�#��w��-N1��Hr�O�%&�*�;�
 �#�%�ԿϤ�J��c|L�0Q��{W5vI�u������:XύS��B���͠�}�Ԍ�� ���s��y^��υq8�YR���ʵ���@ñ�$�$����s9�s9�s��.g �\��\��\~��� ?~�˟��_ȟ�7av��!�!noo���R��ßp�
=��p$� ��Sfx�tS�M�`t
p�IԖA
�~z�P�NN@���bc�^x�uYl��Nu�u�|�r���Ė7��z���<c�6���^~_E�2�.�,�)�Q�����]Fj��h�b�k�{#n*�<&���C.�e�PX"0f3�#�B\P�Ad=VU`FiNd� ^�Ȥ����M,��9��7�@�9��M[�`Fj�15��	���d��"+�'�IO�g1����N�e������=�3i,���N��k�3����r�6AF���Տ��g��L�2�'{0�ٿ������l��e��ӗ�6a	)!�M?~�?�1C�嫭�wy��{�/�H�4R`"q���]�Ǽc_x�����L�P���_�T�.o�%�z�.7���u;��-���˲D�[�ً[y��Z.f��k>(d� ���et���)#�3$�\Up��v�N�Er�oϸ�^���4��1.�ۛ��c��=�䔉�z���>xe}%���G���_p��j�c���i��黗�B�2^8/�	���4׾f� >�.8����lm�q�pE�z�RYp�^L���ZW��j)�US"�K߹�}D�c�G���b�x��|%�yɀ��b�ȵ�.�(����Y�ғ}���]i���R$_��k0�Ĥ��`_^|�K)���|\L�K�_���!�IN����4��/Pw;�}�4/���7�R��$�t�3�7�)e��dw����s�ۋWf�>���bxN  ��IDAT9��&�)�rAFɔ�:gr��qN���[d�_���SI�&�Yi}����z����)�A.p�7��-e�^I�k�n3��*t�վ5H�k��&��C Ȍ��~#���c�g��Gȡդ���;�k�������B�K8�k_�6REwd�`���R��T޽7���$�L�v��LfF���R�Y��������8��4�_@%"@	2YNn�4���ъ~!�-oke� $C R�Z3:o�`�񵇼��S[H��q�Pr*�uc���Vݜ��;�,w�{��y�+h�S^s� �ƹ͛�e�'Q�=���,4����������DN��N�8��,�IY�$���EI��3��{Pr�U=0�w�A���Y�9�/�`�������8J�7����d��<���?�D(؟�~�����j�k���hH�Ap2��%�<�d 7�5}� �w}�k��%���7	:rHiT  ��[���&��䓢mF�*@�C��;����=�Bl���qޮM&r�|@`d^y�L裰��Hq��p�wk���0)&���dx$&;�׹~?:�����[Y�䡟j����w�6Ǐx�� ���d�S�rsR�5'~�j\�t��#>^��[�,��A����uT�����1JJ9��yF�?���[!�9FUL0��G��I��=Z�nG??��{�t0�j�<->���ĵ�%*�x�����p>'l��!�qH�h��GL��ҜA�s9�s9����˹�˹��?�4G�Kx�,��vEى�t�`#3A���襁)���ˆ\|�@1��Q.��Gִ�q��c��  7���t��^�q��MY�܀BN(�] �m�xxYw�6SɈ��f%yi;Yl*�"��glV����A@���I_�=BM0�Fp(H�}��;I��I��$"�Ƒ8g� �� A�����f���f��TH�5ZW�>c���"$�F�� 2b��fJ���:�"
L��oh�A(���%������oY@��	�3�`sj&ԭc_�H5x9'������yn �mv�&���l5̧%4��&�-h�m|ys+����2��X�&I^��8���|.-$��J"�s �����背����Df�\S������d2}���B�!���'y�����4C-��fJ��q(�;�~���Ӄ\L�zݖ���g_���R��K���^� �AY��z���/~�G�?����������33�mČuw��;0���edN�}��k����D�ļ������C�����ޠ���I˶�wY��;w�}�>�p����:�Aqv |&���� ��?����&����i���pjh��K/9=�A_0�wY������u<KA1�x����\�T3����V�,a�?|spD�2J� �ZoD���P����zh��p(����o�����%�(�H�j����;�~��C �=n7�m�$�-��,Y>���¼hI�d�M��W2{�R��Υ���ޛΧ��Q������έL�G&���!���i#�"�'����v+���e\���^g+���xHrMx!���W�7�#�^Gdq���u�z�\�/R�z�ymr.�Sɒ\�v%����2��#3mG�u�y������1^h�o(�[���\^O%���'{�?R.��N248�W�n��[��M)��)�v���X/�~Jm����zq�*���6�G)76�)HC���f�C�v_�[2�VZ�Í~lY�A[�LIyC��[�k� �jB�4��]Vvm/��``�����`$��ytG�=X ��9�O�\��Zכ'�-s]st����Р�V�{�� �Xs-k[�0v���k*���������@}���0X�q /�Sq��#xO��Չ?Q���{?�D6�������G?�PJ�l�Iz�@�g�����u��tXA�{dc��W�#������`
B�
��8/�"|m		��vh�₰�S�!}���ؘf�����u�����f��\_�{G*׳+��;�K�6��$�lϞ_���5�JF�1�	[r-A	;���F��mW����!|� ��Y��G��u<�#�'�Σ���p�`8 �	l[�a)T�;F�#���8���d`����2(֍��}ރo/�g�gj�
��k;>=ε������C�g�n-X���a���a�|DB8|�/P�	x��yY!vc�a��	�I�d�j4�j���o���G9�Ss�@���K�^˼�>���*7�q� ¤J���z�1�o�u��[sH�*&��G	��*�'8��D����1v% �ݶ ��H'|�m\2U��`��.%��{�u�#Md>=�>M�Q*�S�<���˹�˹�~�3 r.�r.�r.?x�f&����^�O2�θ�A@�ݛ����7�)�QG�xd%N'zܥn�������Y�;i�c��d2#k�9Xv7ˌ��A���/ȱCp D�`�������U�H�ZN/y����A��$�5��/�(�1%�['rN��Z�H7�&SQ����I�&�d&I���t����n�?O���0�,�Ӹ�u����> c�e��+�	$�$� &�wC�u@3z�	�?���Ny�ד6C̦B���s�LV�opt5v�uʑ4���=4���(2���[� i���&�#D taN��i�hɒ��=�h�7�՚���+yZ<0���/��B�	��쑕�%I6tRH�,�\�,&s���A��$X�����%�O�7_#�|������ϟ˅��7�[�S�O)����l,� ����;�˿�+e�k0�\_�#������hx����|  ��q��3�-�Sv�97P0���8N�LF�27����� ����=?NY*8�#(=h:����e���/>�4����b̐a����������\����C6�u��3�l��u_���:h�C�����ؤ�u<�,���)���Jd���
 dmb	��d����L�v%���ݦ���fYӳjJ`o �^��&g�={�m�`=α3<&����|+=��f=q�5�Ɓ�x����6;��v#m^r�Y>n��=��X$�@�DLSñ#H4��y�3w]鼲�O(O%�$������������Y`*�Q� @9�	&,�f�+L�%��lA��-e��;	6si!#4�F�J�y�bID@2���v:�u��#�k#��Gl ~�G�Ty|��e����V�W������(�Hh�=�_`�+)#��*�.�k]
���/9����m伞�ʮ�����e��v���c]����83x����c(@6ϱ�p,�G�/(�Җ� �!!�dx2փ�O�n}|0Fi�]I��y�8�D, �DAԍ�#�js�z���?yo�$�k�}�r��dŁ���q�n��̞����J@4��	�u��`0��PF�y�Q��ݝ��L<��x^�!��kY����_:C����������4���L�x��V~�_�x_�����^^������� @��v'#�,�!$����1��3� �B���_�t�1Fʋ��9=��4&�v�m�}��5)l���ވF,��sPc�Y�Y�5�E�G¤
?G�Y��
ߩ���׾Ug��w2kB�M������x�2 �����Q��:��rB��| �"�s<�a`F�	����p��OD��S�G#�c�/�.��I<}�pf�����ab�ux���|�*�[���^�+�m���~B���� Lr��hC�z6�:yJ2�q���¸�{�N�ò��3��ז.!r�j�����s9�s9�s�S� ȹ�˹�˹��)_}�7�06���<C*߿�����������62O�Ff�x<���B7�=9�-34��.tS���_�/�'2�\HO���ݎ�������fC��9��t���X�;2�u {�3�v{��:#�W�xd2r������C��:����J .`�L�;���׍m�aV�|A�YƑ<�����]��=O��
�Xi��F6ulBD�/�P;݌f����n��;� 7B, ˎ�����š��� �ѿ,��T���&���N�$M,ئ�T7mwn�)�r�"��h�5�M2a��p�"����u�:����� ��2|�q;��Sf�6��5�ȐF���L��b��@�O���NJ��5,����kyZl���5����Zn���@�D���l�e:k���L��n��0�>�e_���'�y��a><@j���������+?��'l�W�>'xv��#�~K����kJ�����J~�����}��\�-7�b��iM��e���A �)�{����.����;��S�������ϸF����)p��A�4M���ऍ��@FTX�Y�<�!N&�����%#�{XY �B��|K�+�,զ� X�,��\_49y����F&���$�].�����<(�:\J࿢�h8��52n�D�� '��`R��NE ��$L[�(Ij��"�&�ɚ+d8,b`��od�^��t�A*l���"Z� �֩�_-%_��;�J�[�o��cB?د����"{���M�\v�[b:�)�FZ��� 2 `L�"��JF��R�����Jyz0ZJ������(W���#��n㚀Y�Q�f[�����o���-hs�"7�L6k4��g����������U-���?��5 �F?/�#���\ʻ�B7Z9�R�?���Bp�z��ZO0��6����%��, lF*��7%YN9�&��͇���~䙎=��{��:v��(1> ��'{�M
�aH����ã\?p�m
h��t�j �����J�k|k��� �4���J���W��?%q2T5=)*���0��}2ڰ�|8�C��Ax0y#�-�=�V�`��nKYC�Y~0�c����}�cn.!��ڃ�I6�;��ρ$��\��Y��q���g�t�VNr�_l�!O��`*������(˾��^�z �Y�p�=Z��[��@�z+[�� l���5�(���Y�G�ν�#a����l߆�TO� ���0<ceA��X���?��������Q`���YQ�����21P���>A 0�8M���j<S��B�J�9sk�/��vqy)�cO��k�w�%���x���%�e���Ǫe_d}b����wc:`_��[��O�>���#��ӵ~S&�������F[�>q �A�sje}��#m#����Nd2��r߆�_$�+~����1H��HmRW��%v��q q�A��х"G�{7�{%^z�H�gG`�y�I��^��{���7���A�\Q�1������N,${��۫	KK2j�ԁ��<�l�O$&������mDn�'�	t���{��)<�L?N�9�s9�s9�s��.g �\��\��\~���UD�U+_�kNFr����ӣ|��o�?�ǿ����x��Ŕ�}�?��o��u������J���\ͮ��d9_ɻwot��(�rg�4l�K����g<����k�mw����q�28O��w���r��'�v�t�S�ڤ ��33E��F"̬U݌�ھ`����X4p��68`����p��s���e�|�ˬ�N=��7f��y�j�{)��g�JL���K&��T�I�TN߹r�Ct���`d �v�I��N
	߃<AXb��V�d�]���1����軲�������1;/��4�#�A�lD���v� l	��U.�O��(��0��|C-�����&�1�����j���b)�~A��$�d��$o߽��س@�4/v����|%���^�ӛLe<����5��W��"ߑ�q}{+?��O���-3��}��x��+��O~,S����W�;ʍ�MAl�c�s���|���c�v&��t�V���Ll��y
��w��1��$�����3�=C��;ÃUe�R>�t�,Ԇ2�/��y��k  y
�x�����d^�t�5}���������|�\�o>[��/��|������|A�u�`���q�>K_�v�,jM�`���@�Bt  .���"x�Fh\�|�N.�g2y�Jϓ3bB 4L�%�f�o�2��l$7�'+����}��&j���Rf�c��5��L�R�j�CB.�T�t�����31�M��l�\���۪�|ef�7sd�^_�����H�Ð̍]����38�f�x*��c�X_J�eC�˫T��3>��@��	Rf�'�D��a��݉| ��K�jT:���꺳)���t)*��]_�
 SN@�`d.��֙�,�W:������*`]��Dؘ��Ph�4���h%�i$[���4C�V
PᾸ&����zcu�z������u��"�}A�
��:6��Ґ3�Y�E�;�Itx��u~��6�R�w�F{��:�z]_l��b 9<c]�5��Z1�i'�Rcƙ|���Ei���O ��r�i���ǟ��ĭ10G� �qN�y��"~����?�����#�tc|�^�����0�eHqz���d�P��uL?��$Mc��R}����K�̫A&\���}X �5`9p -LУa���/�u�:c]T�r�������ɾ��۷����4��!7�U���g~A�?�)�lx���L!%���ь��t�	Z�1����R���~��uN_��xHi.�I��A:B&�2���4�����T8�Ս�#P6k\ml�#���������%8��U���d�|j\��{��q�?.�,5�c���7�/��bu�)i�a�pcl�O�>���	6Q��� G@��4�ѣﱥ80��!�m�Sy��0w�|�$��#v����͎r\��ؼ��+�5�	@z4b݁�1�:�s�qt~��&5���E����{:T�ce6�.:�l+UE�ov�7�c�}��Bx����U���19�����������˹�˹���o9 �r.�r.�򃗢���dȐ�z���_#��i��������_�!����\Ng>b���e�-)��d8s�6�|x���������˵����]��5(���&���Zm��26�Д�v�@�%c����������rf@�d0��N��m=3xsdC������h4��96�� b��ld���@��e��^kD��wƟ��/�3�ߴ�y7��i9�Fv�N�,M���tC�~#4˅��>Md=�r��I�y�X��8 ��g��4>��0>:%�#���a3/5�`���� y�A
�H�@����dWl��#��E�h�f�BFJ��Þף�p���,O�·��F��t�Q?��+y��&�S�B����X��RV��^G{�`H��db^h�uoÌ^�����E�&�;\kW�?m79�b��,�dzq%�_��s��� ����cy��\\_�����Wˋ��e4� �fIMɏ�ir���#ٷȚ��������e�bg"�@R{��B?�k�ksvP�x�� p~.-��ɹ���*��	+�* q�$�@0Y�ȬFP�%6��]̀_��� ;�Y��3����g)���@9 ������x�82�Â��<������ ��PG�����jqAX�I^�-���5mɠ�����H�� ��0�OVNd���Y8�#3æ�Gm���,�!OG`ò���w�]$2L�	d��2��!��I.�/ 6�������k�k���k�k)ۥ��tNK^ɮ�����򥔽�Tţ>�V
<��딞 ! A��3^�%�Բ�G�[�\��I�@"
�/���R6{���~9�5چ[ëR��X#��6�萔˛L&���懦�|�SJ�� �:��gR����[�M��,a�I��Σ%�s�.pO��x�ɬҌ�#˥��-|	"�M���B��?��ŏt��sY�D��2��*g[e��L�S���i��t���]�a��t���8��G=b�&��S�����kno�yG�{�z
0�j��jO�>L��ռadr5-��56c�@[�ۣ,��
���������d�`�q����-��v��GQ'9UP�I 0 ?7/!���6�Bܼ��8�US���y/ч{��븹��~ ���2���<�Ys�ۙ<V奻0,&��sb��z��Q���x��X��˾�'�}0�:�>�=؏�O��mķA��=��L;0m�:�:� �&92�g�k��|.?��}o������ۡb�³Rn�*�Ɓ�5���T9Pj��X��A!�ĊcAj �eA�U�m5�����n���~'�z�k׌r�	�Cc؜�l���n����*n\Q�〬и���������5�S�ֈ�`�;I��ü���:ad-���=�5LB3�׾����g�����[�sFC�wJ�	P_<���G��(������@|ҁ���ƁK���ht�|؇'�Yx
���� b�����~O=0��hh��1���٤����.�{ڍ>`�V��)���U�6��M*���� �0^��R���w�b&�8C����K&ݸ:��H$:���\��\��_D9 �r.�r.���f.}��|�o%��,�o6�����n���'٭��i	�� ���f+��Nv��$:h>{�]��]@�b����ߐ�,���{f9��;lqx�!�;R��@ ��Ehf����~��ծ⣔$�M��.��#h���n?$h��t6��Г�zC�sl�!k�g `b�ꖙZ��}0c�'���Yp�d�-M�{`Ř>;
���e�Ӥ��Ξ
#^�gJ/�ݎY%�ࢎ�C|�Ghjf'N*�m���wAl�&θ4d��Pj���N��D��y��va�q�<��a7���@jR yl�l-�d�~�}����d���O�Xm0p�Ȇ��Ç'm�	��^�m���c�@���Q�>����b�:�׍�`��(3כ�^cGs�r_SQ���EɬI<K� �M|/	<�z]�3��z�cH��8A�,%�"��&���� m'/el��3��Y�^�3.�d�g5��-[9=�������gP�� �Ƀ��3#N��T�Yٞ�br5��G�.x�z�� �뿞��[��Z���s�x�3�����0��-%Q�s��c��ཷ�yX���^)��q0��{m�=����$�nH��WEK�*vD�Ǻ��	Qx�@0����&ņ[� A$�+���G_#=/�/�2��2�m��@9�O	�>��F�o	z���"�p+�v��B�홎��Z�Ϥ��ۼ�����֓�R��e���s./e��~�C/��4�&��"��"ϟ�2�ٓ��v )� �"��;������w.�S��M���B>L��|�l `l|u���X:�Z�z�3K�UNl�	�ANI-���F�3����ar�����Bt���,�/��D�/����n?�~7�d񸒷�6��Bs�Z����nDf�F���H���,���T��%A�m������2y-�1m�BO�@�y�(��d�`y����&V��	*3V��?gĈb��F���F�;�'Z�I4�:� <�^ڋ��md�غq�1H� '�Ţ*:֕���8� ��Bp��h�౓9��= �Y���������Xw ��=�,t����|�e�< �?~�n���@�YBMu�p>?L&R�\������P��T�o2�x4�k�s�tA����j}��x��,ƌ�y�M��[�(5�;�B�YW[��x�MF2_�(a� �ݳ��l>���V��-�,�w��n�:�t^��k]\1�18�y��r}9�9� Ȱ��w ���5״�Mv�.5`�5�0��a�e,X ØӨGp����ֱZk�1���$>�`�v��(�Gr�N�n}I��`Cf4I�9�lG�9�uQ�o��qu#��{�+�	�	&����f�)_�w����{%:6Ro�^�0<k;	�����(�v\� ��xH$dS��mB��̘��W$�l�;nDЮҾf�����g������u�/��?��)���~���@�?:o���A���d�j�� ����8�ڧ �_��+'��\��\��\~O� 9�s9�s9�����ƪu��>LH������K��Fv@]�����g���ar�M�Z�n���%3P7�������mS��3a���m�� ��,C,P��<&r?�C���>(�)��caҘ��d����������Cn�	RD��gT5%^($Y�g�Ξ��?��Pk��/˨�~6��,`ո,~q�Ge�L{4r��M�� 0]�TI:�3��A�������}���W0�Ld�L� �=Vn�}D?-贡�����j�	jAk^�0|G@B��A�}�D2���%e��W�7� �j[ʻ�Or� Cz�������Y��Ͳ˗? ��QPA��Z�>RZ��;��^����Rʪ�b��͐�ڂa��il���$�F�[ٮ2�F~��\���3G!F�oM����t�`�^�Aj�.�o�Ʉ�Ӡ������4؃ X��b�qt��:eo��)��)��'�z���s��'���x�羏�����gR��V.�����|f7�v���uS�fn`�&փ��0����2����8�m�1�}?��N��?���^w�t���l������v'�a��OKY7H�%�cqQgJZ! �X�79� �LG��&��D�D&�d&WW{i���/�4(%��ެ��������Az���eb���F .@�d�(eve����b�Id��e[97����ю��Z��?�g���ߦ�c��5��pn�z�`X�޶<{ɳی��kP��
�s�������Lz�1��߾ �#����:��Yo &��.�˾\%7f�(�����f�=��2���:nk*�|���x�m?�@B=����8G沮i`N?�`������G}fm�z-�ӗ0�������]�9�����Y�:��~)����	�;������W:�¸~/�������#�z=W6��iY�bm#x)!��y0�b��|�0hPf8�|�ڙ����N����f��ӱ�x4�2��>g��f�,�(��d�|�ǅ�Q�8�Xo=�m� ��pJF�O}u����FDi��dtp��]>H<����n�������W?�;�3HG`�Mxc#�����V90$䱘kBa��&���Ac�����TJ��ÁI6ǰ��/	���Y�M�d�����4��<#��{���3���W:�K���7z��	� |N�
`p�j[�%_��9�l��z�w6��v����D���� 	���z���V�Ow&����~ᝩ0F�`j̫������Ϳ���ͽL�@��U�u=������8�o���x�X ��y0N��u����j\� ut�cg&�1gh�eL����Gd�^��ԮC��Ds�G&m���$�o^�#Kg�.�YDd- 1o{Ľ����|W�.��{:Ƴ�X]x��RJ�V��З�A�D��I;k}G���i�;,7[�@�,"[îg�yĶXW3��~�q	7`��S�\��{�`kZ��v~X��8����"(rmw.�r.�r.�����˹�˹��^�0�}� �VF�Ĳ��TЍ*��[݀�6;nv�1u�sc`gٜA���@ƣ�|� �EN�l�@�ǎ	�|�2����ҡˠC�U����s�7N�)Oe����/;���:H��|RhA�F�Qh��.gP���t,�g����|B�(�l�1�gW,�Z��9MM=�0Ёz����M �@)ӓ$���b���q�@C��c�jx}if��H�AՍ�v��� ���0� ���
NZJx!��e}�� ����W�:6�Am뤓��	S��� ��.����{��g/����[�!�`�A|L)!J7�,I_ ��^�i�]^42�����cp��B6{H��d:3��\����3 ��S"x`����"!�����ł�0��k�!��@62!�K-�� #����=A�/�I���}m�iL`̔��Sy?cjԲY�wGH����������A���0.p�5�Q|64���,���9��8���Ov(��� ��cL�������q"z����ǟ0-x�N�:5 ��{Sf\���A�p��o����x���֛�'���|�� 㜁T �sI�t> �o:IC�qAǐy��E[�-�gj���=I��郘��I���Akv%4No� mD��R6��T�k�w�T�QMy��>7:�wB	���9���k��{1ːS���X箏:/��v��kȴErs;���\��f�u�}3�r� r��j+IS�`�N��#fAf6G �R��Wa4N��y0��}d��Ier�o}6Ȭ�
}D�-�crY. B�z�=�������/G�M#^�̏E$>�@$�d<�B.�}��ze�P��_:G^6&�6Y<�#@3���x����T���O��߉�Wl�&Z��ܿ�����F�ɍ��N�b!�h*�����F������]��e��9�>������`�D���[M{]}.������I?׵��u��`W��7��U�s��b}-�E�g�1 ͼ�y^� =[�pR2C�#ä%8��2d� 	�q�.�K�JhZ�.h?����Ft$PX���*+���j�؟�� �A|`���d *�F1�0!�Ḱ������X[�t���H@0�9��z�ya����.�\�.��K<�dL�#w|t ie�?!��<�8)	p��z��vE R?X'����^���of�nL3c%TU�X"{��>���3J�ÞL�eX����Ņ��;�3��[]�6�����k�R׭� X �	Y�����?�V��k�[3�1��(�;���d|��NjQ�E�4}��}?�oYG~�O�dfBv��맡�\��)� i	>�����N","#t҃��#�F*c�&���P�Ű�G����\;
:���(3�w�^b��+m0ɑ\�7��ޝ<�ŵ��!X�D���Ŀh��JcH����dmUf��NL�$�����*ݟYM�O�&���Gn~�M�U�B�DY7θ��i�%&���qٟ�u����|���;J��i{i���F��.��L��;֖��Pl$�ʼD� c"ulJ�:!�F��d�mH/ �^�%�?a]�D!���ˊ�SCV��wFVd@�ɟ�������vo���]��\��\������s9�s9�s��
6�aEP#J�K�bRi[	��s+3��\��
�����,�<���7�M�z��b����l�Q���̘Ԉ�\��e�X�Y�=��ko�i"�ȧ�����OiB	�N�Mc��F�y)$[tC�,4t�9Af,6�{<��NxC4�8���L�qY�4>�� �[Ld��~o�u�Mb�Ɉ��`0����l�`E%���Ġ�\�"f��@�b1�d�u���2��c��>���+]Vd4�>�净��=�t��Z��Q�- ]`r��s8�Yp�&sQscˀ:���זq��?��+���rz��,A���d�#�����I@�2R�}�6z�������w���?���k��B@�d�����Gy�?Q��(0��.��PU��c�b�l�7 �2 p�O���Ǒ�F�	���9� \�0�%�� � ��E��%�G�#���D�a�d��:��b @y/���;� � X$âϠ��AY }�,w8�;����a�~� G�f��g���|�3t�0�sf�a����"���Ì�*�T�{����Ie}@�����Z���T��rs��r0�>>,��`d���7�; �3CwF�>S�C1�p;>H��A�.w^&4��s#�ی��N~���:�ĭ1�wI�t�Ŵ���uo���r� ށ�К)F�D�0f�똮�x���	1�,��00H���cH����WR���|*e��iD~���f��l�[�+#��z��vp!�q$޼�����$�1������}�9ds�/�f�����5��q&�k��MD���>��6L!��+wږZ�Q$�7CmS�����E��[S���7o�W�3��l,Y=��=�I6L�����<>�<=��������ܭv�k��V�ہ�ͥNnO"ÃLog�R�
�0*d3/�a����Sb@���s�16�ٯ�H��R�T����b�^�b.�w$�H�Q�K�T)�����W�{�IKe$�Y啼��n_����dr�J6ﾖC�5�` c���nd�ث��Pc.�A3d����K���A���$I�l�Q���u���8j�U��4N2r�@z��aW�$��ً��Vf1>��>��Z��c�#��12� f ���eظ���q���}��G�*J: #Юu��G6�[�~�M����hd^U9��b\k����-[�\��� u0��m��B�L΁�g�3m�ԏ�: 	 j 6\H=1�� �9d�c>!��e]�]1�0�̸l� ��9o��q���?�S�z�����Rƍ���4�\�bc�]�ȋ�/����xK���A��GF���ӄ��?ˌ-a�_?trQ[{0P��[�����DF�3z���<�5����Լ��Zׇ�����Z��@�PI�
�8�4n��|�DH�y<��`�*=�~�fC�3 Z("ο��)M�
L[xz`�f� ���$� 3�;
C��^����9:~�N�Hm�V�^��
�I	R �y�1�"bR������p
�����v��oI��}E�G��,�VLƵ� �����w����O�ᨧ�bh�qŁ�o��Pn//�Dz��:����m����wɋ�Lf�)�"J����<�ObR��iP�|�����b~_`�ژZbK�:v�~��p��>TI�m��@���j�9�&�)$J���S�\��\��\�%�3 r.�r.�r.?xaP3fn����O�iA�7|��K��@�h���|0L���Z^�z��	�QF�!֍��������J���������(6�C���2��u�u�q�	�0�&ZFsQfd�di�ٹ���md��	 3�
*�H�ݕ�Q͘�k��z��o��36��K�o�I6��w�������&��v/�܂M�0��YJ!��!��Q(���ֲwNn*�������m@ �W�m�~$�*���M�KQ�	R+�� �d!���f�:�H��y�Y�x�M�ӭh(1RS�� �i�����^�>��c`B�,tKE�C7�`� �̣0��� �7	<!>�j���rN�LUn�m����\N/e�|HU!�c��ɨ�5!���17*�   A�ǧ'y��-��YĈ�	Adc�Lg�����^�L��|lv�5u��Θ�uWOz���B/�����½��虡��w ?4FP�i�������T�����rprV��ῇ�}JN%�,wp�c�A@�DN���X�a2�0w�N�2�X�5����/�Mh�/]���v�ns'��tL��d�{Y�A�t1����Ӱ�t�4B ��V�/ ���� r��^�� ��:���,*��.�&������f��7�~$kA��/����KR:Ond���$���t������^����"�Q/��=��٪m#��;+�W�_H6��L�zP��sN�}� ��S^��S��P���P�=�$ܭh�{q9�><?d+�Qk�KҦ��(��V8%N�)4_
��kx��$���Z�E����\޼�E���3�a�.�|��]��? �YYIxH$��3U
�1�U�||_�7���� NT�/Ki�<����õ\]_K0��3�y�i+�zN�k `�?.kyZ��� |70� ��Ç���4_�/t�}�sZpq!��R5R,�z�����<n���#���	�1@�LNh,��d2���s2m F�b3�oۜ���w�wmRZn\b��)���p��/{��,Ir�������ۺGaf�@�CP������������.H��`������J����Ȫ���T.��nUefdĉ�s�c�L�������hC�z ��RU��x"�`5�˄��ѳ�|C���0�|q>�;|E��(o��+� 	dU�!�$�(�B#M�|�$ bk?!y�=ޗ�Y+%�uN��:��^N��a����??��Y��۸�Ib�}��&�8���D���������>ǟ\�S$#��y��0�~���7�b����ς׆�	r������n��
�؆c��NmMo�����%�y��v��i���g��?��R9Cm?c�o�}�p��	��Du*�A4(���k#�@,���E���(�f��k��B�q�!ɝ��H&���B�����Y������2䶅���]�IS��#u�t<����'��_����ښ���Gā]���qTq5ƥ׉�EYQ}^i0f�3V����Ol�%:FR��)6C_���<�|��_Y�Ԭ��zr,�l�k��;$a@S�VΛ\�?�5X�Y����_G�{RS���OJ���N�#9<�p�^k���N�2���{r|p¤���N�w/lpi���"g��X���ط}۷}۷ߛ�'@�m��m���k	�I�׺�@�u /���ކI ��@sx� C���@ݞn� %��f�`i�/i�#㑔�Mn2(�+J�f�!��Kv �5��	��E�2����N5����]f��X�Yy5s5)��KHć='�h)׍mjil݇l���������F��n)M�"�R	�/Mv �r#�lȊ��Tk���`z]���G��Q4��Oo�2_���GH��m�u3Z�v��L�$�:&`7	�T��e���A�0HV䵙���k��W<�$M�,HE��:�qÊ��B���P u
�A5 �$� _�1�1g%J��3GE	�w�F�&G5 ޸׃LQ)�C��V�`�WάC3�h���K���O���N��`
ɢ�d ��?���Wݾ�#�  ��4�_���(M�)�q�� ��G//^� �4��	�D��u�ݔNޔ�=���H2�(�f�P���G�����������υ����s���ڬ��0��n�˽v;@��g����$6�k��CL���{I#L�%��\)��q�x�`L��j4�fzd� Q�j��c��Ā<�i��Ǔ8=D@^�,!�+F8���&8�xҏ�� ,�c�9��VA"�,'CH� $����*n�q�q�T��uL���1���#�?��^��z-	=�5���f�R�/2���,�.|�*EK'gr���V�N������YK�[�Q��Թ�N�}���7����j!/�k�kzrop_�p	O�˳)�J�:>�M.��E��81���V"������:�Z��JJ9�iL�o4^_�E�B�׹YG����Ksz}'W���a�s|�1XT��kְ'WӅ|�u%��_�M~{]3�� �'�9���$O���D�X���R����M$�����Ȳ@ś���kG�d"��n卵-���1�M������\�a{w�/��..�U�A_��B��Np��#�����\;:4���m�X���gd�G���HZ�R%,L>M����c��Aw�G��<�Cf� ���XGU�s�t�s�oO"���I��4��+V�`.x��K@y����Q/�y�V���3O�l���V���v�9��q�\�@�f�[_L��K8w/��X��'�u��2W���B�*����&+������-��c��[�+O�z���&�.�'p�z��L{����q��U�9B�W����c�'���a�\�� 0�?A�?zx_.//���B��.)ׅ���kt���o ���b���������s�$v�UA{|�7e�R[�z�����Omk�U��z
��sD��v��H^Am���#����N�ڪ�����%D���kX��q�����W\R$\O���v��sݺ��,�����{���qQ�z"��ڪrZ?�*�����N�U�t�ؑ�����U}�26+ $Ť^QeXr� Q^���q�Ex.�F�23csTL�*�^\��1	��A�έ�b&S}~�=��zBY �"��c]C�o�F�C�V�\�F�N����
�Dy�gZ�S��'7���ə<y��L�&�9&���{rvv�s��@���sV~���;��;��������"�r�+��H�ݍط}۷}۷�˶'@�m��m���kП��٪�h�&y0�Ofd�Ƨ��!$�]l� ���Rh}�����6���13,�I������@&��ͅ����r$
{4A��
��*�IZ���t���wl���G #f6�0�>Ff!�&AT8@$�d��|EcS��c�LƐ ��d��7�������*����#�S��$z@�x�0 S0H,�Ṵ�Q�٪sz� ��
$�G���F�n����A@� ?�!��	��2M��\83�^?H�E���{E�o�_@�y�k}I�I7��k&� 3 1a��|`p�>�LW�����=&o�f�?!���S��2&i����LIM�ُ)|Z ��z�/�ڀo@�-2a���+yu���G�ފ����;�-?��H�0;�D�
$�bf���:�>��H��]5G��dK����$rvzO2HHX���: �r2q �@�H���l�6�l<>0��~�h\��=2�v�-L[>mA:���_�����#0�]�̓�ެ�g,k�M���v�0���ZU�k��v���[-/��� J��Y�
TTt�z����,�զY�m���u�Zz�8P�gR�x��1����`�`,>˪)=&~���1��g/�:ֲ�2cޗ4k0R�
�ː�@-,�>�A,il�C^%�_GL��:*em�g�ŜJgdz��2���5+/xz�q��$��r�ӟc����;��/����5�U�z��N�ռ��_�������2�I6�����N``bW �#�Gi%�z�ǧr��-I�2�z-`^H0��X���yJ�>=W���}�J"	��q�'���מ�+��\\V��k��*}q��H�k|�,�-e���ړ����IMY.H.��;A@��I��j�ȅ����`Mr&�W˹ܾx.��\���w�J�a�'���}NSx\#�,��@��r〷����i����/$ͦ��Z:�U�E�Ug�K�P�<���2x�Lhl�
�0!��⫙ˆ�6����!��_9E1�A9�@q��@����U�1I��[�}O+%�8�^�[	$�B���Bi�^�}���.�D�'|��แ��VmE���1���q��k�]w|
粓Zb���v�NO��$7K#?DZ9<����C���]b	�q֛�{��Q�f�J��� R(ٷ�����v���]�y��sҒ:P��noh�+:W�G�9=�t��B�U��*�:tĸ�4	}U�UY�~C�#^��ʂ��%mE���hx��/�z�~{o˪n+vP�g"��� >�,�� }�����}6p��f�ظ	h�M;�=L� ���R�N5�hZe+��q� �#;^T�Z��r{M�è%G��?l�� ���S��shڒ ������������KiV[��r�xT!ј��V����ao�/(V�l$S>����sf��Xq����4Ya������X{�׋5���J))!��C�^�ɹ��U���GfG��|���ʟ����'�l��>Ե�3�?�ɕ.tX����O�I?�I��ʃ�y�;���o��o��o��mO��۾�۾��7��t(��Ery���n���@72��v��t < ��.4������}E���d�t�t~q������x�M�jrxL���ޱ|�y"��o�X��z1��Zx5Hӣl�:[8�w���@�%B̴��
-��Sb�0X�F4��<��CG���Ga ��3�B�!�$��go���\_]�B7rȼ��%�,Cw��$" �q@2��u��22�������
�U��F%�!�E�Į���C��%y ���:	`��I�A#�?�z:�#"�UI�2�-�Nđ�%�c� ��
 ���k@����A8�� ��
墠��{T�*��4�I(J8 Y�.5�Aޠ
�^#ȜGfmm�0.$u7� Ri�dz7'�:��ӓS�3���A� �����~[F�!�$h�C	���5�5'�Q׉e�WB�D�T/a���я#[�<Ϯ���u�I�h����v��=�7�OPX���X�̚Uhd:ojJ� ��r,��Ԏ���=8�2(y�M�k�&F��.��3�=��+#���kb/�b�E�fj3�S�V.�@���J�\�o��VVx����n4Ε ,��t��1ϓ�e�o�Bz���}���8�����&�Cf���YeL��~.`Na�z���& �(R*�$e?@�<��U����R�Mj ���(;ˏ�U�uD�Y��JX����Zrs��W/`B,zD�
D���T���H*f��x�=��ѣs(g \�*����B�P�I�@�~~-�ru�H��f��@?N7�%�%��zR+�tl*3�s>�ż���\c���,�Z����I*#K��ryY�R�	�� Q�=�F)�U�}˛y��3Yf�%�dr��H��I,���!q�K@8�(��}TJ�y`���1������]�W���|c�w��^!�<+��͍2��el��,�y��̍��L&=���~ �Y-e����k=�Q*��r2rFƨ@u_�s] ��90�F�[�75�����s�0�bil"9e��`6������@��c%��	!�I�n� �M�^AC���K�yY-�ons:aDU���x���Ӫ%N�z�Z�_�b���!V���X�@`����$	�#٠�X%)b���[�-.����<�,�k��d��iҒ9�ؕ��a�*mu<{���'���^&�*�L��@�^�7u���y�s��뒄_?�p]��Iw}c)���?�o�� �ǵyQU��]_j��Xk�,��e�#�kd��δc 6�Z96*'�X�k�[aK�0fG�;�fg'+|����R��y����dyM��2o8�dXH4Q�3a��:1��m��_��$m�����
>;�K�(��Y�)}GՒ�΃f�
x�9�#��k� ���0x6�z���$��u���D-想�h��V��}>>��#M��q�m�� � �g��r��(3X7�V�{v3�8�$(�!��XY.ϥ������==K1R�lS�����v|�=O�#�\�H�繳����,����{?�}�?������2�ȑ��稁s��G�c��?�Ƹ�Ⱦ�۾��N� ��o��o����!;�6�p_��i�	�P�0��@ґ�h �J7y�n
!Q�Z&���T⯞�ٽ3��9>�HW��X7���;y��n&��Τ�F� Y��.�ďmC�,Hה57�8���ˍ#7�.%R��D��	����+�����2���/���βgY��^-	L70��{���`���A�l�G���jH),��(	N!K��h7�) ��B�yƬ=Tz`[����6������fkV�\&r༖�l�c#�wH����Ì^7�K�N��'���J J�n�YQB������k��J#@�,d�@Bªט���4!������LJ�Zn�_W&��ɏV��� �R��\��0�h3l!��ͭ�of�g���o�ӧOy_��.Ht����
�M,����k���>�XG?���#z��7[/9 � A<T�l�A�MB��^;����`H�qQ�Q�{P~�Z���r��ﱪ���<9bUy���=�Y�bsȁ��;�ut\{�
��9����	�an[��V��4 �W��,�I�J�y����W��A��iy�-� E��H�.�Ꮕ�|���f�k�7 ��ߙW�� � �t.C�<��Ka} ,�Y�:&q�`�^B0��(O%���UT��jÔ<�D���GN"Y�L������5���;"���ru���V�����ܗ��%Dj�/��&&��:s����l*ӛW"�gd��f��4�}/Q�)�=k(�Ǣ�s*����1��P�)͟f�����m.ח�N��̴��Ab��#��W&3�� >�����jy-�<�W� �*#jq�[��׿�_~�S)�V���B]3�9Ծ��]S;R#���yv�h��A.˵0V��	 �[Y�f��s�y��;����
D�\z=]�c��o�+�KT$Z�z�M�6��n+ޯ~TIW�	�̠ym��1��#�V�*G"�b(`���?���?$�\����e냰��C�	Ǻ�+���F$��9A�\oR��Ց�`H��R��qԂ�4�rr����˝c��s!m	Z �~]dLi#<��;_}L��MM�)���ʌ~Q�yGx��k��I��,�}��
��@���;ä%u[�1%�*�<	`���*������UgF�wz���Q/U�c���5���uf� ��BY�� :� b�>X��y���=��y��V�9_
w���yd`Q�$x=�+��	�v+��;M��K�<w�H��/I�g��p��N<��e]9���rM��0��3ɍ�bVW��(5Y�����|P�0�Z��֣-��̵��qA���Q�@%�*��an2X[�C�ꌶ�����0l�1��_z�,T��Ո@���a���L9o�܉������L�߻�$!�g�9^urr$G'�<���=�pͅƺ�r!w��������9�,��ՠ���#�[�@�MF#�����\�5��ĝ	�d&�@��ޕ}�˛o�-}���������LuQ:Iֈ�����2��T�$�5B����#��w�H~�_ʾ�۾�۾��=�o��o��o�h�ǩ��#{+э.��!��Z1�v�θY�hd]���o����Cfw���|=tgO ���_�K���=�)1q7cfj��抙o ڡi\��Pǅ�QM0�d2��L�L��J V��6�'rxx�l����C�����n�pC�,��/�s���/��Ͽ��/����W���s�\*;�}�wht~w{'�%̆@)uӗC���x�������F����$�e��qL�QD���L�$�Ѩ�����}Тh�w��N�G��3��RdӰ�"f������\~F���'9� wdP6�эl^;Y+�#���kf�^:��LI��{f��ex234$(��`v�a���dAv��>����5eA�W�d�3�N�$0��T��L֊��Ġb����O����@�jS.)��݄Έ;�f��7 ʨ�����Zm�$�<��A$� +�LU=�ָ����Pt���U成-��%��>f��u����2��rF��U<���/4��^�s���]8�^�b�~TE���@�4�402�_���q?sjӇ��Ό9�n��1�9����$0(?��m<h����&^n�~�OBg�\�U,i� �BJ��YXm�,F6�	�dpld���Kʇ�"�$�w�m�I�Av	�,6	�f�0�5��<���pnU �y���k�O�r���r3��!���"�c�B��
>���1�w<�8����ޓ�2�X��Lo�ɸ����YA �|��v%�u���"q�	@�ch
Z�J1s�}�t�;uJ���j�sL���X1B��jl��p���#�.��,�����v��z�4��Y߽����k��ʋ/?�ͺ���+�^����z��x!����t�Xil�)F��>�aG��a�~+��P�2�	 ; �S�ӣd<�X����eisDlD]�gaZ�[��Gz�q.�~ld���kA�K扞����g�=�uQ�qkV�tpu-��ex0��r{}�cp-���pr�ߑ���1ވ��V�WV�9�$V��&
۹K2�ι�td��orqe[H�ڪ������<o}w�|*��f��c��֫�dh�2�C#�}5��"�
_I�s�>BACY9T�!r<���A_�� �Э�?p�`�̹'���!�"��'�7�	"����İ�1�<iS��D��� ��F�x�/���k�Ѯ<��F,�IE���c�{�������Uux��>�I͌�{Oٺ��n�W�Ǐ]'Z����n㳿�~���i��B����!��%� 5���D	<����Xp��9�7I�lZ�,T4������մ�����^'%��s�k-d�H��ma�*{���^9Yа5&��IH9?)]�F��ޟ]}��^[�9[��i��+��*���W���ڱ�J���L�9��~p�<{�T>x  ��<�g^<���g���ϗ:F��[9?)���|������Y��R�K�ҕ=o���+��5`<H��rb<Ig�5�����ٸ\��x��!����ҕ7�~���z�}��������D���;xF(�]����A��_��/~���C��۾�۾�A�=�o��o��o�X�3+rf���y@y�u���R�_���₾���f�?�3��w?�t�`4��C���_���W�/�B7:���|&�n��Z�s� ��92ICK��
ir<��2���wz&�����n��R���̲4���&( #n��%�7+�6����Hƣn����f8Ol$��o��O����7������G�����f:���8���Z�	'��M��X�\Vh��D��SY1��Ր��D�����J����+3g�66�����-���3b��g"���F!���eܬ�p�#�XN˝z�E�uF�i�p�&ׁ3�L�^��FQ�l�2�S�r.'6B�,�[���Oa�E�h�� ?�ͶU��fFMCXT�x��g4��dxy�еq��4(���x@��%*j��5*^�WK�<�l	���e
����aP�q�U�П4ؠ�$h��w�� ^.�W\xR��_�u�x���Ȁ,d��uo�楩hfY�@!_E�s�̈́6Y�-��1�|OZ?_�����������v9�d��+�4�}f��([���[\J)�%d���q\?N�?���u~�I���+=�*%�i`��K��E��h���ET;��7�ƭH+���'���m1!�d�S2ҘS&:�����k���o�sו�K�~~	{	y����Zw$�y@������1�Ôq�H��_^H]\���3il1Q�Q���$�q:�,���l�ӏ!�@�4���A�C~chS����D<y[&}�3��O��.��z=�7�,�L�"�B�p@_�����-��~%/�A$���M/4�W�0�w$���ȓ�CJ[��A���v&s�zTu@��3��?4�S	�J�=K�Cۥ�xa��rY:7����L4��Գ�Z�־\N�G�԰$'�ǒ�H�������S��S�7��z�#��$i%z���T���R��U�*�L������%<xH���e�/s�#���(|�)�5 �U�u^Q �s1b�ұ9��By(ąMi24����x��/����iH�l����[�����㏟o~��w�U�A�������_A��t���36Ǔ���s�=_�f�wU[)ƪ>��^G�
 G��@ލ[F�[i=�+�T9B�W���;�1�VHxi0#V�x�2����/ʲ���O}���V9>�y^�5�'	����3�n^Y�)�>x~��R}$���We�������??���A@ 1 zY���&�'��='dȞ(KW�5�A���M��a2�f@NB��XM{�\g���p�Q_hR�f�n���Z4��X��[�>#Y���
R�����?�H�k� ��0����ʭ��ר�Z��t�e�B*��)F����G���<y�D�={&��G\��Y�1[�F�9dg72��F�̨t�;��1a=]h`~���g�~$�|�J�~�ϯX3n�����Uq�ޗ�˪�Fc���Ŗ�����uk8�E	�F[� !�1�LX���{����'r����@T�o׺?�>����m}�].dzwg��6��sW�LP���R������/��_˾�۾�۾�a�=�o��o��o�X;<<��_I�;�)06��G�������������D�?!�閒�'�t#�ɷ?����O>j�G{�.rT�){���}�_����������F���rzz&o������cI �n��k݄1yp��D;�_>�����o�fꐴ*��U84��$u9�ݬN�xu])|A�*5�RZ�*�.���T>|�����~O7g�*���ɯ?��l�3V����.�eЅ���$]�h��;����n�ˊ�l���F�����d���l�jf��*��|���C}�Ͽ���־���'ذ�p2�1^;??g&�h<�9�����ΩgY��lA�Y�k�0@f.�p�����A����� ��¨\	:=^�_T���Θ���������;��^h�}}ڣ�(�J��˞�LC��z���̜0�J_�@�z5��Q*ϞޗÉ��2��l�s�T�:�����}3d�?��H��C�uHOLh"�c�w4	�����.Y�Ad� �PR9sJ��M�!O`�6Ȍf��#j`FJ��1D>sUP �p/p<�w���R�����Hh13�Qb�G҂�x��{T~@O�y�s��-��S�A@�e���L�0uf�13?a�j2:��,M�� �������ev,��zμ=���C�?��}u�U�$$s�ǉ��������%b����!!PՑ��^3�@X�f@�H׼�R�$�F�NVJ��Ҥ[jGD+�a�h��s6�J�M�Pv��ӹv9�Cd5帿�����B ��ȀHC��B�>����rY\�)1��,��$֘�(%_݉�J���_���%<y�H]��?d�\E�μ����� 4#�Ҍ�Q=E�rR�uI4��5}��3y��}IG @�������d�X���Zt
J�E��I���?�P��H��@��.���v-��<C�N����5?���x:?�e-�L�ו�.�;Q�����X�ͭ�&'$�P$|�֙��L��|J^+'{��bW�JP�2�Y��6-���+�r0~
]��W��>�N?��ޏgo�r٬r�ZGzO�R�x���/_�r�RX2���H��}r\�*��t1�<����*ApȚ���t
�t>�4�Gq鱘e߷�9���=5�&��> �uNVҴ�g�*��촹	� ̉����?�GXӻ�2*��E��[�3�hW������!Ɛ�pUY�Q�U6V	�~֑�^�H�%MQ^��C<�r8>�;���x>@���l�A����2��YoV�/c�e�H隇��e�ZB�U���*߼<#�+�K�֔ r﾿�k"��k�c���:��rY�8?����W6~�s�y�4m����O 'Py���$"�˒$:�y,qL��!>ZEP��$}�i@ٱ��7y�dB5,d3��>C�[82���>g�6�Ʌ!�ԕU�����fc��T���Ȯ2��<��,��[�MvCT��%*p�ʞ/v�8�Ȫ��<}T�v�����^)�NkGz����X=��$%�T�I��s{�h+?�'�S�r�����G�����6�1H=���Zc��**je����������Y�8�O��>x,cN������8��_��j>չ����k���q��u��}~���O3y���8~5؏�R�������_��_˷��]�O��#�����~�k=ƅ�t�<�9�����ū�Oȗ��*uU�����^^��?���m��m�����	�}۷}۷}�F$!Jh��[;�P7go���|��Z�?�X.ί	 <z�T��?��o"GG'ܸb��e��	x�3M��3+�sݐ}M��n�#�?�.uc��_�SIcd�x�����G������flt)w�W�� ��χ�ځ}�¦�sI�� �Ii������f�kY#;�@ 4��]y��Mn���>��O�Y������W?�+=O�''���1%2TM+�����$(#��?
IHFljYW2_����SX`J0�$�1�k����f���#��H7-���t&7�7<�>��A�0Z-�3|-�p�L�@ w�iZ�<�&8u�?���Т.m#�`�O��^��"3o�ײ,bƳe���:��G�׹D5�zA����	���)�� @ @J��y욺�:
ˠM�5x���c��Z h�/��P t&/��֟Vy��V�9Pޤk��YoM��\�29�@��:N��V��#+W2"hlʊ�mU�o����Z� ���������<�X����i{|/���za�V�x`�g �-DS�	�}��{��ؙ��O�ުZ��+
�΄�g�{�qY�^��_��`��?��#��!�?#��pi7��~\k\61��/bR�8Ckj�4+�-�� ��Z����C��Lv�*e6��N�������K���h�(kYܬ���S��0��ԍ��TS��QA�t����2�>�dS�+�댙�0=ǜ�Hp�#5�&�,-a
0 ���4	�l_�Ю�B�� :Uz����d��d~SQ��;�3�ߗa3d�IE_����LPus���V4Er|2���c��H֐��Z��s=��z��Xc���\�z��j#��m��i��lƙ��FC�*��(�X�wk��1��CaOca���J�=��+'7�W�jWj3�/7ff>U��5v��ƱuN�+W��U���d��v��o��:�zM��ɲ���8}=_ɀ�c2{>[9����CJ�(�<�L�t#��<GBW*���0h�	a����ƣ��K�����@��ɢ%@v��L^N�{iR~�u ��h_���a�l	&/�G��w6�3*t��plMH��\d���d�|�IS�QE�3��_U�e�W	��Dm\�m���׸[R:2x��Tw�̡�-�&����R�K�"���ҵd��t�`���ޟ�?K��՚�[|w�W����h���$���@z�_���7$9�k<�[���2X���$�KJq	���_�İ5���qN��E����ja���82�$<Ӵv}�}����7�U����ھ7���EY'����}�����թZ�����2a�d�e��d��t�,=5�ey�n�2u�Z�JT5˓���t�ϑ�����|V�_!;3���^����N;���������g��P�x�]y���=����O�'��O��z������Tj�O�É�?&a�)Tf<8����"/��2��\e,��N�w����Ǐ�Jo�7�H=Õ~�󯿒��?�ǿ���z�0tG���Y��v&���st? i�l���s�u ��+�7%��o��o�����Ⱦ�۾�۾}����T7G�YEfף'(�C����,χT2����|��>����2��e������gN�wH�F� ��K�����}1����k� ���>ɋ�t�2�6U��dad���G������8s��sVyp#Z5���`��9p��;��H7�L����C"1M�׺��p��&�'�8��{�����G�l������U��n�{�; l� �PCZ�S�hZ7��*&�"@C�GL�5�W/}�FC�># zi�l= #�����_i�|}��TA�s��u�H�4�IѬ�e����" o-뿡$	�&O~�T���$���e�
�P��9Mk��M�Ҵ�� ��>� *���*J��T�pF0�^�r�d���(6��G+�?��/I(�J=�o�6[�, �@Z��]���_)=:�b��I��d�����-J�� W��*��@����໿��T����rW^��P�|�@��5�Xk�%/ی�����Q�����V�sG6��ƈ�Б$��E����tI ����f{��H��!:�Cb�� /�~�^厰���h�@��AF2y��S�Q𺱼�b��V�q���.�M`D*�t�J�bʥ����?�-�1��RuƏ�1������sU�@���l} ��EN��_�'=y��D:=ȳ��Z���y���K�:>x�P���d$�
	�tƉ��qs��Pc(d�b*�yE���и\o�0%
���'���.�]G��OJ��Կw�rP��0(u��wC�1�q(�CE��V8��Gڟ�̲�`]�>*d�Y%�(���R�#gf�X�Iu��$^Ur�j-��]7��Ct�X��D�{u�����[�*��r)��J��Rǧ����]3�����L��Jc��$IW�X����յ��HJO��#I����4�+���$<jT,HE�1�|@���׭�x]ф��Y,5~��W��P"]�u��J�)�o2'���`1�g�.���.�f�2%h�q_V�IX��]
]eO�%����c�W��>�
�TnA�BU(X�RWR&/6mE	�э��U�X�V�<,�J&�3�=f 1��~���.^�mƵ�K9��4���\?"'��1J����@��zi@#W��1�;�{�n���{�=��M�}5*�	=m�hF�_�hbm
c{�lھ�w�l���J{���Oֱ�H<���@���:"K��,��k�D��ɣ�Y�P
r[���"^1�$��^G4�O8�BVU|� ��4)��o6����u�	-�"�Q�."���Dv���0(��Y�%,�k����9�5x{!�GQ��o�k1Bd���5٫�UY�:B=�^!x�й�'����<�i��^ż�+j�,���S>ˢ:�w����$LW�y�u�T�%غ�e������K��d�ըR���7�g�y㍷�ܮ�Y~�����g3���IN�u^��=�����EH�Ae�z��sX7q�M�,��������?ߠ���l��7���/�����_�����o?AV+MB���X2��n w�k��zm�*L�m��m�����	�}۷}۷}�O��x=x����T�WI�^��Y]��x�w��|G�.��w�������l����#I�����n��?<�}�gr���܈a���g#Y��~C����Xp `� 2-��%�ؘA�rG �ys$p<h�M5�;v���U"膷��AH� `���R7N�����Ʊ@� K��?�Kz�Lo��O?�s�8�nll̈́y�jxC�*��;��;���p�'P���;4�Z���4��#
}p��V��
C�>���	(d�&���d�����g�G�iL��^��1Y��� !�~h��gpzẩ#_E���A�⣢9���Bc615�����O%�0�U��K�?�(�F|>�(��� ��#��1�� ���6 ��x<�k�����x�)uSJA-]�0�' 8���Q�M{U%u֭BY�^;�g6�y��u@:�>��!-b ��P�Y�t�@����"���ތ|ל�k� ���� ������ַ�:��c�mFΌ̓��0�����î� �j��F�lZtG������I�P�%�[y�+�D�/�=^��g�X�r��qU"�xm?�ȷ�
�?�-bWy�k�G���A�k��{KE7���\�I ���",?H���_Ϧ�l��r���ǰߓ��PFGGv`�>��s��f�
3����Fօ��t.\U����4|R�KO�3<����t=��kl88��p ��޻խ����'� �kPй��j�Y��"�^\��b�\�j���!�44����� ���)�G7�Ȫڑ��y�`~�C��G�1��|*��k�O(]�R\DO��h!cY�p�*�$�:�`<�����|5�7$3V�R�ӍLt5�y�i�����zO��Z�~��T�|'��٪��_���V�s4��K��e*7z���K����Pz������)wЭ��t�[erq��"�$Xٿ5�F��k���zD��W�p�9�<���b�����YΓ�|#x�2����Q�d�@�8�K�u�+�lL&�a��u�?�]|�@��0���!���������=Gx�u�����II&��}��0onZ��ʞ�9�+2��C:Ջ�ǐ#S�w�'�!f�gǁ��k���ה� �Q�i�����f󹓀����=�
�,��VmGN'��;x�]刏O�;��1�ذ��:��]R?��˒y9B^W�:��O�tBn����^/�k�O0 ��c'+z@��
��	�CJ4r�X�˅>/�K��Mllᙥ�9�$A*_"�7HLC[�3�"��$��%N4M� I��P]��� �Cxv苑kv�v���&�1��?]�Xo+?�͉Rr>�v�v�;�*?��[�����`�G�xr >�����޽{�,��r� Adk~����y?+��*�Y�b�m"=�U�؁8b���Ҟ_�����`,�?�����±���y��^O�����R�4b���)�us3����Pa|z|"O?�3<�@}6�0�&��?�T�����O�Y^|��+��B�'��jJx�0�������k������?�󿐟��gI(��o��o�����Ⱦ�۾�۾}�����=�0=���No��y�T�x2��96K&�����˫W��p�!��r*W7O�7��|�]��ѧ�t����	�x4�G9u���]���;o���SB�0��5 ��VM np���4@'h�t ��I�(m�-� �.�<��(,�EZ�a�j��.�|����_~)r~~!ÁG������p 6�k�{�@FNn�2a+U�T������4!�ԁ@I��yD� �'�D�D�B~�T�/������8��e��2#M�<0��A��l3!ӎU~����	� ��Y�N7�'b@�сS �@j ���oc����T4� �7��ٵd�1>�hlខ�A�D��?��8혗��',C֤�P��|(v������U���L(`�*��/Z���x��2/Z�6�>�S���U�J7y9�]#_O�x ���k�~��q0?�'�y0��+�� 0�y�#�kO
0c'���N@y��2��q�	
#_J��$7|5�ɍA�$�H�m}����*�Z�����V�HO|'*�@f�����w:Ns/w�����<	����V����l���^�m��(uܦ�I_��rt|6��̮?�[v�2{'1��C�ZB; �Vk�f+�ݮ�#������!�2���Rz�X��\� ��k,��{W���_��ý���Q�T�����t�똝�Y��k���Wzn���N�����9�X��*V��q�A�i�A�}ҝH�L��{z}k�H���R����T�cs��:��T`0��_j�|x-�u����ר���W�i �X�:Ws�����ra^���s*t\��0[�`x��S�P�ls(}�Y�~D4�-s��Z��"7�"��UP��`���a�����l�I/X@��Qǐ�xӀ83_�Uf���8�:�����<�Qmf�y�Ɓ��4�B08�X�Ǌ��2�q?�Qh��&��LR���:�,�b�A�J8Σ�d�P�W�U�����p�w�+|���s�����Z�G���u��4��q<	[	+F�jW�)�ߗ���CzW���PaRr^&������."3�3�� �-�bm1Cy/�T�ﵵ�v�8���i���+K�ԑVrkP�����fX%�'p}���UD��J��1��_��>L��
��c������w�'̓0��`����')�ĕ׹_[[p��>O�P�Б%���u��#V�5x�)��Xҧê�:|���J9��2�}}�Uy ?B�t�6V�W���Q�A�*����,M��d�l��N���P��誛�x�:����wC�Ҫ1�otbG_�����R�*o���] ?RG*��~�b�$Ҏ?�+�7���3y��7���_3��a�a��󆮧 ���sg�3��<���X��!VӃ�V �����qV�M�5c���������T2<��7wޓ�>[��������\A���s�W���$�\���Bc�󯾦VN��.<�9!uŊ$�>װ���Մ���^Ϟi~���ˏ��o�8ݷ}۷}۷��'@�m��m���?E�裏Lށ� ����jd��M���9����N߻�O�Avo��#�"��Wܴ3�4 �B=��LKVE<������{��� -��g���p2�f`�����@�� s�Y�У�	��u��?Qd^ U6��wS�`Q+�����F�����PK��K9�ȣGO�?��|��'2���Z�K�8r�@(+``��>s��E�|�@G���M�Bq��L�(r�!3)���R�I\���8� ���.!ce&��n�����HQ�g�⼰�dP��f���ZAٹ����J?�l{d�V�b��N}d�M����`@��`U�ᰭ��i��sCL�� ��2���a��D�w�4�|�,jd�cSo �j�izf�#��W�@���r�zS�K�p���<���%��,����H?���ij ��4o%S|e�����Xޛ�������v�jw��}U����ｿ�?A����k��$
*��h�%�|�|~��VBnxE���}ss�z�x��<��׃~֗e{>k�g���bc�>��$�'[<I��K��z|x������@��
3�������g;�0�d���q�l�2*	�a|b.S�I�auٽ�Vud�' �~��S���3ߕ��5@I���D�3���!ݝX��Fw�:��Fr��
@�:���_G�2n�sY7��{�����7���+�~66�-��������N�j%�����Y͑8BˤWP��D4��d��i�8~M�\��1�;����`%�M_V�!� ڀ�B��;[M��W�����÷�a0ֹ��[��f���ru��������n�RʨDA.��:z���4#��ܸ7+�,YՀ����cf��"[��Td�t�,%��T�AGz��a�&U��������ڲ�[���Q�C�s	��7�k\$���+�_����0�aWש�d�(?��ӈ�a�U�yr�_ޘ,��0JGf�%$�me��\���G�˸���XF�u�)hm�-���]l4�m�1}Օ����;y$��!���8���=0o�Aw�b���l�ϘD�B�RQ�jd|��^P�r^x}���1�ǭ��~�`m�*�D0�sC<	�cL��X�s�&�Y�1�$��d�'v=Oh��޴�}��w���Kn9o/��5 /v�BȘ�� �K�C�+N|��?��;^20���}������:���E%M]���0�]E�]'}E����OW���y`�l!	g���p>$P�9cҒF��K~H
O Fey��I����+�5ɏ�h���Iu�lEQ�s����U �P��4��~p|zV�YVn.�{H�DV}zO�o�<}�jf4<� y��z]���eՎMȖb]��Qqs�qF�B�����2���|~L�$��X�ks3`e�d8����-����WϿ�/��T6��'9K�����'�5����W�*�`R�|1���;&'����Ʈ�������[��;���`R���$�Iv \5�e��D;�~��U�����/�B�m��m�����	�}۷}۷}���G����?���q3��j]X�&_��5>#�� qX����~��׍u��gUD��rq}#�7��\�t#xĬ0�����r6��䀾�8эUWziWF���ѐ ���T���d�X8�BGrU.{��^>�F�z�c��9��<GY�,�4�n@x���z��M��kY�n���ӧ�����_|�)ϩn���V��Y-%�����C�;t�5�#V�T�HѾ�M���0`Z���&T�! mk��ȷ�M�Q�U;�,p`BE"ě�Q��|��，*=��B�� ����u�*ʆ8�O�(A�D�S'hAy+3��z��bv ���e�:sU����|@��>B[�nz�x�W8i���䉆&�J�@|@ T�t��
��+��Zƣ�,���n겆fU�, ����ͷ�Bc�I� ��&0�m�LX��d��k�Q�
Y� 4(�fਁt�ekR��Bl �,+<������� ��X7�-��KҘ��e='q���N��H�t}�}�~(�
���W�$jrw��#>� ��w���� 
r渾����g�z�(]W��HT�xRtD+��T-���km��kj���:0SW�3���G�vÊ����^ߍRF�����Ϋ�4$q鯒�g��Q�1��g�� H��Er�S�S	V�&���F�۪���O�cY��M�KH~-('�	Q�Ve�/�*�֍^�\cl=�����.�G���H�Ъ=HU�D�U\�~O�R����C"	֬t	�;�#��HϹ/0˅�I����"�y�qez�\�����1H�~���lQ�J����� �+��o��(g��5���b%7_�B�f-Q���$�nRJ�]I��1���!?��U(���J�\�:!�:ꯙ�������a�9I�~7�n��[\�;mzD�w���:�{�E�9 ��#�!j�fh����+�	�~���L�l2�S�#	�p��h��zZ�^[����zͨ�'��1�C�b��gRN89$/d�Y4Qn�RX���޻�r��5�S���V�
>H|.]�瀪)_� �W�$��E�Ib��<)���|İ��j�+ĸ'턪F��7L�����f$��Uݴ�����������#[2���a�=/�씏�F���O���%ZI�p�u��M+�Tw|j�0ck�oO����|sU~��)&$�;@��(i�+O��{=��'�����#IL���}�U����C�ȏ�h�ѣ�l�研�g[�1[󑈲�s
^�3S�-�a������q��1��ǧgώ��r������4�φ>=�٘ٞG��Jv�<)ǉՠv7���Ge|���	\�,Ͳ�������`,o>y"O�<�l,�%Kw��˕dy֮i��t�����&_i$����pꠊ�4��(��1��'���}~u)'Gy�[o��/H��իdn1�I&��OO�r���ӹ�!E:����_ʗ_}.��|F�/�zMϞ��
5x������W�!Յl@D���NB?I��Oc*�P&��}۷}۷}��n{d��m��m߾���G��Y��>� ��d,�?0_	 8Gg�`�r�HR#n�z��������W܌��?ۘ�*(K��|S8��u���^T�tswqq.w�w��O(���A>P� ��=6�>�5a���Y��r�N�I)OE�,lC�\.X)����ol�A�����	�����\���ۛ[�\.d�Z��<���Dϩj���͗WNZȲ�-�1"@�T1�;�b�O�1A �|B�?QXdJu�Y5Js�~tRb��<j�+|��U�5�t�s���U��!�c#׍�'2;Q郍uc��,k���3��F� ��zM�C-�0�7�dB�F�|�d�7���.Z����}B�a@4[��,;@�@�F�� ���,�U>�0���,�Y����@A��h:���~����dL(���J����fL�V�� ��2�����8��gS�?w3x��o�b��������B(�J�-�O0��,����͈锷�F�F�D!+��� A3�j
��ش٪8/ka���c������ӈ1ăof��q�+F>�pΪ�ͺ����<�� ڦ�������g�^���[�`��t����	�S�]x0 �Df9��X���u�[��M� b�O��2���y�0���-(�R����u�Next)��T�^{J� K�;�e1D�k/X��EJ����N��&��`U/�8w"��M金g2�$��$nzIGn�2�L�tLo��	o�^�"�n
n�&��9�>
��p�~�F�z�!\����@5UŸ��C���s&.3�{���^}-=�k����z��łU\� Ҿ�}��P�x-_~q+7Wzy3�{�J׋L��;���|�鯴�n%�<|:��I_�i%q��J��ʑ���b*�~׭��v�r�Kw�Ǥw��/�� �K�x �Rz�@��T�o����F� �C�Ot=�s�Z3��$U<�ӧG��L��i��AmZ��������������"V�IW����
	�ÕşƊ��:3^ �������+�I���@��ǘ"�B[:ʗ�z�x�!T���t�H��P�zZ�-�%7�
�l���(��^�5q�󏠾�[9(A.���Ǽ�e���L�-&c=A�%Ⱥ�����VV���uh�������[����H�V� a��8 ٚ��D���IZ�%��F���U��U�ȶz�W���s01@�6�z��9$c��E� |ic-�lQ9���HGxx���-F2�/�<� �r�|dI-]���X3#�h�c	+x&h�M�<�d�r�b|����!#��З�Ѭ��`�����?j��^���B��">'a}�5_�;H�Ē"6n-��Ύ�\���<��a���8�	�a�g�Э�g��L<�*�^���쭶��x$@�'���#9��k��L��J�-�3pQ٘�8_��l�z����:8��aT����!����F�ij���{�wU"Ϙ����W��;:<���=�����>���R�zZ�y'�9�XBk<�@���$�х���J���y���z�������7����t������}yu�R֫�>O-x�P����y�c4�x0�Z�[g��+����ʾ�۾�۾���=�o��o��o�h��ծ��y(��[��ld&
T[@s_7c��?&p�����2[3o:-h���V�ȉ!K���fJ:\ a.>��5���㾜=z G�����be���Ɉ������� ���L7q�f��7���bS	 ٬�H��!#��*���H/�6����빌usy��Įn���x!�NOY����'���ǿ��|��_Ƞӓ���R��C����M�nt׹D��ƪJ������)�Ċ	�?2�L\!�,��;)uS�!����@�H��X�d��S> +sV�PZB?����'��jS��X��3@7��N=  ��z�~w����C�L�;��э����*Wp�] 6�jJ- �o��$�:N��QJ�^G蟔��b�B!�[�ش���X�ev'���L��,S�ApL�,/)/B��!����z���^�G��X��@E �a,Q+�)v���/�!�;�"J4E���B��4�
> I/�~�$� �x��\�+V� 84٥��y��ڝJ�� ���6���[�0 ��@mMˣ����8<\��[̬�j�2|7*:z����4�H�xec�9�Gc�`ؔ�_�x��*�IA[5X�;��i��G3�������V�8���e���R��5!2ē�I����7��ϲ�Lu +���H���@�t��ȌX��B??� �:�8��vPq��
Kư|������p��Z�.�}�ڪpm���,K	��H�H��}�ŅԝPr�'��S����%j��
0s}��Ij�Q�]\�o�ɶ��������h �@�^�J�/��L�qp/�I� ���L��E#���R�aA	�4�A���迁�xPR���<TO��4�F%`���d���Z���b�s*��X�����
����ߓ��-�ru��Nl��{c9h�[�>���xp��H�oa�9'��5��B�u�!Q�z3%���ǿеc*S����<:h��Q�,�r{ug�ȣ��3�%����ڧ����7�[�=9���1�K��ԐTo���A����'�%mH�7��Ay�J:�T��*Y��60����%7�0^���1�SB��n:��릑����`F��Q��g��G�%*bD�~�
��䚕@,��"���:��(u�:W�x�g2Ne6�%��2�Ѥ�@�#>.f��0r;
"'g��y��P�,}Ɣ~�?��+��1�	�Gޓ�����0g����d���[lK��<���yoXEd6���8�2&ayh`�	��a�l�wIBu7 ?�>1Nfs�ok#?*#K#�aV����&T�,>!<Vz�X{����2}�@��h0r~)�PܒF��3vw�m�"bVĈDZ@�j�.�������̬Mz���ױ����G�h�uR{&C������~�,�IL�*�$'�RBcim&�3�?$�@��O3�Ј�Nj2OHl����+���c��@C��>��|.�=��Q������^@qj���ʡl�XeR�ʗ��X+
HC���.�������{���lc���5~C���]cI
!��.X�W����7�h��g��̀���+xÉIa!�:�2'%�.��S�Ƀ���Xb��3��k�
<g|��sL���o�`� �B�5�9Y7�g�T4�8�{�
e�gH��hclf(�zz���9zLH���9:�9|�@��G,_�qwyMO>��IO՚D8*WG�ν��4΃A����~��ɨP~���H���Ecϓ��4��ȷ���>_�)��V���[�z��áMXe^���+����o���dU��̳o��o��o��mO��۾�۾��7�"G���(&����e�c�l��e�a�pr�����>��~�����&��w���R7kG�Grtz�ٝk'�D��B&
Y�����> u�$$�N�A S��5��6TؔB��p����>VO��6�Cu���u�x�����6� ݔÌ��ݱ�l�IR]��2ӍeN ���P��������gK^.���IM'd�ij^Ȩ,+zX`�O�gHd�y%T&婧�0�-2%�(uY�E�;.�%�I��@��%+K ��r#����� �\E�e�5�0��u���f�C�Ǚ��ܘ"1K9��N���ޛ6�qeW��w��#7$ w�,V�Ԫ�U����ll���d�S=K�%Y,�I@�-v��u�9�yd���|��*�� 32���[��s�98O�|������d��~�h5K*��|��i����,h3)X}i��5�( Lb��A����^=F�ͼ�]�m;[\?P\�`�B#6PM�l4�t��ڃvS%,�v�,S�߫:;K��ҷ�V6����2�;�.k��!{h����y�#��!ޟ�>-�|�*�~���<�#D��>:_���H��c���Y宻��2R�e�濥�[�����
i�a�%.k�AG�{{N�bׅ��B"�1Y��س�s�y4�=t����i�X���5R�:�8��0Vt�Ce0&�|����l}p/���U�����o� j��fk�;��::��*
��s�7����<�oЅEH_n��b�����+y4���f!�f&�n���}K��E�h�Ff��7�lgF�RG:'n�wr;{.+�c�K�Ҏ��0�hK0�qT-�f��fa0��M*p�ˈ�J�aPد�" 9@�+*P�;`�9	X�@�;�-4���a�R�_ą�/�p�7Fn�
)w��o�^�t8`&Sr��%�G2=�Ye}s�׾�vx��sVY�t!��4c�:��V��Fm/�mN��b�sw_o�(m�?\ɋ��$�����z<Su������
���2���n��?�%���I,�!� @�u}��ɉ�raj���J��JRYI����2��Nj$F����ƫtLV�X��|���]�λ�G�5!�y���Ź��>�֜�I��D0������i���S	�^'	��k�A�<kyP�>�	���2�6_tJ�@����
#hEW�u��<���} �'�H�I���Ij��ء�8�y�Jv�.xN��]W��m��[������]��I`v\�tJ�f�@Ltvz�;A8���iI�T����v*<W����a��"���/k0p~�.��©��g�Ud�
�h��N':��2wd��X�j�*�>��\�5b���o�����p�����`$���`h�:��KR����27���~�0Pf#~��P������gye]�yIEk��qJct:�3hZ^/�E,TE��J����sq�o/냩S(&$�:���MٝU�4�}�����	.&�#:�S�ix߻�Nw�����3��	m����<�ty^�N�ȄI��G<o��E��
Sm�����Jb�{��xA�P���΃��,u��;�2�,��{��e!Ul���X.?���/t-Ă�+�LPhǑ=�M����ͤZ�y�ռ��?D�n�>~��FC�iĽj������t��ӹ�;ƭ)[��?@�,�.__ȏ�q8���3;��8��p�����~�w���7N�a�WWA�j��p�pD������"�%�/?��<�7�����e���d0��G���'��O~�K&���-��uA{��$c�/�U���i�v!���t0H�k�55Ce� V��-�-�Y4P�d0mS�{?m�(��F����6)��l�!0 ����r�$ k�X?���&���X�wt4��>�H������Uw!C*Cؐ�Ii-ۦ��� эk�^��0m:BZJH�r#=��P\���"8@��k��#7�q�!���Ξ�Eހ�x�$,@�x���.�m\դgj�
 ���0k (;h�����@���rg�ё���8��ڪ�W�P2��!`�W�|�MYDda���|t�֝� A����8oo+Bk�Ƚ��� <u�Q��GL�xO�4�o݀�HU�>��Y�l;�����{�o�U��>��˵�,Q�{�}E{�������8{-�<�U�ā�S��a譽W�M!X���e҄{b��̇>vvS��Wg��LQsXF��(��;2��_�'.��ջ��k �}Ϫǥ��䵀���_!��a@� '%n�іNߧ ��q��ÑW�-��3j�A���ȏ��4�,T�����q9  �{2菥�L�+r��Mu�fH�M���n��r��k�yq�m�O%�ť|�~#����Q֮׉l��.�M{���\��+Y���K��Dz�c�dH��`��\J[�XE�t��F�r܇��j�����) q��CBo���D�x/+�zk�/��ZF�H_z|K0vKbh���f2KM���?}L�H\�ep��/^K6ԫ����Ka�0�=�ԑ+��ٱ�>xP�,�\�1`st<���HzӉY�K��JX�l�Ӱ&��Ús�09�깎u�b���v���\�{.��'! �L�T��V*TL'��#������gM�F��&�E�=ȎĀɺ�,_�V;���K0�i9g�ŭ��k�o[>0���/r "\��vc�qDj��-�����Rw9>>��n�������U���Ip�Qq�jyg��l������z���tރ��2�=����L�P�*}(	c�ح�7�m�<��nfwzO7<��
�^�kc��;�X�P���ݍTے�f���z�l�s샠X,�hO�t��n�E�T(����K�=�NR�/��������]U�TzP��.КsacJ@�9u��̮.������j���,�@��)+�7۵D��g�1bm;d��pn�P���H�9ۻ�>|�[��֊�Wq�l<M=���B%��4��-�X���1Ԓh�4I|�X'��Ѹy�us��π]�S�9�S`�\�xvo*�,E)�O��Ŭ(�<�(�����Ft�����Nz�mi���@=A�^L)�g���
L�BŢ�#�o�2P������>�������,�	������X���͖������k�X�s�V��%�@�����D�r�O�x�k�ZS�@�F=m딓6�5��;���>M<P��̸�MY�:��	�Wt��&�����ۑ~��Ի���$:�����fG����o���$��|&�������*qt�`. #�F+l��2�^X��Y��s�>��|9yz.�o��p��q8ǟ�q @��8��p�l��~��!�/^Rzj��0`�TϞ=�үe0���cT������B����F^|��|���f}���)��7����c9��A�f���</��,��*�����v�݅�b#l�V�Ta%M!�͍�@P��wՙ�t@�#Hx#���V�*Ul�Q%>N�Y��^�ބER	`6@�y5�.�{��$g�i&~��~}H���b�*�^=`�I��W�DH�mWX$,�.D�`P+@�=��f��N�6��.�3n�[T�:�k�{��!��fɵ-�h��X��f���&� (�JQ��� �ڵ�)����� �����}
�j���э�{�+�w>�U/��9&��N������]��}�C�
����paFD�mj��~�Y�� �>p�UԲb������ F����ڕ�^ �r���NC��g���N�c@�#'|ه��ک!<3��#���l���~��s����w  �|GƠ�Gwߺ�^���7�����	��L������L-Ґ�yPq��:��)TႰ�۟��U�Wl����Ļ?��&��;�>�1���Y�u䓁�l
����\����׼���?�U�$�̔����o����x�ġ�+$�}4 -��Y������n	���"���d�t���c�'��T��$�L����H��捾6�bY�r�����R�����L�E��Z�V<t٫�+���c(29�$�aa�ZnV�켾<�K6�G�B�)����ϝ�%�W<<���0�1D4~�*b�� ��$`s l*��;I��	����Ke<��9��y&I��9?�\f���%�5$KK�{��xF��oz�s	3(Ar�*��X�<� Ctm�\�p��?�N���m�}�I�=�'�~�ǖ�Q^J]i�k��|]�:W:��HD&�X��)
0�΁\�����lfb����zAzS"�Tka��j�u�?n �̺���e�A�"	M<|�rY ��X	�\ŉ�& j��Q�죁#H���o����e	G_G~��N����R���SFZ��=	��!���B; �e^�~�k�S������?OυPw�B�m����vA��W�^k1{H���NY̌�_��<�xĹ`XZF	�(��[xN��q�9�8���F@0t�VG�#D�2<�\������{�j�$��)(�&������Ȳh�g����]jX��"�i%�K� v��Yx��6�*�2���Hc�w.O�����J��𙉊ł6b�>�y@y[΢��g�Р�w_n�)�*�[P�������1Ե���q��ʑIV �gH����zPs��Јe�O�����U,����P
W�;���1���n=ں5�rj��Dת�>�n�6�M�ΰ)l��׃�%�a��w��ݫ��D��g�vXQ�b�P�5ӊ d���F�9XV̓�n��x�����V�(`N���^�\CE���+v�=S}��2�4�Z�cԃj*��@nbME找���D�)��O���ؚ��B�^/t����9�8S�$RW���|�R�[�=�ֳ�O������S'f]#3�wd�Yf���u�S���n~|#?�z%_�{�c�|�+9��p�����q8��8�*��򻿓����Feߎj���я.IҋH����ᲥJ"K2y������f����|��O����Ǻ����啼���70A	Y�P� ,�0s�����g����L����6��*Txc���h�k=�3�(�2y�sf��f#ovW��ŏ�1Ɓ���{�>��wCU��Q�M�m���k�=��O/�y��{��otsibش����-7� .`�B��6� �V�A�pȇ$�	��x̘U��*Ec�^�e�I��WT*Ы��.��K룀�g!&+�}��ٝu`��7BI|W�8p�Ul�ւA��2�䍅��%T��@�4�Ϝ�9@��\�����S ��\�۝�޶�ʂ�56��Q�
 T��lֲN��P�
���S���*W^C?sS P@����ɰNRf_�כ�t�Wۮu�G�#�U�Ah�C������K�ui�C � ����Y�{�n6V13Sv;���q����fmx��~o�Zv��5WgB���kOi�RF�v>㍳P�����"`����;"N!��9bS8:�r߷\�nG�����ǀc��ߢ^W���b�z�c��Q'��۹��ݰO�c^*���U�Qh�0�f�d����*d8��"v�a�Uu�Z�f1Ϭ�Y!P�E$Ur��
)��4ۙ�I��G��,@��U	�g�l}��,o�u�(����w�,�+y���v!��L�=�7�7��ؽ�rt��,�VR����9�E:խ���#b�=|/����	0��8g�d��-�C�so!g���S �G�%*�jq���Tm��ΣY q?'2g29��̓X��R�����]c�y{�V���Z�'O��'pw��5���ʤ��.tΨe�<�����(�@s}�Y!�]�Q�7RGS����ɑ$��t&%�Ĳmj��
LzM�ǡ�zY:u�Z��s�ϭ�a�U�d��6_�M�$LjZ\�7��/���::��/�}I��b:��M.ƻZ@�E.���D>�􌊍��F����f�w���X�%r'>D.�d����I�#����!�Y$�N����A6�{w:�0'b!�(w{)*;`����|��t��r?`�[��W�t�C��9�P�2�o�����/���k�����eĘ��m��w�y��簺����Y>���mbK�a�tBE}j�,J(�=� r��U��.��|)�
�o�(�����ʁ�>�l�*Gu�7��=�^C�Q��$��&VVN��	�I�sr��j�Ԃ�����)1�8;���9'���s_�Z� m�d6��u�� �)�wx�X'������Z 9�RA��xe>_���3���&�*��0;dFE�$OϞU��ԁ��(KK�987�@�� Lj�2XY�ym��|� �W���6�4De�H�U;�-#Y:-�02�D�~/K*W꺺FB!T!i�v@v��?�{���l�r�pq�7�Y�ORNA9�L���L��c�?����F6��"2`�esWs*܆�́��T� �+��%;IGC9;9���c�z��>�
��Yqс�9���6��[oVTLǺ�b>X����Ͽ���y��<{�]���_�ɣ3��P�����.f3�1s�i�������n���p��q8ǟ�q @��8��p��G�^�n���Z&�	���n�<�B�NǺ����
�ډ� ��l�wzvNۋIO�Q�,�������믾�?���6��4�|�R1aj���s�j?W:�`zYGȟh(ˇ�(��f l2p�����;�'9~Um�~�����v6 ��!��${X��f�߮Zu��e������9CI}���
u�`8 X���n�$GI��ηV�=< `�
tl�|�,T����U��mQ�,' (eiJR� ����W->$5 �w�K�*�� ����qj
�>�Z�
i-�$u��0��툕�h�]�p@�����ϩE��,��N�N��MePZl��If@��
 �a�;�e�<�W|�����A^�f�/r|�xb� H���bC4sj��	R;_�ܚ�
�H#ME�z�l��ݾ��`V|���i�����^��x'���4]Ho�=ڱtD~"@[����Ŭ���Ћ>N2�]w˕����r����ho��}�C�gOB ���䭻��e�Sk~RMN���,k@~N1��uq�Ȱq�����JW�V��*�ak4Z�D�S� l1�N��) 2�AO�$���6��&iO�3�����R��:ҫm��Kc*2�'��:�I�x���B�:����]�rw���[�S�>�P�$���F������X��*pt:�����b���D��5y=�?K���M?)	خ�ޘ���UL���\�G��cҁ�Y��m��g%�ș[(�屐�� ���ď{��S	�-�C_b�eD���d�3`(�j)����2U��b"��S���"�(��n3[zn�R��,�D��Ahz���ׯr������E!���3�K	��^6�\H�N$\��jVI��⯥
j��IZa.��m���u!�z��A�x����N^�����?�|����GSZ��[��[i�����@M+����E�@8�}���n��MY��*�j�qlB0_ǂW�~�ES�	��kM��Z1B�	H[]�V�%������}�̮Q������9�v�������/�O�Q*[k��_������*�{��^� �d�����w]���}m�y��|�����s���� �{[;Y�����_k��"kIkc�9�'ϩ5K�]M۩+V�<�Ԟ|�,Ǡ��x��yʵ�` ��:?����T+���BV�����r9;< z�\�ã S�m���n.S�ʵ�������i�:,�d����[$vkI�z���=΃sk��)]�T#l����}}�
�,��ڝ��1�����!;>��ٍ�>��j¶�+I-C��97c}�s6�.��fʎ�fYYlM!��$���\�I�W@nw[]�6,�lϢ:�9��b�3[G@t9T�ܺ�\�0�ua������%��6�>Ȭp�b��ɉ����p�����@�N�jx¸��(�}(�/�O���"�/��8�x{uy)o޼�fY�F��.�ه��+#@�����@k�	 �ꧏ���\~|�/f�,O+��d��u�9��f��<;g�ܾ�޳Z����L�w$��I� ��P�q�⧫�o�9��ﻛ[������}�K}��G��_|�c���q8��8�ǁ 9��p����جW�������y�V|j'1Ak�ݴV�]��ݓ�t�0e��X?��u3�Я{v;����W������?��d��P���d�>-� F����x*���	�����Q�Q�  ۣ�3��'ȯ�4�,N�Bo0�1����D>����p#�JzZ;�r2=����������29:1uF/cF�����Q���H_.���H��%� ��!�#���J�J}ߣ�c��Sy�Ѝ�ZV�5�?TV�8� �Ȱ�Y�$c��V_�9�a�RT{k��!�.�"4��dEI5
�,jܟ��E�n�/���l�.�^����0��|�Ya���=@���(3ۣuK#���Y��w�ţ?�Y���EU�X��p0��9 ���/�sh��N1B�ڬ���t 3���>d�@0�;*à$؆M���z�J_ڄ �9@!��Mٓ r�I����Y��J����P�,3b+wQ &=S���g�d�Px�<��*�뀈P������'W!�y��svvO �@V��dڤ�E{R��"G�$�
E���ݭ������CO��̓x^��G���#��}�z�u���~�lt �y�h��T$��.��P���vn#�%�wê�ʭ��L@�*�(��`��U�@_�U��d�kt��b#Poa����jG<
��	�_K���b��r!��@��
���\u䇁��v�����}eu��F�)D�0ə���������\^_��t�<���ɓ+�ɑ�������,�/%,q.=m��Lc��R~�J7�οIU�e/��'��j�1x:�-̈\u��{SQMz:/��qr-q�M�'-�#&M�@�"��5��_x���` A�V����$��U΍���*���ܾ5�rZZA�����GZ/�{���o���K=���:�P<��� }6���,��%?R����`ϧӴ�CsI�^���c��F��؟����t����!�B쒫]-˅~-sy�L����FۻlY,V�.7�?=�3���KO���$lt-�oH�v�8>�g�~vLU.������/�Ʉ_��2�r� ���,}"}�T��^7u>��C�������.JL*�hggk���Z��6 L��"��B�QN%��h�'�˺�2�Q��lM�l�HއbԎG� ����� �7 ����H.�'`��6
*�\���='	���>x_���� �%}|��f�F2YNVyЪ��
�d�g��Y|���؀{�a8j_�[�^$����)� ��֪�?1��F�h�y�>.dn��c�C%��~�Ĝ]�Yg�y�5|�e���kB���B<S8H�7+A�2-'��+�u$�=���jG[;+�40��wYR6g��x�u��ID@= b�A�]�Ai����<roERp�ǳ��E\g�JXd�YN�>�Uu��!)m�me�Yl��f��[�2c��-�/f��k5���t(��,��v��=G	�\����XX��Saଯ�zo��29�Ԑ�Mk�PV����続�VK2��G�(���oSh���T�?���r��3y����L�Ndzz&�of�]�f$��6xv a��yntX����S����"��G��d����3=ױ�͔6oFruVv[&1L^^� ����������2�L9��>G�j;,��Hn�@�T�4O�}�Fl�sy�ϸx��,U������8��p�?��@���q8���Y��r�?F����歼�|!�m��nl%AntU�m�,&�Y�����o�����,s�s_�|%�~�Gn�����������~"b~T���h�0�,�׷�� �Sm�qc���2� )њu �8'�UB���9����Ӛk26��p����{�
���O�믾���vS�>mJ�rE�Ȍ.����\B) �&M3��-����J��FX|���٩�'#����KJQeYu�
��l)�+Q�Z9EFC�+*[ 6F(��C� (���� ��aS��MTx�l����d�t�eR���}��"���$pa�[fW �!��y����{8��B ��5��}؇x��O�H�C� K��/��bg���6"�DT�}������|G�3<Ǧ�C��A�����]b�;�K����oo��x���R;O{|n��1�I�jHV���7�J�َ�>K< mY�����7���/I��aON�H)�&�b�2((��3T13�2�.�@ ����	�+���{�fB����˷�� _��w:���j[Z`���6_P\^�)�T�z�`T�!� =��ڷ��n��My��&6���V�2��������Ux�Ե5�s�V�Y��iYP��b�j����9�
_�����bAΒ���U;ɷK}-HB�ܗ����32 ��	�	6ه1X~�#
<+j"��াp!� P��5@��Z��wY�ҟ�+��Lǥ�ޓ����[Y��p���������sb�PE�P���K�k}�G��N���X��5��֡9��5�9�ʿ9ouʬ��91�#~�(	ؽDFE��
t^��\��6������ኪ��<�uA�Q�8��!A�8�]�ss���3��~�M(�hQmL��0 U��jS�<\�DZjs�����[ ����P�ނb����h���,E<��h��tą��B�oky�ƲD�1�?A�ִ�*�ձ�l7����
�V������3k�j��j��銝}�lh�c ��U�@��y|1�<���HS;`=lu
���c!�̇�ڊy�<5����86�?ύS���lB���� /�.dK���<�,������6�vJ4�+��p���U��U m��a�6�ER�r��		�:gܾ��< ���L��؀��s����=�81o��.�9�'��"̵��̺J�M ��9�ULX�m3�"�KY�����$c[�S��E+�劤D�3쭠�������<FN`]�h{ɹܷ5֞6�S�0���<Զy>�>��g��sz�W�t9���d��OڟJg��,�>���85{�v?�5.��lź��y� ������{Vt����첞�������v�>ш��?�T���Fo�,xƀ"�����fME	ȩ^�s�C<?8;-N$��%�e�
:ڽ�m�0�1��Z	�	T\�ϸ�b��{U~+�L��h�3�J��/�<��%۽�j��A��gPx&��D�=���<c1N�q�kA�y|�X��3�YU����ko߾���+Z:"3h�>�+�ϊ�<S}�v�P����	�Cm]��]���}���h��c����/����}�&�|��c�'�¶�ME����y2=��.gۼ}���s��\��nu��R~���� ��p���'��q8��8?�@�����}!��+�a���l���tb�
`E����l����+������w��{��np����Wr{}eUj �{�lt3���L���-�U��r"N$߮e��s������|���z`/�	�s\� ���G�&�&��c6ັ�����L�={&Sݘ!t|�Z���cC��v����$���mi;��A0���'	�kj�v+���I?p�Х�P[���I�<�sz�å�n����90ͅh�z��&�dd�9�CK�p��h2%��崠�#(�k�!v>������(�@V����p���#E�:w�͹y�
���Ԋ�u�y����Ț-.롡z�@9�:���0�w�
���[ }�O��ǰYV�	�AM+���~���;*������1?�֪DiRSy�&����\����QY^l�$C��p�O�� �,����.�7�@q fo��R�ڷQ%NTL� ��Vɝ�B*5�oq�a��זp�&�s	^�����~���� ;z����2�Wz-��H ��� ��ڭ*a�	UH ���{��o��������<b���!�f^_^S��^~|4aN���T�������C�-�8X�y.���.'ď�_�r�afU�1U���@9�6�_��<IJ��e�j׎ �!Ҵ����B���١�I��]S�;������f�Y/��u.k�tlZIF�
Z�)�k)J*00�[ z:����:���K�П7Ֆv: g1v:�]���e!W���X;��3"�6�ϼ�)�ڞ_ �[�:�>��W2��h,��Fg�.�ݏ+�����\D#٭��1ڃ] @d6!�6���s��-wZ���K*z^���{.�z�A��c�uC֥�I���d��a���YQ�b��+��b@:��zU:?޼~.dNž�A�<0#�Gס�S��R
m.1��<_�R�d���Ɓ:U�����K��y{v)�t+��HB�eQ�>j��,���4ā�]>
��pIqR��{]�sy��kM{2���[	��B��(`���9�ԥ�}��W��g�$נLX�c�>_�g����a��X(6ڏ�lJ۫�z-�s�o:5��1o�X��V9��Y�D��*�AA�lO�M�?jr���v��/p� � ����!�I��c#�i�d��T_�p���8�=�l�����̕�InVa��-�,��srXT�̄�`H˺�[����\��
(�P]����h}���ky6x�^o(}��_rD5灰������=T�lu΄RŔ�	r�8�Ev� �SmK���M����ye8�J6��L�π@k��В�'t��-�xq+��B��)�G�<qA�K�FO�~0:b�xg�êc�(a���;��8n��Q��@<7x��3v2NI&���a.�s���(TU��@�Ld����4�u����o�Ԩ�j���1J�6��C� �:����n�+P���lx˒�
OtnnNNH\�^��\�y �b�	L�E���h�U[a�N����wĺ�Z����dm��E�}���g��ـ��i۩m��0`�)QqVs��ù�ρ81��g�V_@�N����֭''G��)�A��d�R�7�u_���ј�-rY�|��}��I���HChx�a������J�\_��7�i���x �E�)�����k������>�P�Ɉ�4��hC��u}}�!�޷�|�:.F���V���{���+{�1=~��_��8��p�?��@���q8����Z1�P�P��� T!�H�B�G|����<��1e~��In�*ݬ�F����C� ���i/!�_�fn[le��oTk�Fc�L��H��&�^�$P�]8�6�!�BjZd��&����~���Q$�d�uV�*���z~(p�fa��n� MF�|n6[��k3oe� ���j�����|��/��}%86� �i7�� 8M��6� T��a6$Ŷ��8��v-�>��'  v8_u �@5!+�+���h��=H��]5�U����m<Qu�
�yx���z{5�7o��o@�q��O`�yN�a`�g!��uӍ���V�r_	��#X�q�ܸ��B "�� 0�s�>������&���p���m]��o�D1���w��F�]�P[�C�}���_���@���``S/`<������5��@π�b������QT�/�0Aݦ�:�|�"���	j�����T��S���)*����|��%�h�Þc�үmC�*���f@�a�I.��� ��?�i�Jn�� A�{�[���Z�
�{opm��� 'b')��.�����'� ( �+�S�C**�)o6M]�-^WU�$�F�n�-��g#�S�U~�J[j��D�+��a�^ZnK٭�^��B����!�#�K5����}��l@U}���j}��a`7H�ma�"�Ζ�ۂh�ߋd���D��Y&P-h�A���	d���v&rw����ec͎
?��qV�ኑ�R���,��ʱҸ�'�y3��*�[��v:&r#@�� Q��mV��n��Ϩ��0�o����Y,;z��`%��N��^���/��+OG�������
w-,�@�!�EϿ?��ي���a[F��XO)����K�/��R�ғ��Z�݆���4 Џe|T�r|���q���d[m���W_2о.�{~_�a���#��8L÷�>��--��s��1j]�����:�m��
��o�F��k�[*cx��D����~$Ux���������^!Fq]e�'��8�QզD�B����.�v����<���@q �m�xAs@��m�l}S���`-�T�]QlʔN����u��C��JA��zP��,�ڜ>�	�жuŋt��l�a��)'h�5�@b��5VF�(�|\�`t���7-�&`�Ҡ��3�B?��ܙ�����F�_�cq�lY��{�S�������� ��)7<�g��P���[*{@A�G"��:��F��&YܓPa�uϳ0����O��5�ܧ:C�9Nz} � p}���ܨs�x1ۉ�,{~�5��0ռF(�|g�k��Q
�nc�\�XY|���c�8|�o�yC��\���{�1 /��$`�v��u��0+��g����.���{_>O	l-��9ӱ��y3���:�M�܃�|��:�GKA�5H�_\\�������I��6�bq�����B�y���)+A��wzx��s���}�)�Z�_�mO�9�]���,ܒ��bx>�u\�ۓʓg��/>�T�y�}9:9�}g��0���Y��Bы1�{�+�4��=g���q�D>��3�lq-��|�ٯ��q8���38��8��p���X���Ջ��8�7t�r��Zn�J�!���Hڝ��� (�nt@~������*�P�����0@v�\rC\�5+�˦��+���Z�0���o�X�;==&��&��2o얠z��\Zy�{���a�*�a����Y�hA.���hAA��=�@@���#���}���  _�7+�E�>��	ڮ��'qf�;^�p��6�)+�͂
�B�_k ̹��I�)X<+�ׯ�S](�U� B% a =�B������A�4.��n\�)p��������
`��{�q @Wm�� Cc[�ȩG�̧v�@|w ���B]nn��~[?�?�m�'5b�<1*�I\��<�Le4�0�.6�]��c�D��B��L�`��7�	z�j8,��,O�$��w���~e L-��H����J��������|��B�� =��%|�l�G�e�$�j���
��J�~LU��VWPWpT�$�1��3ك�5-�Z�����-�G�n ժ����Q<������kA߀�T�Bj+o�����9������z�=;�V` qI
�]3�
���Fc'�n��B-T8 dY�Op�gF�O�+d#�q��+N����>�zK����1�3?0k C��-�j wA�A.Q�s����jo�d�&ky� jo����g�K,߁ \��T;�:�f�;�9$!-���W�/��); 6��PR�l�z)6�j�d����f=ɫ� wE�0
��􇡾]��|�7uA�Pg �*GP9��MTh;��j���6����[��)Fv�&[5�y%�1������_;W'w7&he��O������ex[��,^_��/���Q���7���d8��k����5� ��2�L�x^�,�9m�J���,���c��l�����}�w3�v+Z��^+E惾��c�V�yΜ�f���T'�1x��\����[�b��L�b%�!,��~0/��t�-l�}>��%�ܶ$h�����r��]���\�k}����@��P�=������֍驂q�:�#¼���@�5�k,*��PWޣ<vvF����	�*_\���Um ,�w#G ��T~̯��K]�P���k�.\�k�,����l[�0_b���Z�.��@��߆�/��`���N���6�y�}D�J���a�6$Wѿqs����w<���Wv�q����CXl%��Ϭ]� �'�5�R��GR"�k�;�U�Cy��������l�5s4��g@5�.�/�b���}���� g#{/fO�� ;��hB��S�m����(j�ثC�g!	��TA,���fA���`"s�XۑIu �c����D!CL�G��ɥ���	�FD�v��s�B��]%�y��עH�ٔҮ���ֱ��LӺ��mx>`��O�����K��4�*��0(S��bJ1�WB���z�s�O��|V�T7��w��`oB��on|~_��~/������ޑ��#�Lp�J���������P瑠���u�I��Q���x���-�mw���٠������s|V"1��Y��C�)I\7|�8yt*��7!�|�+���҆�gZ��}{�c?�7*w[�L��_��O{V/t��y����'_~�{���_���8����8 ��p��q8~�� ^ë�
̻Z�d:�0�q~sK# ����؞n���V�\�Ôo�}w�ʶ��zG�6�}݈m	#���52|�����w^�ɾz��Zpj~�l���Mv����U�K�*��%�1#,������pec , ̞+t���A�]u�%#h᳢�U�J�вh�U�w�/z],�^�G������Kn���8Z�λ cWS�9�~��T��#e%�"�b�]�'.|�x�;q� ����` ���œ����{"�d
𥰥-W{K	҅��u�re2ɐU��L�&r~~F2�;�v{5 �9Q��U�����xKo��H�1�R�\�P�?����W˵�,zN�8�-p �yVA0�f�*pQ�B���~Q9����2�S�,�Ї-L�e��dd�iq���=�3�Guv���l��v����d`�	��&PXe-+�ۊ��;gQ��c��Ǌ�rPV�3xX�
������`;���_�z������J U��>��	���}���bT��^&L-ܸ1UK�Z�r�cQ�@DE�Z&�*G���:P�#Gu����ti����e�n@R����$��u��[�~"����M,;6p��'����O���V�ڮ���k�*hT<O��Z.V�#2з��B͑��w$o/n�u����:N�\��
��J�nL�����(��O����֬p���&g��Fڝ{bR+�!;�=%2/Ne��i�O��$a����ۂ௠��L��S���Z�������SR�Jh_d�+A����@߷�Mo�wr������\�W��_X|F��j������P��d��}N����OE�ի9�Ev��%a�r��\R=�a_t��t|���a5�!�shk�h$�s@�
�<O�!Q��yE?�d*z/9��\���H�ͼ ���$c���L�V�*t����^|3 @ZutP���r��U��5{�ͺ]�<�`#2<4�����*!�5��]�O�����$��Co�j�ظqG��օ��n�9�
5�-��s�o�?�!������a��S�.�1PIG$X�8M��Jӳyc�A��^1�1f�x��
�+�m�b�Tu��^]�.��r67{#�R]gG���hi6�5?��JG�{.�� l���`��fN2Vr�I8��y�_׻�ف���`,���ї_~)���e2>a�����S��3jp� 3�����W�^ӢJS�>&�	I���W�oh�B�x:%%po	�c]l���5��\��}�E�g�]�Eט��`8�',���uf�R[�KJ���z��al�`b��K���S�v
����ݒ�ǿC*u}�?-���!�]��B���L)]�,�9�)k���bsT���0$t��;��Z��"ŭ��L��
Г��Nk:��N8�)@@��$��^,��Yn��,�B�;#�cw��.��t'ٶ��P0�k4�ˣ�c99�矦)$_-%/א�ꔬϯ����4�%߂�1�R����vSz꜡�֍�Wɤ��Y��f��s��s-��ڗ|O�&����  Ep���|��g����z~l��
���y{)��;"�Ÿ�c`�f��9;�e|�F��yt4�_}������8��p���p��q8��v���ŚЪ��a]�;��Pƣ1�|�,�}��lPt��`mx��LXS݌E�r��W�hu37�J���n�wE�L�����O,�6��0�dl�A� ��z~/a ���sa���x�mB�˽�N�x�Z���3D�+ l�V�-��M� t���	�s�⠨tn]�a���U�� ��*�6� Q�FBe(Im�����jGs(*���s�y����3��-Dc��Q�
IT��[˫����<ZC�8��uv��%�#t\;VFd��@u��3�\_[�=B��5��$�T9"y�Pb��7���b�c�A�j����<:9e���Y���]{�9țI���U=!��b���*7���2A"]3�ق�-X�3��ix����X/�V���v��m�^�槡W=�`Ue�ǑAa��r�}�CS��k�pe�&I�-��mE>,B52H��E 6�C��G5���S� &,��)p���j�j`�Mi�o�����zQ-���l��lw�� ����� ��ݠ��h��J���G999�gO�af�8X���Y]�ޓ[>~��dT���+�ũ�@x�{�G���
-s0�Q�
���+la��;��R}��Y_׷�klx\9��'�ٿ�ǟ���0e�	�@�z�*�3V�#�`ZB��U��:��z��f��-un��`<1��$��� cG���l��x#77�i�[��o$�f���_����界��$��v��0%x�V��\�|~#'��������L���T��+������KXf�0�c�w;%N��k|ǘa|��S p�e?�OT���v~���KP!�Ad�����^C"�������\/��Wp1���������NN&"��"�' `[�9`#+]7f798)����z�$�T&~Ā�6�e5Y#d%��4���(��  ��d��1�.�����9r=.蛵�R�{]Lt<������-��N�|�)�I�<{�.�����+=���&G��>Վ�}���R^[%> Z�/�ԟ��Ȑ��s���Ĺ�  .��J�[�O�Z�&��S����}���)�ʮ�͎�!�3���8���g�y�ٚ�0vּ��FfSksq+V�u8��ܕ��'H��M�q�X�jy���=(-3�I�ZP:i m�N��{����z
��m��h$�|�s��b}��7r��5�ad9�Hn�P�,�q�y��s�1k�8����T��"ԁ9�5(|��6���%�����זu��<L{}9>='psu+_���������	�g4ֱ.���\R���}Q��z��o��N�ur9:>�����I��\�+�����3]3~��<�\|�a�zkj�?5M+�T��}Lk-؈%�'�ʪtk��h�Iip��=}W|�Ӽo<l�����:�ٖa|�E�ٯ
���1��@�~T�E�~����e��Nk!���|�x��2n�;ۺ$4eS��UA%U��?�w��y���;B%��V�"��*G6�zT��m]YQ��܄g ܛ.��s!%��J���}zt,�g��2��b�0+}yrX����yaz2 2v 4j!QV�}Cch��<[�@�d֜%.���k_f��9���:��ə|��_ɻ���A��8�������?j?�Z����3����ϩ�ѱ�j�<{|!���|����Q���<{*��p��q8���r8��8��g?|g�U�[z�����fE�Ve�f	^�x*�@Y�>�<!�X� h���N7�cy�Ï긚�������9I�PA�&߷jWϳ|��r���a��<"����ٻ����t�Z�A j�v�N��(IB`c>�R����kG��8����n:Q�ZT{[ %TY��VR��?��nX�^�e>_�@% T�nJW"���`�p11�d��=���
+|l�˜�r��~'�M,�-����(�ܨ�*��d2KO~�3o-l�T"���i�,:�C�������rf�Ժ������ ��>�f�C��u�5����*1X�Y=@�aNV����r��2!J�aӒ ��j�Φ����޵�~�-2�&
}
�P����	��~�YD�0�P� 0	����@�XHpg[�s�5<�} �TZX;��U_֍�KG��oűO��rf̧[ (�#[����!���e�f���Η��h7�
M���f+�"C�)�J�ꏊ�Ha0*:�u y#��Z�HI�J8%��Z\�yk�IOgߣ��s����d���ڳ܎¬x`��MY	��dn�|+L�h=��h��N���%��w�xFx�ek�: �B���׶�ah�E���b_)+D�#(�,t�Y$O[* ��њ�	~����^��0�@�}:B���{.�_����j*�wru#������or�~!��Zn���g5S��?�ys%W�oe1+\�v ���cOU.iO_�<���o^�)T:��K;w�9�Y,m݁^�����Y��=S���3�ǳ��ƫHh�=�b&U�A׉UC���g���v����=�ɤ��F�⭬�����>ȏ���L'�+IC�J�(H~�n9�oo�H2A�f&l�7)��qي$&��#�)�E�J�� ��+߳b�ˁG�| ��J7WR�W�ŔF@��;�;�_�`˸�s��Yh�M^I��e~g!�^\���z�9C��m$� ��J|(Ę���;I$���m�G@�:��͜���$`q�^��������QOGI�J� � ��˗�:�6vYo���9�o��yz�x&�n1ׁ p��rB t�C�#Ać��'��w��[� r����1��N8Ay`�������ӹ���+<���y�j�5�1P��i�\��@�i�,\7����z�\��]�8�$�AP\�!��{�>}W�	�WP��sÜȌP�\^���?���ou�.f�~���*���X�,�{� ��=��>��c~YKK"��B��z�&Y���%C�O&�\k��� oAxw��ېkR�OkL�珇��Jӌ�;��}�W7���O��4�ߩP���\!�M��0���ҬJi=�g���}�$Z�9�YfVV����T�+nh��O�"�!z�>ߣ�Bֻg��2��B��뤲k��v�x�D]�?�tG������P��9��ީ�_������C1�����֩��%�+,�q����Ԇ��P�>;�����/]Ϡ-�[VӒ�u�i��	���]dx-�p�Ȧ�X�uT�5{��I�iYW�9VN��0����I�1�9���<}��GcSz�k`��������?����/�T�$�_��D5�G:�\�z��;̿��8��xDE�?�����_�����8��p���'{��q8��8�:l��Icnrngs�^I`��(��=�3w5@�Bvۊ�:2`��d=S��ft4��?����o�G��G���5+�b�\]�F7l L��|��Q�jn���]U�T͡Za��X�H��#�F<�M�YTA�yi��OQ�[�]��A�(��](�K�B"Q}0�³=L](��M.��\���2���jl��*	i�M=�  � ��I�!��YD.`j((Xa�X8h �p %��Ӎe[���3��ê��`�{r��"!�ɭ7"�v �+|�����	�[zڎ�g� �-��a���J�m�V�&��F�k��Cݵ3~'�>��CԵ��g��E3n�⊊iXLAi��F���A�a �e^���롿�{W5v#�¾�v,�ϐ蓄 �Ȱ����`�f	�%��e�C�}F[5f�� ���6@�m����մ��2�) �Y���c� �TT��B�]hlMҠf�|I�G����-e[�2���q"�]C�'s߱��?�x];�e����^o"i6d0I����7#@]Ս\�#� v�7��Ţi�$fr|�u=���\�m[f0N��V�;¶�<V���*Y�1��[�47 u���4�r�}c�oD�IS�w�ɬ����Z#�7�،��DTxx�h�50��s*�#o#Q?��'���X_��������ۅ���f���p,�9 �Tw;��]��ە�n ���g"�a!��e=�,��G�Q-�m!��k�G2�ϝw�B�Z�q�}�w}���p(a�0]w�e]���Α��[Z!q�K�C�Y�����\ϱ�J#��c}�P�R�:H6K�I��eq{%w��׃(���L&�P�X�T������Z�\
I������sI�Gzˠ~ӓ���Bze�k�ZZ˻������[��Y��N�oeA�Ȅ�mJ�V�D'��3�u�3��=¸\K�m
1MO��͢~�~�g>/ľs�8�k���HdpD�?����� aOT�k�y���<�dvdZm7{�6�I�:H��뉧��,=�2t�Az� ˡ 8�p��	�G�q�I@ґO,�Cyv>��)���*��$�#v'�2�U}�<�̢�Ht�#�n$@�l�9� W�%��}��Pͮk�d:���3��c/M����ܮ'O�ɣ���&B	PW��ܙO���ŝ�VK0�I����K�T'2ֹ���V��5��qY '�s��O�^H���%MF��|eVR���������A��)�f��E���hd���5U��ט��Vnnnd~��u��cX=�iV���nwT��i�e�|�B��o�^@u t�Ӓ����~˱���v</�>[Q���p��E r����|]���;���kN`�%<#I��3�l.��o���a�C�Q:s,+�hܚ�3F�<�d���gW|v�]�W@A��B�Β�b�ZW��/����'T0���)�Y��rʞ�r��a�:��DO�h��e���)�Z�[>�\1׶� ��̍]�^U&%�m��Q��\<���4b�=,Ɛ+�sZm6���{P�yQ��X����#�*]�ARA�x�h˪�aI�r�p2 L6��l�Z["�&����D�o��i���
n<�.����/��'��/e�\h�u���z����/��?�t�B��?�^>��3y��=[�,��~������q8����?��8��p����,�J����n��#� pTQ��VE�-�v��9���3[7���\J�,B���W����V�}�]y��sy��������-7\�n� R�z�>+�}�I4ogo� PV9G�!+���f܀{��A�ji��	�ăU��Ei`�l0# �`dM�b*;␛�}�+7Ǯ�a�V	���A�T2�H�}P-`��u���HG����:�ڣ,aE$���8�@�(�@�>��  ���¿�{҃G��m-��o?�~� �{��] rh�	Ʌ.S�H�fui��N%��g�&^�;P�5�Lky�G��@�w@P�����}x3T��^�]U���P�HCO��O�;-{��п������3�H��\X| [c�� N|Z���+�M�|K���~���� Юӣ1���̵�^��"���Ta����8�h�B!�̓��ZR�?{c@d�����网l�P���TKծ���kH�Ж�Lh�B��=�$J@�}�g�,5P�I�R?�*���AϷi�*J(?�|�
��j&��Z�z���}��� DpSt	@�$��| ��-I�+5��Ty�jr	d�+�NE���Y��p���0��2@,��6���� -{Sˊ�jgDc�y��`B�v.�)I�g�!�[ �u��t~.�aKZ���ޠ#�(�  ��IDAT\~H X�i{hҿ��o��+���J?��=H��S�����͵O��]	�*N�3��گ1��<7���^��e1�@���G^^�d8�u<dz�Hz�\���|w)��Gz�d��]���Z?$�F�jb���2�`���{ŉS�y��
�'��5	�cK�R�s=�9y	��\'��L�׋���ɐ�G��Q%Q߲0R�U�c1ؑ�Z�\_���bx4е�L����Q�G����2�_!��sm���tz݃�'l�b�J��D�\����i�>����KYlby?Jr2�5צ[�p.)��t^@}�,� s]�혋��J.��l|�.z.���>�P��$�F���T���fM5X(ǀ@���.|�#�J�h��f���j�]�~Oo[J���-��tm{no��	̴
;�@�׃�@�CI��ǹS�B��U��c 4�B�K����r��u��d��x˔�۸��'1��'��F�V���*s6�ܪ��__&ӱ\<9�9vJ����7��b�s>��`E����`rD;��Ώw��2�I#�7w���
M��ȱ )��� �����y��Z��3��s�  �X��0o�=��@˅�=��;�{aqx;����+���Oi�W���L�n�x2��x*��gzOb*Y��h�^�&X��d8�<	u췲�G2	v��8��"+%�YE�Y���#�zC�/x6*�\Ź��Mfpo�I��'P�ۜ
��yo��;��{-?�5@僙��-	���X���� ��l��4ڕAi���vӊ�3������bgsj�j	�Xl�b��Ѕs�#D�5�ޣ#Y�g�����B���]���\P0ᚬ���?,T��i�gG��ˏ�3�^�@�dDR�g�����l�-�����|�u϶A�1 �ǐ�`����A��3��@w�ݳח�:��̵�> B�1�F\�{�U��^�23$��N�MK����-�D���l���@�i���=:/�6���uկC����/��B�ڗ�85=ۋ]M9̝��a3s��f�CN�{������Z�� #��Pc�1$\u�dʊ5��r!�~/p�2(}_��[��c9�c9�c��/G �X��X��X��� ��������٣�����>8�"�	8d޼��a��l&��>��R��3�qZ�裏�����ԧ�S����3`�t SVA\ΤI ���,�̠�iT]���n���G3��_.������siBi���5�MPƘ�!�(=��H^|���y(ۉwrf�����ؐ.ʙ��1�ƾ��z�O���l�L�&�#���&(\G�옋G�(m�\� !3MvǞ�����8�
��=� F�%�а����^I�m6�����z�ՃhV��u�����<3�.p�KG�HV x��l��� ���"8_���G�e�l��e�S�A�^�cst.���\j����)����c��|��Ԙ��1nR��*z�)����nN?���W��~-��} 8BY}& y���sh���E]J���SɌd0!�Ҙ��˦��G�V�]�}���#J� Hrr~Ƭ��3Y������g���������ӓS�u�g�����  ]`��~�rͣ������$}3wE0���5����K��8�7N�:����F}�=�B��'ܷ'lW�$� �T[���g*���uw������B3 ��t�k��n˳���V���� ��h� #�c����n�KP��&c����{B��`^ˀ>�g�L��C4- 'He�|�N����^�g��w�C���A�33%q�+�˼��U%:�&�pce<�gv��RA���;n�[�;s<K����GM��Qbmό�1^�K=f�2��k��K�/v��[	TB��F�TƏ҃ŇN��|�����Q��V 5dD*�F�[��-�D>��}�8����ꅬ��>H�ep�L�����ߎ%b���z!Z;R&0�F�*en���S��4��@�}�kq�sd�!���$A���d��nC�@F{���D" �Z��_������#�<��KIou,���sy���y ��ѹzE&��ه�N$�5	V����ˉԛK�t�U�\�N��t�s��%K_��|��X�d6�	�ݼ����z�X~�˟
�H�����R�q�-�i���%Ye%��nJxY �p��ߵ���&&�4xqv�$+!��Ț���>$� �ܱ
�=C�ĉ��槑���5h)%�)/��/u�&2� lB��vG���@�ƚ���ى1�5	��P�<
=k��"� �C���U��W�}����,)�g��)*�{��b�+�� �h `a�L��@]���B�@'�}2�
��؄�
��z���ܚ�pdN�=���n��Ӄ�\:����|-��F |�#��׵@�y�{.��>�5�+��`o#]w�~���Ɍ����D2��rOV�Jn�B�/��G��JZ��n�FÜ�����~��D�����{+����k��|�}�?i?��
�����D[��1�u��y1׺��#ͦ:OO��	n0Rt�&�00&$�-�U��l�R`����`/�0�x�9�d7�m���9�a�CNtK8��=�ױ��4����Q��oc�I���L��x6HR�a�؆{�2bMr�mS}W�ӻ���h��k� ���`6��c��x?��;�́��4��������$���^�yj`�E�77W���9��H�-3�'�tά}�N)Q�X�(#�	Tf[�#&�@&��VYlR��Q'P|�s�+��7��Þ�m�{�^�.���^n��OJ�t.ZS����$�~W�`����?0��C�^J�T2}/x�`}��@�`8Ɲ��]eL$��t��uN�Cnt[��#,�C�#�}�v�.��p��({u,�r,��U� ȱ˱˱��
�w�7��?��#���?�����a�p C�Y�8(��gà�H��و����<E&������hB;)� ���Hm��,��R999уtj���CpU,��4��y�.�ѻ|�C�n��A��bYv=�����Ļ��P�5�a��
�EA� �����jَ>��(��03O� �Z/�Wd����Є4�3P:)pٖ��1cR�\��cA ��&"���]�PZ�y�C��FF]�Dǁ1��-Y;`�t��8�#��""�f�=/��1�ʞ�+3�#jI*g���xm�.�������8�I�l��6���2{4�b'���[����l���l�g���٪�{'��@���/���[]"p�|v#H/����|~줾������4�ύG��0��`��q�j%l tAP���j�f����6N�%�m'3�f �o��6�'�m&�d �%����2P��p������Q:�a�2[���X
�/��򻙽O��=���w��}?|Ȃh�#`�y^3�����  �^o�l�42)Hp�h7(�زGK��2}�_0/�v�ˀ�n�X�1�`i�Nҫ��,����QY6y[�A|h&�$����A01p�4 &��Y���8~�C��;�@��xӞ�ާ��[�dLb��W�vRo��mq]��������i��?��5���|��_ �k!�/����:g�S2NP��~��h��i��6(��숥0`�e�$����s��|�ɾ�h��I4|"�~-��hם����{�[Rά�L���T��,f�d�f���b�ׁ3<qE�g���>�l�����l+����B���N�0#��	M�5hM����xe���F�ۆ��n-�{}=j��;��Z�G2<}�sR�}�q�I󵤣�V�١�S�\{u]��W�\�� �x3{`�$�Y#/��RF:V�O>�3��m&�#�Y�Q�_D����"�y#���b�Ϩ�`���:��s<�3`H����%ڏ��Z4rу���u�����F�)2���|!a�'��S�[z[@:��ڑ�ZE!D9��6[�z4�
�@�x뜑Ķ��Gה�D!�. ��Cک�KG�L�[g�]�	r?�f!(�5�k/>�9�����~��X���e���h��?�~8�:�N@&<@sx��t^�W���P�AA��(P����t2  n�B��)�������F�V�9DfQ�d/0�%����'�G�x23Ct}0��h��'܏�'C��i,��F2�5�kL��bO�����������Y�d��KV<a�`Oƌz�� �v;�;��ؓam$+�r���K��U��
:�%;�>T��Ι�s8�O��&��=Eg�;����O�@�����Z��+Jb!y���B�r�S�>���~� ���ha�o�-���ݕ�`fK�o���F�	(`��}�`�6d�]���������Xß=��%H�i�O�Mr`+��üq�4�0i�4�Z.��l�/J���sb��c�I	Ų�=#';�ߛw�%�5+�?c��&K����}�8B�
��5�D$ �����*d�2Ǭ	��~�>�	�?�/�7Ƅ�دr��j����gȌ껔:�Ѷ � C;���.���n�(I2����>.��먗�ٙ�Z������r,�r,9��˱˱˟�P�����L~������7�^�.�Hl�~2͝i�ڙI*u漢�L��Ђ�Y�R��F����Ȝ�Mв.ļ�}$���
\N�9j��9�&�-� J?�OJ@�=0�]�B�
g}������oa����+y��5���a��ds��v>��B@�?�3@�Æ�_�@��!���*� ��D���;
�)	R3���ס6#oO8@fd@���9 S<=������}+��@>0��F��f��駎RU�׏ށ"MmAx� 0)��L�� >�y�X[Ŧ^�P����I�8e�[�-33C�wREN_>�
y/�e� B`:�� �#{t C}���8�}�i���Cگx��j���LȅJ-�ہ�sz *��<~h�s�s�LQ�m��trv*�ى�I$#�?��,�3�1����.k�B�w���A�����`J| �j����<�H-{���{.�t0�O1��DrRp�F;z� �[i?�1�0��ի���@��b����{�D��>��< ?dto�{2V�	��nHV��%���ę�V4�m�
J�����$���g�Z�dd��L �r�a�m� T|P֪3u)d��&�y�h/_�-;��R� @2��53�C�
z��&S�� $;H{������ tPc&0O�xΪsF�`�Ѡp����7���� �fQE�:�́1���'E}&��T���H\�Kgڦ�F?�f������Y��˫����~��{}�Gg�r�Y/�N#�ڱ��^��C���ڶ�Rg7:]kUed�DvZ�Eb��� =4�y�Ʉ��dwh}ƮG��
���D1LCmH����`ed��߁5t#���t.&�]�;��t|�:�joր�2I$�}�߻mq1`"���`l��l�V^�
�G������W��_�֣D=�0!��I���>�r]�ݭV�F���y@��@\��2Y�k]-�\R �'�x��^����h,��	=��sbs�vz#Y�@�B�Sң�RK!���HP%��{��@~��~'W�Lخ�h�JT��H[��7�\�3��x,'��ɍ�p4�d^a�BMw0J�����2�#24�o���@��3 ���`��9��<�0����|$�$��F���}7����ZB^I����π=<����0>�:ښ�XHX������!�AZ���d���,9�Ϡ�~��>[}<��?��=ȓa��rx�F��<���FN��>�Ie�QǱo��D?���e��e�!��&qBYC\��z�� ���~����}n�J3��R^�7x��pD�]��$������ O����[�@��j,�$��իl�K
lN�6R����(ZS���}n`�Bܽ���l�'"���t���>�/k�����}Pd{�Ij�q��d
��XwS�i�K��u�@�s��]��_�ލ'S��`{@&A  �Z;��9x�$?1����A*B�:v �d���Ս<}�~�?��2�!���w��V�=�1�$�����'6�͸�u_�&�C`��N���MRr��PV���K���R��-Y/:TA;F�G�>I˛�����#b�o�31$����Z� '1��ͥ�s����?h�g�~��\2�V�<�h_��C������y�?��gϹN�Q����˱˱��# r,�r,�r,�2�e����dz!~����6�]�'`a�$���&/̄ۋa�1(����$A�Ь��p��(?&���z�&�`٢=j����4,���"�b��˘^�W<(?~�����x�LR*;d�A~J�y����_������tJ�>��# �̃!8��5��/$���%�F���6��Й��-N��ى����X�����/x0�N�=�K ��#��Π�s�o��dR� Oc��yw (�������Trz��1`� ��l���Z/�p�(��6�����!`O���b ��i��d����a]x��{��2i�У���L�!exX���Rw���B멳lS��#��؎����Gq�#� �t���w��c@�e2����(G��c�0 ���*A�.�x\�o�r{{+���z��{N�!`Ћ�B�0Ʀ�N�xp=k#Z��l� ��0�:g>���v  ��@�$�0N�-�P4��cj8r|�z�ϋ�첒rĮWYm�4��]�,�\�޾�<����#p�` &�<�`g�N���`����������	��ʇlcԅK�~���v�C�l�&f�A&AB?��j%6?��N��vA�VL�Y��!d�J�-W�<�?h�x`M1a�%�"��-pih�w�ɢx����!`t�V:�%e�̝H��6Թ�j{���ψ��R��d\h�/E�+����1�����V��������er�T���^/���)��B��H����>i���	oyP�yt��o�/�]hv ���B���uN6P0 �1��0�zv��t��K�H�~_�n�B)"��Lu�mS�5G&3����#�
�?�0p��B�߾�d����(�s��Ѷ�t>	s��?�~�~_����6�\yޘg�^�߃/��`��\����_� x�s��ڎ�9n�BP�YO�Q��S긠2���n�n)U>)R�\)�5�Q:+;O���л����a��]����<y"�Ph[�WKY\~-��=� ��6`Q�}����~71Y'}����Ҏ���2�C��I��na��e�y�|N�Y�u뼈|3ko[g�lcs���~o��̭K����|�y�� 	��O����I�g��-���9xF�Y��³�
d�Cf��N�_� s��G� ��r�`V�|g�BiG�x�̂{ŧW�3�F�A��	
xWp�"O	�����C�	 BO��L�I=4����lYHX&N�L�ى�c��i��:�u���\gh�@�es�lJ���1�[�Y�~�k�/�*K�cE���'�/tj�7 �8��| 2�g�p��T 
�$�U�۔&��%�ܾ�����n���;�?�2��>�Ѳ06l$�����ɒ�v��0	HȓLi�7�����[��^����x&�h���L׃�
�d��Ӵ��ĭ���p�^�y�Ϧ&+���y�ʌ����KB2.V�w��W_R����)��p2���3�5���3B��_,^&��_�I!�f�%���9#x� A	�k�^�J��z���N����A=y�1�!�us�V�>{f��6����ÿ����o>�U;7�-�0>�^�^���'����k��_��\<~�g�sn�k���O\���1˱˱˟u9 �r,�r,��/����d��P�=<�p��	�Q8���ޘ.�ى��@� ���=!� dhH��/��� ����h��R���̶DVa��a+w>IS��nM��oꃜFn�c=��dq���ǎf�������F.�����J˕���{Y�g� �$�?�Zf�;���'=:z=��j���k�7�#���f���t�|S(�YZT�К��a0W �ӈe�B�
��1��K���FvzHn�3$dV�e-��KA�u$�A���Һ��������q��Cf���{'�)ÿd�T�R@�>��p��?ٛ��k� 1;�zAR=X#��a0	2&��!�� MćH`�؇��
u��ս���U�lv[�a&�G�k9�@rJb��4��9�3Sr&|�̌�x�'?�7�qd�"sLJ�0Tn,����`N����2���k���ϵ;����Jx��3�ˮ5)D]�]`4ϓ��>m��zA�'����&�f��/ID�	�@F}���,�),BY"���`� YB�	�[o��_�e���L�	�M''�Ⱥ��7�g[>�d���g��E?.�2���D�z��A�(>�a�ށ4):��h̨��h^�d���k ��/Nb��Zư�l� ��	J�9`Ay��8co�|dI�s���4��Y�Rz݁�ϴ���Pd@
��.��2���̱$�A��]|�}�\�@�6�{�?���GR�S���U來�:V�z��Uo���Y��83��Li�C�X�+2��4��@��AO��tz�f��X齜�Rg�.� i�;����|���Vg�����1��y5�&�L��/e����@fÙL�����rAzj�&IŘ	��Q&��>[����\>�d<���o�crG��٣���I&�uYK��KB`#f�r��ѣ��.���{�r�ƥ���	�3xX��rZ�\���K��%fC������EO⨑�m).�� '���$��͍�c%Ab׀���? ?��;Y=�B0�)�M�XEd�j�#�	������+���&S�}��+ B���_��G �
�H^Y0�xS�ru�GF��NʏϹ�9���A��Xo|#{���sr~��[�U
�Nl/�9_\r�"(��{W=6GP��6� X
��������B}�� ��0��I�
�5��$��
�����@�j���tD@�}�JY�M6m� �yĔ�? �e�h>fac��B�i��f3��J�NbE�A�?�*	"�l�#�"�ҧ$! Э��&�|�I`�t&�� �h��f��9Swz׼�,�� <�4)�z�n�1tv��0�1e�=���u��F�b�B��4�7����6�LLd�eTc���� <��ц��䠍c�� Ǧu��q]ҏ��=֐ �1��m;�_	��om��"�HڱD����=�| 鐍�̘mM���k<�����zd+��M�Si�T���^�f�2�]�X�����79� �`�B�-���JV�f���)|� �`o=�7ur^؟q<o��0D����/�+�/�u�� �!uNZ��=�Jv0B�6��j�Ӝ�G�ph0b�����|��'2;;��~�#&"a���#�ۿ�[Y-����kY���u"��r���`BB�/�K���ɪžX���Z>��g��_�B��X��X��/��c9�c9�c�Qp�ԂC�˗/e�/��þ����t�//�������a���h��L[-�~aF�=�}�#9?;��r�9�~ԓ��=�X,�Pv�L7�������Q ��А�@��WZ�?���e�5v�ğ���kR�Q�1����k��z�,@&:5�y~:&��C�:��+`V,%�� E�y�Z�W�g�EfB�r
8�O��I-q�P����m��q��>��8�|���8���垚6�/m�[@��@@Y�N#tra���r08�@	�F)�ih#�~1ސi�� a�~(q;�N����b���@��A.��?d�p��F��e�v|w�#���/����%�v&C�,O/aP���c�v�^X&$���9��d�����m!�\6;��g�i�(��S�LȺA;Q�*2�����'�������b��(�K��!�� 	M`�w��:�~���b����j}Pd#h��#���7(CvedٹZ�0�� ��Y
6�fC�2r�0x�ej�4������g�*�-�0p�"MY�D�5�[R�������������D�2�z�O �����6Z-7�,�x���8��@�2���(�;��?���9�/p�� ��`�}�N�ISe�Cb����8�֘^~K�W�K_�`��2�2����̼c����-ۋ���o2)�"�K��2�չ�φ���k��~��8/w�ޭ$�4��@g@�x/U��g���0�9�jX�H6z��
lx������{�X�aL���A�I�l	0���`_x*�_�YR΄@xY=~���"��v0�X�9� dd�-��A�.�J���;�2 i��X}��y/aO�����Y����ʶ�Ʃ�;�����Xn/s�^�9d@鴟�r��_���������k��pY��t��{��c��������T�$�-��v����o��(�Te_�,�D��c�W�S�6w����8�b���=t0��9�ut^�9�����F���������� ���$�{`�=�#�����>ֹ?SV���!י��;�N�kvr.��L�vKٴ0�&�d��)W���1y����n���c0?`�N��(�X\���!����p��;6�dU��蜘�&g���~2�+�{dL���� ��O���1x��Lz0�i��9!�`AV��"ɤ�j�Vs.!(i��t�)�/�h&H�(%+!��ן�2�L�]g�?���E��)
rI���Ijek@�<�� *�۵Ιw4���F�5�`�u�)�$yHc�{�$7��{�#�v�,}��� �1��6[�A�U�3D��X�c��N����\z����Z�|���o���p�I�t�V%<��!��c�"c@3�y�xY���Xk��@F���ګ�\�Ntwe����j�מW8ϩ���kX#�~b�H���7�>����e�,&N�$���� ��?�>)��}��Ϳ��$w���0p�1 %oto�����{���7�D��Z��l�H���\�c�Ґ}��k]�3�!a5�/�E��L��yRA��y��H�G�O>�bz��o�}��h���j���##`�&lm�?��c9�t%��7Wo巟|B�{���C��/�c훨7���(���s��Ʌ<�\�
�� ��z~/�}��7���7�_A�c9�c9���r@��X��X��OW�H� �l��$ru}%��	;H-���rҟ�0t���7_})���)�P�\a��2�x���3������p��P?�1[pE���l[L���޾}-''�zpY`U,���md`B��3�~Y|���M��`#�_���|�p�g`�
�.[1�RlA=HM&'2�HȠ����m� �Ar �w߽��fk�2|�Z(a��;2g����@ @	�#����l�9�	� 4��	>xI@���Kf�L6����<"� ���2���A
4Ԩ���|;�W�-�`���SF7ۭ�n��02,,��rzv�: �ss{Ǻ@ ��Ʈ���o��?h��0�e�3 ��z�}��@�g�(�b�#=O
��;��w����X8�S��2��ivN�;�GH�1+5w��`�%�"�
�]B��] ��%T�r1u���^co��MIv���:������e�MU�QJ�m
)o��%Nv�Of ����0�Ef-2D1�̔V\f�1`0n�O��M�2Ud��\����gXpF�Q�X#;2��A_�C3�ܓ�$6���J����ӓ��y_ެ��^.9VCJ	���1���N6�y�V��{F`>������ ����=�k����t|�)^���6dc�@�N�&0���̣&N��XM#���q�"ȫϻ]��gڎ�\d��ki�NY*x�t%?�5�cf�|Ƞ� h�ޚ��I���v��y��}�fײ����!d�Х����Lb��J��hIU���L���:_�"��H&�Ae7Rd������!��2���c�J��x"�a��E��7�k͈[���jO5�=�Cc��x�O�=� �E�P�0��2�ΰ=�1�ZK�xIЗ�'X���j��|��2�HɾaO�3��k}�4��8��[����w7���=�к8	d`L�՝��L��[���I	2{Z�9���C�E�O��Ǆ>La��ZUr�(��se�H fdK�^����l~ዀF�J>C�l0�h�5|�Ӈ (��}c�,<�<� �`�:��=��8����Q́�7���� c�a�!�s}s/��=��A�蚖��� =�67�!x��������aq_-L�
�V�fd�~܈�P�{�wd�'�vr� �,s���:̚m�w@9@o����\w�W��� ��7��^��e5����xl>]m��ƼC�"��b`�}�>gO�`l���{�X�Ӏ�Y/x� ���&�X�`RX)��Қ �x��2�ހ�F��\^����[�:zl玲H1�8��w�vL��|c6�-�*j�!aĵ|�X�l�}%kG�mA�3<7�d�T|N�]�5k� ��eQ9��>�%�� |u-%�,�^J�q G � L`�	H�|��Reҟ�1���+�Ƀ�X[q`lI }��a�����u�bI �O&���~sx_�%%`�$#��.�ٰ̼;H��/�qM_��{c̘Ʊ/�~��'�6�i��ӈ3�nm:�!��*��X�uBR����¼_FSQ��`mF{�?U:�D�m�{�=t����h1�L�JYr���Ę� ��y�)�ǰ�&����>m�<j�ޣɈ��g p�����K��z�{�-�~Y��n��^���c���R޾y-����B���#��>!p	�W�}O���e��X�{}�!���~.w7�ܧ����_�n?��s���L��X��X��/��c9�c9�c�S�m�Z/��!e DQGmg}_��^����ͧ��=�y�i#�x~q.���"o������\��Q����RB�� g�Dz(���b���^�vT�kl@v`)@VC,�b^��w{٬�q^�}��lv��������:��D�0H�1���p$'���X�̄Ar\)S�q/��`�|��7ZOkf!׃�2$��>��w��!A
(���uHsi��E,�������hU�Z��������n�;��Lڡ%�!���xk�E~��LI#uiY��G!r~vA9
 9�o����D?9��>������5M�lJc�8�	2?��WIK�������P��;�����9�4� h����6N,�<`�ł�53��i\���LXg�� �!�ՐAc 	2�Q����M��`'u�X ��8�`HWi�u+Ek>�w�\�)�s����0p�Q����"�>2}�S�� oZk]F�����<���9y�pcO` �kf�Z7�̯C&���B���|����J�K�'��Ig�;Ue���â�q���������ij�v:��l����)s@SKɪη�W��!<7��"��0�͂��S!q�1	��Qu硒�,�u>�T8J�̋�g�Ώ�$|B+J��dP5��]Ւ����0a���`�әMYŤ����p�����;	C9{t*Mq+��]��I�w���t��k�Wr!�<		$1潭�W����@bO�����F��LB���d���n������䉜�����<�{"�`�u�s_����?��=��~ A� )6,�u�>�s6�IMGI��]c   y�n�d�z�]��E,'1���z+�F�M��Ji�݌evҗ(mu�49���L~���y�b���Sz=�}�?|"�	R�3>�v����d��Ѫ�$������:�W����I�]�r��U��@�%�gO����޽�cc���г|2�Gd/d��>�V�~,c}ﵾ�d-�=P&}�!L�K�Y�Gp���s��C�ژ% �Ƃ��T�����õ~��0�=����}�i����/�Z���������ܤ���`�a��#[�id'���GO���	�(����|<4of�3�9���/d�P�l�Y�@r2y=c� �����BP[�/�F2�y�ڠ�Y���`pn��>���G�� w|�;�j�Ü��cq1_�J�Fc��;HHt��?f3с�2����k�tl.GP�mP#�}�ep�f�E���V\3C2m���
02^����{�� ��9�W-�{0����a^-Ȱ���fx�u��2L�Ǔ1YseQ��k%@�^ �~~׬��xڞӳ�wm��$��	d���^���������$0P����(�i����z�v+�������S� ����h24@A�o���;��s r��>c������Kb���1(=�@�`�7�V��	�:<� �		<&8?�>�'�!�aN�R�{S���\i���4�*���ZR ��X �nvw�c�G�O8��- ƒR��� # Q`�&J`��1J<�����bi_?�8��lb�3�c��w���������q��ݪ�^ј�د�7��}~����g��uy�{ޏ��G\_�x!�����r����ֱUS��}���N~��_s�d#H�����˧���a�~�g�?�c9�c9�c��-G �X��X��X�EHK4U&�������(�W/���o>�\>��7�Z�i֍`!3.�]2۝�`2�r9_	"F_|�kz�����2+�檍LF#=���n~'/_��	:Ua�bB"(�� MO�!$9�c�n�����׃-��҃�@�lR0T&H�d�2�t:���ޗ;^�u1s��	��/߼�O?����-���+������� ,���d�p��C������x�K���F%� ��(���Tf8�j���g��r��v��4��ᴧ�XWC�`��������x���4~���zH�h�j���:?��� �,�7z�E +"[h'�~G�� k�d�Z�q�G����0u���xԋ�9-�!�e  OE�d}d��a�̙��7$S���,֜�I3�>� �B�噽��d:~�~A�G-l3�h=}�X��^_�jy/�g��?��������i^�
�(	})�W���>e� ���Aj`�a�9��p��?�����6|3E휙t�'�*���R�h�FF7ޫ�ό~�
�6 �� ���E�.h�b �w��)IMH��<Ȣ� �6C�:G��0-�*)�7.�@A)iP�
٦A�N�y#�m�}�%K}��P������9��e��kNI�hA�O
�]���N;�ѵ��D����mV�����Y ��3}�>M� �~-�,_���"�=�� J	��@HM� �Q�Q:e���0l���y��3�S�i��RlZ���l���U������g��iݵB�lϵ_nZ�kɖCir_j}��2c�h4(e:�0��6
�7wm30r��_�}%�h!�"���O9���`�$[������.J���X��S� v$c񓑾g)A�c��6	3s��2&�<eD�3�?,�݁:`�x:�� �u�����&�wG�M39��-c�4jd���⮔�^f<;�A�H���㷐8�d|>�G��\�;��jty���p�i��\��y Ӵ���ՙxZ7� >R2�������V�Y6�{p��G�����o���J._����諝?�1x�GC��L����F�r-y}/�G1�wWچ3�uJ��:�u�C�
�ĝ�I���Y�~pp�7��s� �$�T�z͞ջI'Z�s�x�a?����'��3y}y'�7s�+I�cc8sl����W��Ą��KAZi4��3��Jڀ�A�B�s�����?��Cy��3��mϠ�4����� ����[�����˫+� d��	R��?��p�]I܃����X�I�gbn����zH�$~��u��e�ٞ �@n���c�`.���AV���{���m��	s8������c-���%D�}q��ع5�����%�8g (�:�s�ߧ:Wa��u�s��L�bOv�%\<bW���#s�����O~�c9??�z�9��A�Q:����t���՝,u������3H�$(IN������ݓ�I��3HR�0�u�)-Y�&�	c�\�D�'��x�������`�Dd�^_�q�&� ҔZ��bG,�2��i�,	���7���\�� ׇ�CdX�H�}�\���n��R�u<� rX`���$��VrxZ��M�� :�@N��.!�����< "��+�����ك5s�P^�,AGp�%@�!}���W�W��c�NO����ŔW���\���>3<�b�N���_�˱�#&���=����,"��&7�Y��i�  A��Nࡅ},����o��Jkɤ�;c��Ô,쵐C��ozHY�^,w�7�_���O>����`�i�C��:�!�oa��@Nt��������O�I��������	@��tα�G$��X��X��X�|� 9�c9�c9�1e��d2�⯯��buO��������fc{<�!�
�E�m k^�%dp ����}!������0@���\���݋<�"�m0�3p�k���9�<7�sqZ��I�+�!�0���-��`/��I��c���NƔ�b]d�nc���ڳ�;�`���k�4��� �d���	=l3tz8���4�����34����D�������%��8��Fv���1aAbq�-��:f��Y�A��A3�Y��oR)��q�ͦ�Yd�|��Y�XV8����h@����?��~Ͷ��Cl�����º�����#sҁ0������g{�qń� äF�֥�I#�$� �U$�M`���@���e����]0�r������B� �w'�>��Wڶ��dN��V��M���Rf����q�����I�������3�W�	�U�@����2V�YZΗ���ρ�W_<�����}�7C��<@��h]\��v�Oh�wm*���VU!�;3�`�G5,���k�A�0H$�1>99�,�O{ӂ	JE�ø~�/�OPKht����l)H��i��m�����C�y<��ye�$Ґ�`D������
Y�ᘤ�<d�L�������� ���䨝�
+�ܓ��u;� T�=a��;ɢ���YY���9S�I��.�%��������<YS@���h[m�2��-u���z^6���r��d��� �1�[�IF�MF�X!�.�_E�������:/�|�!�m��Ih<�T���~�,<� �&�ҊI���2��w ȃ��������:&��^ҽ�y{��Td6	dv��A_X�8 b@���7}&Ó &'�|���VH�h�_��7�u���z�Vzq#�����e���F�Q�(��-���v����B��ڟ{�t�FR�+�.���d�y�!^G�Q��jސI�џ=dxR3c��X�Q�.o8��;�fK�2��0�+�&
!�p1���j�!a >%�'����v�&�2�YךA�A�G����ɰ/O�k=�P��#99�'P �M�B��l��λ�u./ T ��ɣǏe���t:�������=���z
V�l6"�G���|H���G畲he>_�1�,s[��\�����`��[D?��򓵎W0>�p o���0���!�xd������չ�1���{��@zCK��!zU��)% 1���r�]t�;�N`�+��`�9��,8����ۚd�gki`�A��('�@HO���Px'�3��Fm)M�R�*Fr��=�b��e�T`>�D��	�����f;�$0�z�G��J4���q>��k"��}�o��u.���r���;��D6c�iç6�1;�g��̪Y����^ʤ�zz�?
-p%+�^�L���b������:�/�� `�b�ƫ�l0b��x��u��
���3�%f�w �TmE����)�� s�y��n~3���B!6���{�
90�b�'tR��K}���K�>2o8J�E�I���L��)C�y���#cO��}0�8�t�ίڏ�� �� �v��B����������>�Z�� � �F��L�H�)�C2���1��%�̗s��I�kx�@�u::��s��}z��1�-��' �A6���W��6l @>��O���2��X��X��X��� 9�c9�c9�?Yy��{����am��ɾɶइ Ea2 �I�l���{O�^<�)�C�n�Cٓ'��:�L���n���?�ׯ��ի7����A4�H��SSc;e@��J����~�w������z�e�@�fKd�:�j� 	���F�&�d83P�����眝������p���`�#��C7p�/Ι��cf�����o�e�8=A�Ad�"�C��D%�3!��F����n�����'|��5�(wІ)��"�t䡼�(�Ք�y'�w�R �J,;9,��6��67JzH�ԑ7Ss_R$L�;��4��	�ϟ=�Av���z�#��\�xhFഫ!�䓝@�ԏ˺��(*�*~�3���Zf����'�Yx���B��lSdL��Ҙֶw�sp��0��6o�P��)0W24�5����p@���U輏��1ߏ��/�m.u��Wi߇��9UI�B��_�5�"��t�ǂ�cdD�� ���0�T9*xYx��
�_Jd`JJ[w�/w���I� X*����idr`A��.�	�P����	@bO�[N��2.̈��U@sg�U�*ږ��bJ�@�+�_����:�>���SJՌt\���$[B��ׇ��g��~d���u~��AO��!c	�Y��.����A�0�t�B����M�M�'��FEΤ�"}��@r��97�׊��l�a����5�GP4F�@�=��?2��a�B0�ka��8}�r$���$�:T��d�``6\�_s����/��3��!R �\�Uq���{0�f@��f���賷�<~�J0�:!�	�2H�W���:{����}&% �h&��T� >5`�xfJ���h�+��c�-(UES��I�y���:����#��-�����ӹ�W�\�uٶ�~*ul��z1}K�E�ǻu#ח�,�	��E,��B��?�g��^.e����'6Gro���￑��h_�����Vb���~�e�,L��Z���`8���D��ÇQ�C��\*�����@�{]���F�<0�D�1IF�Yg�!;{R˓�'zMd��;��H���^���J�Um]�e��P��#dǵ�s�o��8G&Ke��m�;Sf�¢�X8q�����p��Db���֗���$����%�d�����KJ(A�I4tO�u�96n�ߕ��@��Ln	uY���S�)d0���r�5�Sڱ���+�|����7����u���F��ڌ~�2�����T�.��z�s�*~�*#GLnІ˝�)�ڂ����`&@aR[Nǜ�^�s�Xױ5��5���zA��P�<@Z'w����G ������s�+�0b�g ٙ�dr&��X6:���?M֜Ѧ�]�� �0������d�@�A�Z'o��
鳑�׾؞�X�!I����q���:��K((��s�(2�!mCx��H(�#qc�@��$N��e������`�$��E��No�I�WC��s�o������ޜ3I7s�f�� ��{M�G6Xk��f㉜��t)�d���j�{2������ft.�Yȏ�Az��&�%dQ��|�nc�u&�&��,\���0F�WKy�Lɟ>{Ƥ��?���*J�.��t� �X���!ĤJ;1o����2i�`��O)W�ɦ�,�틽��鄦�_�����_���I��B ���霈Ӈ�c���	ٸG{ ���I�ӓ���d6����9�>�\���`k�5��9W�-'`�����g��?t.]��H~��/�r,�r,��Q� ȱ˱˱�Ih�cdoBz���kֳ�TV?��O䧿�9�䞟?���s����s�<yB� ���^8�|��O����O��a
�:q��h���^��>�K+o޾���``r��F��3$��ѥ�PS�"�	Z����x��dl�8(z`�q4��b4$����p�8bF��`@�����?�;|��7�Z�h���05stj4�,9 �:E��pxfv�"���f:?�7����(�/Č�f�2W�R�{C�Iq��(4��ᜁ� 5�a|�:��?( H ?QU���C'���˙���8�s��18�$�1�!�����Gd\_��W_}I ���ւG̀GL�6�#�E��������N��3^�)q2n�2 *�.��)����L�ρ��*	����` �;�|���%��|�L��j!{�9�И�u�B�>�T�O��10�X�_��aV���/�ݎ���l�F�'=w�DEy�G%@�r]�F<�M�=K߂�<0;�G��mЇ�IB�E8&��KcL�[Hy't��bX��� ��E4'G�o�,H� �Y�x�0p�Bߒ �s�����Wii�As�e��20��W|I��b pb�[���~(��Z-(�,��}f�|` gF����>�<
Y(A��U�4�!���R��7�{3^��"�`��K;��{��MN$�����!����MA�5�����_))b�4!p��� �L�v�L\v2����@.�Uߧ)w��EO�Y�{��/�Е�w_����M#�$�&���J��SY.����,֯����I-���=��Y�m��fy�χ�b缮��`*D�D�g���G��%M�#��m�H�������x��Wg�gQ@q&6�9����:�Y�����]f&A��^��]�$E?�7���ݛX�}+�E#����7$��( ErR�X&��$:I�}!��'���KbIz1�#��;�֙�u��`.�����)�2�4r��_����e��`���0��\�fa�_+�۵�?�O�yf��X-6�����{O���s�e8�v�K�nd�n$�>�_�K*h��8f$8s饤�����TZ�D���VZ�2&�<A0~���#��`R � ��Ha�M`�-YD��n�dZ�˕���s�Ef�Cj)�$/L�$�0N��Iɝ>�.`>�u�W9�;J�XƜ�1�u��>'�SJ
�c(�E�"��ɣG���L�c&@j�V��L~� %�	h��;�� 	���]� Uո��LB�������}���S�ws�>���6����E�  ��@D���\"�\!! o��?����`���3�_�e�c����_�x��c��՗_s-ž2����;`��OxzẨ�V�>��@$�d��d�	#׆D �l��s�<���<G�=�k�>���\���y��������0�v-�)�� ��a�����d$��-K @� �1! <&�=�1�4'�`Ա�k¤���\����|�|�)� x^�k➭���{�p�T��=!�W���3�~�{�;0/7�@��:��W���|��!�Q�>���sn��TZw�ހ$(�8Y0��1iÈ�D��3�`WT�;���tµ�}χ:���:&�>�h���յ⫯~'���_q�C��ru��Xa��犸�E�v+�/��x��s����N>�я��ޗ�l�Ĥ8MLF�?e�������v�A�n=_���������[c��1˱˱˱���# r,�r,�r,����C������L��?�@�ݿ���_����n���[�SY&��cMj�����s�>��cy���p$���W���i��L��-$��(5�[���F^|�Bƣ�|��G���i�����f���3C����@���i�� 4�<��Hzz��6�0=p��y�ǳ�%�8�^��3+��o��_����}��l�sː��HD.��>�`���0Ns��䴐�6����g����W; b�3��L��F���8�d��Xd�tl��wM��t��:� :�˸3j�wٍNz����X�Npmʅ@�`2��Ȣ(J�z0N��ӧO�O�v&��X�d��Z<I�e���R`rM��		eBjF��c���H�] ��v�w8".�`丐�� ��'�~��㿙��i�3���T���,��|����*o(� #Wlx~���}'&� =�����t���#crd��j ����7�� ��g��A��=�F�:�[f7*	��s&���;#{8����� ���ā<��{�� ��w��X(�4�'��K��rMe� � ����(�[f�z&�BfE�@%ҏ!��`�n�cqw/�����A�Z�W�� EAS��Ź�#�WhB�AL#Կ#�E0��ϡr&á�3�Dh�1�^Ǣ�-�B��➬��p�|<K� ��c��ak@p�FB9#�'�vY�������Oi9��T"�	�|Ȳ�s/�-*2��>���q�j-r����k��>�Y�T&�J��}�u��O�߿ж�h�d����C�� ���5�4���Y�D=�����CV�k�mW��1��B�8���]�UI�xrrW���kq����!&a����l�}3�-X@[G^C?��m)�+�˝%w�?��1� �Q_��{:��<0�O$�A�p����Z�Ė�U&�ץ��U }����x��>�}�������)���hkAO�� �n'q����eQ�-��v}+3P�k���#�xE}�r�d�!��)(0l��r@:��C9����<�m����\N�Ѧ�fڕ�T� ���S�����4��5��d ��0���j������k����-���6�(WuN^�w����4 =t�:=����w�#��qY�6�1�}&��<z��{��ٔ�2�������wHx0#��Y�^8�{F�D�u�g�s�y{:v��  ���G!��k�I�������s:��~ &@_
��!���I���-bҖ��z�<�!�w��H�L&�$�i��!���ՙ�x$�f�5{����o�׾����{ε&�%6�u%�B � �������W���@�
����~�֒�����O�E`M8�2�Ǖ��C]R.
I1�M�w/�n�ի7�ŗ_J^�Ƅ�9y��[p��݁yP��� ��RcT7-���k嶀LV၂��d�W�b �L��,A�|-W+&o`��>=���$$؅ڷ�&-]�:�دV1���{��"{�Q�frr�Wx$?<�Q��

��b� ��2��p\��dH� [t�%�x5]�\���w�O�j�.{���=k֔��4�o� 20_��V~�٧��7_����l��� c���:H@��+��������j׋��?����+�o����dQ��U蘝�$� ���qƱEY��dP�5��'�����>���c9�c9�c��)G �X��X��X�d��m��'2 ,�p8N�G�D��?������C�)�8�.A�.+d�` ���q��xF���������L���������;o߼����pX �SR���Ȍ���o�*��O�p�c���o�x�͍,Sj]܀�gl�K�L>�e�#8�d�)M�d�Ȣ�\Fÿè�����ɩ>���/�|�+��g����&�/�'���Q���4�!��7HU��i���w�@�3x�o'kՙ<��^��U�&�Y25kd����~���e1�w����e1��[@�Nv��6�y7�J2=���l�4a6�>�lC�����)���[y���l�;�W@��^0>�^�ߛ�2���:�)V�a�D�{zvB0�߯k>3�D�����������k���A�"��J	�B{dY)�Ȁ��>�(1����T%�i����H]�?C2��Z�Ȁ�ʖ�S����B@R8-�V H�-&G㤤��eo�R��q�Le�� ������-�mÞ�ϵ.]:�L���,yǬS���,,�:ٱ�$��h\ �f�/�d�BFɔ�Bvy�\��A��i�뤴<amQ�ï���{�g\28��V��w#����8���J��R*
����.������ ��/��{���e�xV8C�211=I�]��f����l�zy����LƉ0�(��)^���@A`�2R>����������C`>A%a�FpL��f���m&WoIJ�@��$?���U1��43���.���O	��$	�P��D�&Y�Ky�Zd�]��[@8`2=�S���\M54�1Sm��U��	��`d��;�	 H�����G�V��٣N#���.�mo�����1��I��5��@t�T�wC�!��2�M"|rLl�ؼ_�ϝPr��*�o��1���#���͵�{:�JO�} �����7��ҮM��}a���d��|X�p˩^�ݷr��ln��h�MZʍ�9���I�������ҙޒ1i��Uf��IA�r ���b��?b�0���<�����n���EÛEG!��0��Gb ��aOP`��SB{q>�dG��ID��#�:e��2�Z��9 �>ۓ�����	Mշd���u�Ř��kn�,�2�з����d4弉�	��5�F�?"m���p���oA���6������3� ���?4)!�U1<���{Ϟ���9р���O��#�=����I���:�y�dC�	5�*�͊���e0����I������_��>���b��ۭ�~���(`� ��)��P��� /
mx7�_��a㼡��z�!0F �I�-��ga}��^;8�mK/'>���{]�s�T��n�l�{JS�cퟱ�q!mf ~��?�\Um~{$* ��'dd�d;c���9"�c�I���Пun�\�}���ݘ��ׂ��ٙI���?�ޫ׶���+�N��nSQ�$�-��n���b��a����_�[?6�@���d5�L�"Yd�������s���>�(����N��^�[���s�'��V/@����ɔL��.w`��>�w��o5��';�$~{�.�FH�a/�MzJ�Y�K��b�e(�
�0o����a��Q�G�:���6��?�6��Kx�x���P�Hc��G������?�9�KN�d�������ȤF�&�9��3p�,�k?�>��wߑ���[����ѣ�	t`� �/&V�LA��`@����,�l���g"�~�2��O�O��2�e_�e_�e_�8� ٗ}ٗ}ٗ�[��w�J~��Ju�F@t4<�o�{����KL,���i���w�Bh�ϘQ��%���U���t*�z��[<l~����ų/$�6z�M�C6�pb��V��q ��N�wޡ��b����k����̰sM��x� ��l=JZ��e1*���!ݷ�J���� 2 �V����?�v��Ϩ�R���P���Qd�f��6��$��6�br�q��͛����(P�7B�w�R�'�S$����3��{z8 {���������sHE�甋���SE�,Н;�]���:����B� >%�j~#{������p _��{lG�8�..���9��'X:+a#�f&і�kH+�(�B��zQ�f�"H���`�Ϛ,�
�.%�w��i+���\�z�~��ip���"Y����2,kߢ\��ۿԾ�sxd���8`(���	����Ǿ�����6B���H^^���11<��x*���f��^ J��,;3�Q喕�J+��2�XiM��Z���oRK��j1Y�����׻̤�hbk^�,�OEG�+MZcaL U�"���l���X�����72������C�㠨ֆr�.�)�|�,�o9^X�o�I-A�F�^Ei��Rƌ�5f��sq7Co��h�^[&~��,�<���/�ّ6l����}����-tC�l� ��?�<�L&z�~��?�2�-����d7��!8�9B�e��ͅ�re�7�02�m�Ӡw{d�K�I^�8l+�h=/![I����Z���֧�v�"ɴ/C��|'J�1���I����X�/�N�z�$��h�m�Aw��abF?Ǉ�wZ�J�d%u��,�І4���C��0���F�J%mG�m���������I$��/�c@H����(Y��JƧ�L�:���Y�k��ã����D�_>���J��'�~�wd4�A�L�a�E_�<��֧C�V����^��	�@����]HwP��P
ϘN�2�<��@,����scm�F 3[O��j�7`��3�pǟ\�N*7�#�&��K{+��gAW'i�\��R�#��?%�k������������A��	]?!�9�1�9IIG_�ԡ�G��)}+�o8�@���ͫ�h� �������z��u.O	�)���e�^��זu���|!��LvR�eB�d�A�g��9Xzߨ�t/��  Y�V��Q�7�n �'�4'�>`|O�a�\�mH���� �.o�dxeF�}]���\Ĺ���۹\�:��4��1e� R�F�7��д����k��=D��j�3x����'���� $� �����Z�4]��X�񚭩8�m0�h���l(��VV�TV�[��r�G�2���Q�_Is�B`{A��"א<����L~���,:lN�Q�y�c`��}��~e���W�V�	��U[qrc���ñZ��@z�vw:� �ܗ~$����C&8�=K[1ט[Y�M�ؤ�;}����Y2�բl�;�>��=0��j���g����	Ҁ���Z0�֛��&��uɄ�a�� O/$��g |�?H�A?�N|� ���	�c:�3��d�̗y����'?�_�������Ü���=��x����S &��0F�ۘ��Ƀ3��������J�����Oֺ�!��t.X3�c+K���vDXDBrml��c��km�����������/��/��/<e��˾�˾�˿��C�`8�G�����)��6�x󊙙�A7�����Ee&Aq�=~�c��G֚���d�L�z@�����8�Pt���E������4[��w~�Z��j��}���[z .hh�Z-����f��tN!���yȀNG�};�fi+�JX �#=�R�#O���X���?�1� 2*i�)�'M���t������43u͇�Ff �ڮ\�.���V^<{IAAہ��e��^8lC���8�iA��.��p��1!�d�	(y���ֈ��!�2���X��E���^�� RgY�p����u� 8���S����-��M�F�n��Ӭ��H<[����9ωXG�|�a���m{�0�\m`�@�B�� /p��Lq��O-�����,3%l!�#`��<2 ,���� ��K��C�1�w��redY ����'r-08L�
M���dP��d��`�1�0I*ˮvpخ�Wf�L��d��՚j��y��%�#{ܳ����I�w0�;*�k];�ޣ��k>�Mo�%�Yڨ���~)��c}.��{�OiY��1mW�k�$Af�o����K3�+�+O)K������y̜Vc��� ��m��X[���]}���J�1��re�%՝�>*ԫ!x�IB6��{��x�}�#XL����A�f�"��!)�JA��+	Oh�w��>�>Õ�Y#�6^�@BSsb��v}J��c7������$�1����Dt~x]_�^�% ���`!P1��]�5�hy":�I����;[�! �a�܈em��1�FS�澭�� l�&#���&�T����u��K�% A����i�L�ɚY��>�3�u���4�8]��J��2$ \���dy%W���������|�y�UEێ�G��b���5
~7`LL�	�V�jgV^2���c���ϟ˫�7:�t.�� ς�E�������m͋�=L�7��G_�����lS��'}��w�����-�PIw�������m�Զ��WK�r
���1�	������d+�(;�)"1?#�9<��u~���r����@:��2�n�� JO�2�Qg��O82�Rjg<�R�s.��j�"�
6&�m�����L&�C�]�Ԣ�5y1_��Օ\^��?yK�����${M�^�Ud�qm�KG�%ձ
�	��4�^?��sL�g; �sx�(D�����l@M�%AyO����e4�<�d�(�2u�X26�Q��J� ������i�W��e<c`������3���c|�k!��o�� Ոv��;�1 (`1�oMט�����X+.�8 �Y6�P|����e)��F���u��JK"�>����_���!�(��tB���?�ɑ4��b���L=�
�f ����i�@V	�a|dEL�[W�ؾx��N,Aĥ'���n������x��-X�2@(Y؂�b�Φ(8G�w�U��Q�L�[�|�
�y�����p9���&]P��2�{��U�N���J"s%� [f�C.@�$��$x̀��\&
�By��7�$��yI���;�H�@_[j3�l?��?2fs�{"�(��z�a����8q	l��%���T��o>����'rq�F�:N"���m��ﻔ����t�v�
IJ�>'ƚ�ա��w�}O>����aBb��������V��Y����R�`�f���7�� /��;�1��?��>`BB
w��h����o�����ɾ�˾�˾��= �/��/��/����w������B�?��@���nE��7���o��g4)_�����KY���顴��4��ñ�^>���sy��;���~WQ]�ݖ�(��d��Wz ;yx*��OC^�}��9��a��W��'9u.��ߗo~�$�����ϭ��V�F���/���@B=�<����8(C�
Y�`JD���O#�lX>�����~��}�-\�~��Bǒ��dR4�D�H������S&�����x������q���&�^�t�(�t<�!�P(�=�q��,��=>#ACW!���Ԟɡ�9�\4t#�0%�HC������p\3��F�ed6�:�����!3u����o�����������,ެ=Y�����(�� �kJ�!ӱO3��jɠ��;�l�����P�b ��Y�Ƞ_��D�Ec�=1�����Ff�e��I.�8g[�Z� 8�C0�C�"���E��bn�����@��1ٚ�҇:�wُ����sh�R��"~�n5�G�_� f^I��(���ɷ���G�&�җG_��wRQi+�U��#�$xrT�`�i�ޏ^#F� ����9���1�L�~�ܮg�$Ǫj&iw����[`��i80���Z���~�~��)�C��K�
�����}��|Y*{o��A�rL!� e�g&;�B��.�A�Q����@k!�0�~��k��ʞ�;�����F�"q�>�u���� K l�N�ҋ!@�ϴײx��=����{"/��~�Mon���L��%2�e���O�Y�}���pנ"\K��K���S������C�/�:$�����S���&4�w����_Q�N��>7�X:��`̑������i�� ��0eV4Y7н��N����������K�w�r��v��@NM�
�̽�ed ���k��u.��y��$�Dt�j	_��1�f)��J��n��s�	��xR���v��:�K +֐BS��hz%S�����ƞB�V�d�c<��A� X�cd4�� [W��J�?5W������:�M>,<zs�쪉����(�I	�4YR�V$�1(M֤�-���b *���!x"5-(�����9���1���I�+@>���C�GdQ��6Lj]S��cH%P)�x������������i?�ծȣ�qͿ8��N��:�:b��o�k���~��e|x,'�Grxt�v;<:�g:�/��\�Y�a�h�d�� �e0'��C�+�p��� }��b����_ʣ�oɠߓ��]�I`�������b�N���T��Ԁ6]����G�$+}�&�a�dȽ1��� �t�c�� ���O�~�׽F:���)��90�#�~�X��8' ��Go�C�c<���~�`�B)9Ǥ� �ԅ�U_�:]?{Z?�G��M�`%��l�Ԗ:�a|�9	l��y{5���,3��L�K�u�^�����`���r]���';SQ�����--zF����Z�Z����*"Ѣq(�cx��S�"^i��L�u8|i��n%�6� ���A`�i��[,��B����j��QI��� ��wtru}��:�c��t,�1�+���/M�<���!;�" ?�w�� ��"|O&������a����%��������j�%�d#Ϸ���7L AA_8:9W���t4��x�{�H��&rt8�gа���� h;2��P�= ɧ/�����=���Sy��^scҰ�F��v*��{¨�_h�`Wb:Խ�K�����' �q�$�$+�@s;[�g�)?������O��5'�g�vC�"����/��<@����>��n�$�������G������˾�˾�a�= �/��/��/��B�H=� �1����z �������W�����p���,on��F,��t�У�D_���Z��R�����3�� 	}�P?g�l����a/���VA7���z�M��Q�ɘ����cO����?���kO��8���#�~��.�>�|+ ?Z7��^]�=4^�_�g�}B�s�5�c�Z���$ �C�����6o����qhz�k24�e^�f��YȂ�D���=H6r�|ɀ3���vh��ڤ��vަ4�L�dդBr���Z@$h�,xV�p�V.��eʚy�ךFSB�����������<2�=���^��/���r�h��z��7�Ӓ�U=`۬c=S�Ǔal́�لn�a���,/�'�1s�@H�i��^�ݍ�X, Ĥ��ߚ|o�7�d���VӖ�P{���`G���t�NE˶H!DI(��#�	و�ޙ�i�v���l�ͳ�j�f�3#��`p���@T�_���m�����/����#��R{x��Jv ��uQ��D�~����Ĩvݙ�I��:ð�I�-C��fh�U�2_j���������Ӽ���pI`��I�U�
�
h"�Uɬ��Y?v/m۲G\�|�:�Y�P�:tё�-�c|�=�C7�pJA�	��i6���W�`6�40f��ԡw��p�ٷ�><2����N��p��fK/B����J�{)G�L�33�J��L�dn��+:ޑY��wE'Q~����������a(��+�����H�m�Y�d��v3 ��1����xh�Ef�#��ҁA�
H�JI��t�|�A��@
��1�f�]e:WTmx��o S��EFB�_��L@�	t��� s��<{�L`�ٞ���g�i�yE���y)��\_�$t@����3���)7�����'r~SI�Y���%��S��d��C��R �ƞ,���11��?�0(���Q �>��]���M"Ϙ��5�h��5�"#3_��f��Z�ݝ�͞��ӹY�d��V1k��S�,�[�;�۔���j��S���u��I�h]'����)J9�еY�M�sB �[�_���[�k�ۡ�Y]9&å%��7��Q��6�����&(	�L�̘a/_���N�k~��[���` �dz�$d�ט�RF�f����X+`�҅))�͈�ӷ���W����uڑ\Y�y�l(C���&
�'C�]L��v̴���D�}�k���ZvA&1i��Y����.X#��UuA�O��Ȗ���I��.�o�FS��R`=|�����`�}��懈 ��>�=Ȏ 0	đ�p`~YҮ�B������ Qdߙ�{W�.�5����L8&e��V���q��_�(���@*�t�,&����X�Xs�)��]��Z�/zth?vkcty���h.�x�P?_�j]��&���wk#$�D���v��3�2��WEو��5<�
3��=�_^��� �4��d���*��|�\�C�,A�I' �����)���bE�;2(��}RY�<]s�#��!a��F� Ra��x��E�2�.@I���O]� 8lA�w�m�d���a��=db��X �
~'��I��qN�N��hS�deb?�r/��u�&�	 �-��$�I"^���>�<<��������?�L��gZ�� /�>�9e>�P�9�+��"�ޠKFIW��#曶/��/��/<e��˾�˾�����h~�0RLEa>��o�Z�e�����#�� ��@ԃmZ���&����L�<|D �(3p �	 �j=��z�,JǷ�+�8���_ �W�~9X�M:88���X��g8z�\K�Ӆ
��'��/>�y���c����P��_�J?wA�b���=�f����rzz�@��l&��BV��ᠦ����`�Pt���g���6�Rv%���3}���rxx(�A��TE,p��u� ���R�;�RB��O�@d��&�O�,���,E�(�ρ$h�\�u0�[�	4(o�z��yb@���92T�*��D����#98� �}<��т���r�\1(mq�QI��Ƞ�}D tC0��҇T5�=pOZ�y���u��������w
���j %b�*�-
���Z��(Gk����r���awe�?vߣ�+��U&}����[����6p���,��l��I['���4a\�>7Xb��j�������N�^�����Ju͸m �%_�j ���?��ˊ��}A��?+eiF�Ub T.w�Ů�id�����s���y�;����a��w �-����@������`8����\��NֿyKI����NU�f ���<��Z���#nݦ����� =s�>䅺�� �ߓ�=gg��'N쁍x����]��e�����d�J�0���q
	��B�qCPD'`�z�F�W1�$!{���E��c��ͬb�8G��:����k�"n� ��6�����('s���_y��X�z,e��:�M�a�ؘ�����@���ה+KW�y.Wb�Q.�\��3F������D�hr����<���X�Ǔ�yp���Kq����J.o���ٌ~ӡH���#����2
q��[�B?vi�h"r|p���XA�y`��{~�"S
TaO׍���?��(�X���N�Q�T��+��S���ept(�x�����S��X.�C?VG�t��M��3����-YeAP@J�bg4�j#����n�x�Nb������� 
zrr�H���r|��� �	�0J�� ِY�L��� �H׽�� .Y`C�x�`rȹ�6����u*�7�@f9d�p0:p��z !\A�����`{4u;oU6�1�Bh��L�B'�;ҵ���TF�N����lt�lb)��,�W����<<�H�7��o=��ob�B^��7D,}�`� ���Ǳcj<�H�������H�SYa�j;����Z�X�:+���X�S&��Jo0�>�7����D��F��!P����G@s�*��{�z�Hѐ����$1ݘ�*E�@�=˶��Vը$ �uY뾦��Q��(dbNF�k�f��}���b��=�n�lл���	 yO$k`/��$Y����G�5�L��n's��'m�66��#ec����)�k;m�M �?�����4��U�G B��ڤ0���Z+�6��b����4�F���iv�S�v-�^����l���l�#��0��~-�B�s������r����Ԃ̪α�IKH�#�՚�����8�d�=�R��)D{=�� =�\ ��Z�c�n�  �ƒn<�C�����̄e��6k�h�9��d��u��,���q���/�k�^ɷ����6;�?� ��6,�}ٗ}ٗ}��.{ d_�e_�e_���S�E��2��=�B���~�@"<Ҥ=h�I斔�*�8����Bp��K���s�l�%3��a�Dvi����y�B�s+�I�ח�bE���K��V4?:2`�����wu}+?��/���@��
����?��ƨ8��w����dO�~H��U�7v0n��p�0�ԃв�	yE f���z��	-h�Sp�[.7������a�����6���F��q�Y�wW��[l^< C�	��z�;F� 5���m�_�@)�$�A�F�-��:4LG�1���܏�s�%��K��k�_�f��H��[�D�g~p�~����ϟɋ7��j=Jp�8�òߘ4�"u�`5>H-h����[	��p���V�c������H*i�dnm��֭�-n��B���ۢ��Hk~�Z ��o@�k��GF� A��������e���9v�o5�[�
�Ȱ��g��������IqU;��a\fk��;Rp �An*�"�]x+�E6�6XC��C��?��Ծ��Ʈ����Ҽ�{���;Х�,���Џ�'�S���
r�{J���w�5R�O��ޓ��]G
�c�ХO��!P��7�4�H	��7�*Ң��B_K��P2���v�j�D�zxd'A.�q��N:�����J#k\�I����'rP�E�+z��o��3��P
&��鵒z��7:�^|q)ٲ�A��D)�k9?��Gz�nJ����� �f�_���O�u�A]7��������u�a�����\�|z��$�E̯��4�`���G)�B1���
M{'ӡĩ'�,ֹ�P�#��P�ʋ�F����t�p<�㣱�n+��o��v)�_�r}#rzt*'N��+Y,3٤ښ���l`�4G�.}<ь���TƓS��C�G��s�����M��;�w�h�Xל�>#pvBo<��:�7���X�~����s��g(@�H�-���0��f%�"�܃��X�l*Y5��s��J�x�}g.U�4cjL���Ȓn�hpw^�	�u�x���6؏X ���.���N�y_��	�`̅&�&�狁��Ø
��aԍ�U$��&�7h}��X�k��}7�P�c�"�T��_���#}�����5�h�\����i+!�������_4�7�	0Hj�K&8�	��k�O1}6|�[#zb��xt S� ��~TS��uL�R?�����J(u��~��v���М���0�^co�0�{^��1z5t�m���w�k���@�,�����IIvm��4Z�%�z#��2]��{��ؚ�1h� �E`��Ҙ&#�kU[�BP����W �'�@�� �@���6���B��8-�T�?�Ҏ"m����Nc`�n� �A��I"�k��m~  L(�'&{I�m;ԧv�!�kf���r��F��n�Eɶ���=OѶ�1d�2�G<DЏ ��� �[Vw��5,	c�:L��٧Um� �w�[����~�{z��:��]�jǒ���3����'k�-�� >9�s��<Y���c�[�=��s���,����=��=d��#�}��ٵ�Q~�}�� KU�^!�&��}; �v�@��ca�G��ч� �k`�[�l6����Lu��$��޽=;�˾�˾�q�= �/��/��/���ˬ�N3�R���A�  �E8��4Ճ?�Do�odQܚ�(��vC@D���Nˌ�����1�c�&��kA�����iZ�\r�ހT�j5g�q���{o����G�~.���$�<f]����d|.>�C;=f7��Ry��^���Ӊ���{��G��P~�_��2�u����2�ZɁP�$��o�3�F��̐q�a����1f��ƨ�h��tJ�!wz=��'��q��e0�pi�D���M�H�8�R���7�Ѓ{����pCW��C� 	�;��z]�I�_Ֆ�G3RD5>G���uuJ�Y�6�z2Zj��Zn��^�1	����$�����rc�	w�nWr};#A"\�@@m�Zv�n��!'��mY�	�48���N�H�/�|.m; @b/6rZ�Dt��W�����P�� �o);y�DrF�h1	\�pp��uQ��z�I��OƖ�a����;٩�2��A��{(����=4 ��{�_q���T	��Ԣ W���D̺���]�C�{,˄�g�&�d�����N�jz�׬/�d����e�kO��o�#��yu��W��c6ḥ�W�e�"�g�l�ʛ��W�c���S��.=?�U3�MH� l�)Bcv>f�d���jz�ܙg�E��qZ���s�P燂�xQ�:K����P�}��Z��#�^�r�Z6�s}f�����*�}5�t�j�?�k��0�^��C�,x{<u>�e0�:�=���j��jUG�"�߲��Fu���˂X	B���D|mU��_���%�e���tcٔ�tc�̉ ����ܣO��U�Nx,��X��#��߭��w�G�\�h�S�yx�i�;:}�<_�d�y�_"��F�7���T��;�;x,�_&7z�K�!{\+|'������~�/*���D��#}ա�z��M%��T��K��MZ�ͭ>'�#z�H � ڵ�����c�����=BD����^ �̇<a��^>���H�.(�H�2j������$�oū�V~��lG�����Z4�J4B��z�xY�����{cq�S&���c���`oVd���s����$��\����~�q�`��x����>}���Nbn���O	�� �A�`2��dL`�@��&"�=�S�#[�k����E�'�� �M��IjR�`9�i�	̖�У�*�=�t���C}�T��$�)=���2���V��8^1����Qj��)|3���p�տy4����� �� dރ=��A��p8&3������	�G!k��P���!����5 +�|��;�tԎI2	 k7���O����d�,�_I�\��"�(�h������rc�B���	�v���i�ֽ�vMˠ�K0om�3Hʒ2\���2�  �y�{�Oឋ�D��a�B��l��yv�U�+@7^m�:G >G������	 x�8&_��%�����j�K��蛔A�L�,M8~|��M�p�*u��Vk d@�x$OT|Ζ$P�;+���1H�U�R�$�,�3Y�����nɇ<\�ق��L�#�I$��`A ��|����6���i����{o$]���Z�s���&�`��G�����L<O�Oџ�����<hi-�g|�D�ǡ�	&�!Ye����vq��&$'�ݻ/��/��/�e��˾�˾��ￔ��|�L��Τ�)ZɡT�C=�F>3�N�d��²�k˨�F��8�#a���!�H������H&e�Pv�r�fD�Wv �$ �����<x�H��=f�~�ٗ�ZV������,7<������
d���oɟ���˻��C'4��?&'G�����f�0TŁs4�R�I~��X�J��0���y��l9�7��b&ue��=��k��y�L������z-��ev�%��{z��h��38HZ��7���� <	P�~o(��w�ƞ�A� LU�!��ݲ|z����E�Q��p�����ek���WA����������#N0��� 6���|^�]P�D��=�J������4XE��>�R�x Lز�K�/���Q܊���|H�Ȁ%��mYb�� bl�Ƿׯ�-T`A;��[�af�Ia�Kd��e6Vm`JJ�@!&Ӵ{���l�20����⾟�^bܓ��kd+��^(�^������n^ ��x�w�Д��Pb�Q[�)��Ly;lck����ײ��W��ø�ߓ{�҂%yjuK��[]�d�v�I���>��		[i+��a�;�7�����)���@�����@�UO2�L�Ah��qTi�Ap�(����𨽢�)2�\�BU�Xf��������#�^��N����u�'���!�¥^�����-�&�9�P�:���3���>���f�vo��dگ7��s��]L;>�Hoz$��>o�	������u>Ѷn����z!E� Mjr	���6�K48������-�#X�ZVI,A	F
fP_��o^1`"o^Υ�;r��L��R:Y�C��H���uox�s���H�b�י��^�s^4���cIu�_�,6��J���,W��6�D�W/ӹf1�tq�m\K���P��@���ܓa��gr���J<}>U|+O_��g_\���7��m�B�I���y�tG2N��t\N���S"�v�p��CbmP��'2����\�b��H�z�s���E�ɟ��+ 5��_�O�X��|����g�l��xhh��|��������_D&=/Z��)�O��-�˝�O)�0� .�4�
b��rz*���� >
0?����XbE6���P2R߯}~;` DD 4�� [s���`M`|>~�kB�ϸ���<f]�@����c#�>!�)�Y��g짮S��i��>�$�
o靟�km��]$,l������X�������� `��r���^�L�!�d�J��O�^?�l�P�����)�"��8-�&�`�p�p*�&�YG:�,�|�d��c��D���$+5j���e�l�@H����G ���c@z�Li]��h�N�r�|��Tm�x���:���Q��tm!���	%H�� Ё�f��Nz��s۬7�Gׯ"й75���?�����GS����1�н빤u4�ɹW &a/��q�����ײ=�W�e� ��z� 0�� �2>���d>ߢ����5��ң_SG�g�6�"h��X�s��&�� ���1cn֮yx��`�6��Jf�_�� ʑ}�Ml C�e΀�;[o/�{Y�5�s[Ф&�EZV�0���91N��ʩ��W�Ӳ�s^F	-�f�;o�8`9���;Lf:99�4 ������˾�˾��G� ��/��/�� [vq{˃�f��ᩩ�� ���zؙ/���D��KY.�2_-i�X kOO'�����<y�]����/ggg�L��� �H��N�G�`k��V�#S��u+�@ Au��i���^��"/e�\�;<&e��xz o���|�{ߓ�|�;2���O>��>��,f7�����i,k}�r1���4(�B?�4	,��f nq�m�S���#�ģ/���R�]��zHO���@ 2�OZ�q�5�H"@�G�][ű$iBp	���^�a��fPc�1s悒��X�L
�f�y|�U[�8��
�`bP��Ʊ�|߻�5r^��b����k��r#G����q?bA����%k��=ޗo�i�`�IS�����Q�}�Mj��  �� ��~��o,	;�3��5���.f+[�M��"��{Ɣ��V��I��.���Ο����ɱͮ��x_>�s;}A�`����E�׺�lV����km��{�۾ɲR[�)�A�¶C %0mx�N�k[�m]���V!�>*9A�~~O��kA������(]d ��\#�SPv-8����@�-dݚ��d���ym��."�}�w�d����Ĥ-��A��)o��V�ʲ��֎���F�u�U_n���rP��Hǯ+~l #ڸ�c�|���m����?ѱ�ǥt3m��/n�1��:_u���R��\�di}��C}\�DCH�����1��0�6���S9:��u�_q�;��Բ�oe~���a,Qy ���D�g�[���IK��H��`$���.���;�HR-e:6�Y��$O+����V� ���=�wt��X�W2�ʅDyG�>��/0M����5�I�u�w�u9�#q���#K�OS�������>��$ICbm'�K�ȑ����)��ֵiu{.+mߢ
$�<�Q�Ȩ&^n h��_��W���<"}�,�w,��cm�3y4��7�ɋ�>�ls���B.��%-�Hwx"�O�;�k�ӕ<E??�P�!�Ě�d�j�A�@�Fdď���w"�q(�$��|�>�r$a#��Ѷ�^�i�y�[���@ ���-jH�%H�� ^K�l��|:t�5S�6�~e�o^������Yc��}��������H^RHƮ��N��&� �a� �T���3rF���\]��)�' ��	�Wo�㯢�zڎQ�j�g�c�%�Sf�]RZ��E2к�a��#��ulH��"�ZE:��>��Z)�ӱ䅎w�$y�:���AJ?�no�_<{��y����]0�j�C�b:���1� �� O�u�AO!H<�X�F.����N���|�y, ����X�?h�1�X�`�`8�}S3X���@}2�O��<Bokh��]P|z@8���^�٨`�M	%�RS H\�.8�L�6��q�u�ʤ��$ �
̍e&n~7��)֫����s�!�ᐵ�y�Op
l? � 4���$=#$��� ��h�Nn�m��ý�c,��V�҅�f���U;髨����$q�xl۪5#H����g�7h����앴�WƔxg�nn�`����y/X:�as2�F��!�m��&P��7����p�������q�65YЄ�e��_R���<3u7y5�΂�1�ɮܔ��_���F�uc���s����N?���09�駟s?���3،�!-0GV���\���'��o g���F��wNޒ����/��������+��}ٗ}ٗ}��,{ d_�e_�e_~����[��T���|;p�׃�-��������˵د��H���'����498�'O�ȃ��r�o=`:< 6�N&�Z��[Y�Wz�si|��ܜ��8��zX�ǒn�2�/�,�g�ezx,�_��C�^om��i�'��������P��o�V������y�J�QHC�����OB
g�Z1���$Kd��r}sM>2 ���0+�.�k3�-�@Ks�ʫJ;H�ڮ[6� 77���@[@�m�0�){UJ+1� L(�[2�m��	~����m������D��C�'�"��ٮ�����1)
G�&2�!��U�ૂ ��ŭ�� �J��}��r#���7�HVkq�%iL����+���+�U�:=��9i��"��^t�-m�'�#���i��X�0�jd鳁�ve2kQ'b�-����fi�����(OfR�RE+a/dX{>q�{ 8mv���,`Aj?Z��sV�Afn��HJЀ�@��ln}����6�{[����3EB����t0H×�(��y]�q�YZ�Z�- 7w ;�5j%N�.#���ms^�x��k�O{6&���A �r�Z���x������ÃZ�x�2!���h&��$8�;`����EV)e�*f��c:��� E1����l�U�<
�����H��� +R���Rϴ���"���E���Պ�@��#���c ׬!C�v��}�aӅ<`���f����΃������+)H�����~G� 弔�:����LNuK�yM�%������0�re)XWu�ck$�.  �/���Z�YGfq�}����#��׾h�=0<��خ�Y�c;�Q5��#Y����H��u���)�т '��\?�������P���yLD�?:?���z�zG�����E(6��͕v����qSI3�x�p8wt>Hn�y�/���h�c��06����2蝉7��(:��2��s+�e���)�T�4l�Z�+���H�$�纈E��݉�J�Bj(턹����t�
ҩԡ�D��G�ɀTA��>�b��цM`�;�L�v<T�Z9)�m��m<�S�ZX�^�����A��zA��U�����u�k]���q h���Jc}��Xۧ�Skc$p���έ}9�ڡ���+}/�a7��e�k&��e�z��x���$O�����օ;�d�j^^^��I9��'��l�b`�g4�S	���kAeR�&��@I�\�	�. l vV�/��?��~�[Y��HTA�5K+>��t�cs�gӧrv�Pƽ)3�\�0�m};6�׏��G�"���5��_CVP�	> �u-�����>�T�X�<��An�׹��Z��P|�^�fћb����0� D�^���n׸.=7�ۊ��&y�&�D6iM���^S�� z��@�D�z�Q��28l�º9B�9Mސ����եIv�!�mЗ��$5���~��&��d�c���+��>	�*�[����Hia^��:?&�Y����k,�o��d�R����`�E`�'5�+�(��~�\�P&�>�>$-�a�#�?[����vOж��(]l��������IْHz�w���ݲ0��P���yT��V����$6�<\+�{�ߺ[�e �
��c�pM�Ņo�F�/od�����u`�|[�׽~�z�1���3]����a���~���d(�����ȣ�3�'��^�;��}ٗ}ٗ}��){ d_�e_�e_~�)�UÀ �7�_���5U����؃G��X/��|=�/�e�Qo;dp�<�d�Po��п���#������%�q.E��~N��D���{4b����f>c�^8�'o=��ח�?�B���dϿ����������0=���^~����ǻ�'zo�x��i�h�N�w
��L&B��UӼ�9�`J��yM���f�J����a�n{���I'�$�k���m�5�~@gf�0P�}�fsm�P�þ�N�q��4)�l��LM��n=��xco��K��5�����ߡ����`�0[�$����&е�l8#uY���������K2�=��xL �������g�FC2a@B�7 �o�f� X>��e52%}��5@�]'�/B���Z��^ǽw����N�|��a��;)����	�����v|�%��̴��v�h �����@m�Ҷr`��ju�;[my��(A<�5��(d�����u�=J� �D0,(ԛrh�Ʒ@��tv�g�J�|3Ԙ>M���I��3poj���=3�����H���i�m��u�uxOҤ"{i��H�N�"��v��Mb�<��;��[f؝Q��oA�� d�,cɐ�B�ѵ�]v�,�uB���%y���\>��K��n��X�l_�����R҈����8<����i�T4�0�K��0/����D�z �ɘU���~����|�z�?��I���yxщ��X�t%RDR�3Y������a�P{^O� �7+���<��3�d2�ǒ�I���E�10�P�%��?�z��H"�8����h,��H�`(����'����� 3�1��A3}���X��֦*}���͹����W��q����+u�fVH4v)���鎏87e�Z�tIi�@�rM	P�&���< �r��ěL�#O�$���B:�@?+�g��yӣq{�G�!.V���5+@;�h[t�~�M0�t�	uiFc�&��z�@�����6r���3yL����L�Y�m�/)/Fl����8�IW�R�C�+ײ�Wf.��3 ���1�v]{!7���%4s.�31v�s3Tm�ф�����|!���'�.?������'3]k�䁌�����|�\�ߜ�-1_,����?{F�*x9aj>9{lL2M������E]��, �#�k~��T���&����X���_\��h��xAˊ�}�b�a_��b-o޼���gh�����@D�s���Y�7���ZaH���t)����8��v������������ˋ�=��:�Q;��6���\ȳ�t���mvα�{bb{7`�ڡ�|3�s�MLD���M����Ou�Y̗�e#�}���׿�b���b�k�<|��Ȱ'�]V���z�UB�-�_�5���|�-U��%���4�Z��M�H����~S3�M��sll=03��PSFk׵�|� j����Pk��e���S��Q<�5>�����M���Y�X7t��n��*��.�N�U��њ�W�Z����ٍ�L��e��V��: [h��r�y e��y�\g�Gh�ޚ���(|�ڡ�/l)�2hk�wkYݮ�[�;������2�O{�L��+ʐI+X�Ccx�:@�D2�֯ԵV��"��dq�S� ���������m��T۩ۍ�v�sFm��|�C�>w��`���wH��Ͼx!?��������������>`�����ʗO��x��8E�`L�����)[0���֟����o��O?��������˾�˾��~� ��/��/��{+_|�e?�4�8&砇��_|!Ӄ#����-�=�y]��B�v6�@���E ��������W�|��'���H>��G���v���^��4	y=Ht;<�"p]#�3`��@/��G"d�d�IU(:�N��[o�_����������7��_�ӏ>$�0 \2[�t�����F3�� 6 �^����f�8�"��b��tp���a��͸k�@��j)���EȮD�a�!�=����֬�d6�b�"���x�فld�A�Z���[� ���g�pLz�@O��p�	��`83��^�q����l����>�,��r��jy�0w3[H����`�{}�˛�o�Y't"#0���!5ss�=�t�< *e�����SY�M+�D�vGB=P7��@G�G�/�j�2K��V�` �S s�1sj�#���X��Ȥ�!�Dv�o���w, �����@�V��G���۠=���{f��mH֨�<\�6r�� ���옄�	���(�ה6�R�`���uŲ{-HR�G�l��4�"��b��K������۬�Y�h���i:�.��̀<���_U��H�>�{B�G`%��J��:~��e���k�t�C0�^��@�|�c������{�q�J��g�K/бY��㣌�@v��r�@[_���d�*�
�8@C�(p$�: H��2�pr$��x쫅�;I"�ŭd��&ű�)H����	<JL�G%}��P�'��3Y.bY���%� ��#@⪧s%��=�} ��h��}��8am��Fǽ7�z��$q��{G�<9<���}M<��63��?�m6�.��>K�:f'rx���?� �;Z�S	��R���q��~O#	>&�������=�\��B��R6�7�8QD	��B��Z�]m�^dse��}*�d~��r�ZV���pԗÓc�>8Ӿ3�M�JJL��'�t$������M$��k�s�����4�O�L�\BKhS�S}���×	"���<֟WZO2�/�P���P:S�i�i�m��z��b������G^�h;������6��~��&�9����5���7 � l��J��/oo�G�������8O��=~�X�W�3��3�����ƥ�m�%R?���^��qy1���c�
����6Vv#��5<�rjJ[+�w��77ײX,��Cb@V�r}{+�/�- �O6�y��q0�]KJ+�_�h�fd}����1�`��}��F�n��� ��S��h��כ�ou���F���\�<��b��T�ze\�˚ƹ�r�7��G_�m����[)�Z�!��jάw$	xu�9�!�UP	��y_��֣��� ���J�(� �)��^���啼��a�u�H� Ƹ��yF��)8��Z�El�����3	��Ћ�ܓ��޲_#$f�/�d�K�X .�&fz�دQv�iZ�c��'�G"�C#Wpl�1?�۟PR�cb	Yn̟��Q�W�;ƈ������(��{J�]u/�BΪ](�
�uYq?�p[v���f�7 �a��$��5���J���.���r�l��1C��:�ep���[Jcp���d��P���}U ��s�W�������V��Hy�!��c~�g��1?�m����/��j��`����פ��Ծ3׹�ӏ>��2��|�O�D��O%� v��x���z��MZ ��
��������97�=�c �������9:9$�?���˾�˾��v� ��/��/��{+�bCcRd�!0;�h���`!�I/��t�!Ou{<�Ǚ���Lˑ�PH�dyB��*��O?��׿gٗ�B�H@�G �Q����h��LTG������^�i2�HYT�������������_�?��������������_���i��	���$@Pi�Z����B�\�szm����c6��X�v4���-o �Jiڃ~�5�t0#њ���h��N�<�uX�V�@l��}�d ��X��l�4I�֌<�r���!�]J�z'�`3��Z~��l҄A�!�K���-d�R��7;������i`���B]a���u��r��R0�W�l���B_�13���x�zy����:�0ĥy;�
�A��	J�?�=N�)��AS���d�F}Ş	�`�ֈӡ�U���Axi_fko��:�7����lW�dI���6H���4�T��}�[���N0���=f���b���2V�A
�4�h���Hɶ�(�RI���ΧA�o-��W�/��;��P�a��	�* �Lݥy���-�/�W�&s\�Y�u.�g�y^���5O���,�����#�P�2����^��]��h�G�iV�wA �̄�|��p<4�񨧎~�/z�i�r���j�%�0:�r6i=Uv~� �O�,Jkݼ��3�k h��o�2A��;���ΑZ�^Je�oN��精y�S�R¡Σ:��`�s�G:�:/�I#I�+I��R���)M�7��D?�\�j���R%7ڶ3�t�����v�}��(��/e���*��X����PN��%����v
j�*u}�k׋�z�\f�X���:�yp�])�����7�`<���;P<����)��[4|�	��� �x0�.�D֫k�Ǎ�\�&7�����aϤ�u=H��b�'�R.>�L��B�d=�bH�����1���><�w*�7���,2�!�  0��z%MhA[u{#9{�X�c������d�J�]��f��:l֒��R�ʣ�� e��=��n�x2�6�L�a���j�!`k��$��݇e���XĲ�*f`@s�ڤ�|d�'�7?{�##CO^�z-}�Z��	A��֭���ίx��5 ǆ^�� ����X�Y�}v]�dz@V �j���s-D���+��� �P i!�!�h~G.�� C*%8Z����tC�ҙU��X/�n�2_-���dS�`.�`E��$�Y%K��LC���kkVZ��,͘]\�u���\��-m[`��0I�y	����׷dv�T:�non��rf`~lA�^�+�~�}��>��Z�mZoy����օݷ �a�H��d�t�������ں��Z'S���{,�<#��G}��\����	�l�ÃC9��Kp\�P�mݞyM��\)��[�:o�-���}��Z���sp/�w��/6i̠>���k��x�����I(9ׯ~oH�X= <1�4}0��y�(Y�}T���ݲ����dK��	����}h��J��o)+�rbX7��A�'�A׮�[{��ٶ�X��nA[���)���pl�Ѯ�&y��4�E��QH�@R��[]!C�h�B��L�M���.�6��;��k�6�BPt��~q��l)缇$����'�z���&w2uI0����K�B�W����\���|��K99{��K�f6�/>�D.ߜsC@�	)���r]k�B�̝>�ׯ_˫/��20����@���>' ���H�e_�e_�����}ٗ}ٗ}�WS�u*�;����_��x�@q|�oB�?d��r�`P��T"?��d��t�\H��|�T>��#=<����J/��]=�#���1�ɩ��(�	x�̪�27���&�꙼Ѓ��/�Ig�5c���.���ɻO����������cy����,f2���vB�Ys������2�c��ܘ�fn����2?��[�:��xdCF���;ml��}N_���L{ߴ�ͼ2�8��^kF}/��p��rq��L�I�&�8�{��b���Iq�����8��%Ȍ������ЌAr`�]k�R�H�@� _mF�8�#c�t!iP�G�Z���,���� l�z+ � �3�۠?0h��9�8v�mHH�w�������@�ĥ$H���o�q�qi��^�櫥�uN��g^��� =�C�Y6��do�o�|%�a�
�@�� ���f�NS�-�p/�/�L�;��+co�"u�G��+�m�H��q�A�Z���0����h�N��1y3Jo���@}�o���j/�w�C@��"rg�n��b
k�+�\�����H���{��唴F��v������ޛ��q]W�7��=�v�A�i��,���=3z�����d�%�����P[���s�,P�W����BVfF���=��c�������F�i"��)2�!WG���n�C�����$9����`V�u؈�e��t�:�j5��݁$�0�f 	T�a� u��͌|�4y}�T�ä"���]�H�>�*/e���I�F��L��s�7��G�?�J,t�X���:�tn��6�H���[2:,$�ǈ>�jq�ԑ��hF���z-~q%Q3�N��=�o?ƼP�f1��J�)�
��� �\H�����/���}�� "��D`��������D�km�WR-Oe��H�O�K4:�q�Ӻ��l�����2����$�wd3<�
��U�Q����T�^i��$y��{�,C��r�R�R�i(��/e~�P��_鳮����2"��OF�����a�m��2�h���]$굇'4�^�5e�:�U�6��rzr�����O�+�2e��Hn�}Knܽ/Y���>���Ҫ�t}���*�)�G��uM����@	���m���Q�})�?��VTN3����s<o�Hv���9���c�H@٠��UW6�|�B�o�X麋��s��*�!�T퀕�Aڒeu�K���V����Jg��ڹ�3l�����"�۸���`qR?����
���tzL�l*�0���OZ�[��t�з�۱��]�C0cПV���d���s�C����L �3"_R��e�P�L�sw�ycp��s#2i�R�*�[;9�^���%Fx�wdv;!%@�CW�]�R��l�4�g$��Ϫ��1�c��4���yC�}��Wg��Ͽ���R�~�L.��ڟ���M�!9�Hh�8���FگVX+�����ܸuS���Vْ�B�������퍥�ee�}X�Џ������.� 9��-fs����1>���뽾8�~v�?���*��H�c�f�+ȣ�`_�~�^^\��0O��6�˗/��G�&��_����:Ǎt����۔�#��[�V�Z�����u�X���3c'1�,����l�pc����0��2i�o$\��HU��v�Mҽk ���{�y���{�3��z�́���F���5��7�~ �\�� �����:���`ݼ[�!k��c���7E��ы��e���9��@
���E����������0�:��k�f�rF6�a��8_0T�l��/?�R����ږc�g��/��;�]ٕ]ٕ��� ٕ]ٕ]ٕ�_��$=�t����~���=bf @��`�k!�  ��$�@��dh+����y������@,	d��}�gz`*���y�8�UYmn����@�Ya0S�h�}y9g���}�=��~$��[nݸ� �'�������^>���N^��}�H������c����x��K�o2��� ��`�K����6��nPp�l�V~�� D0PL�XV��4]�?{r5C��BfӅ,�| �����64��Sfd8�Rj���ł�e^�渎"ü�߳��gpX����7@ �<}��8��w�TO�JNE�<���o��"#P�;"�C�}�\2�����P�=$�)�Q A�g�>X�t����%�Am��~�zaTJ}����
�5.KS��F��2�@w�eL&����Ȅ����q�g�G͔�i�.i:���������,[֒��Z���=�����:�Ƒ�����	KA�7���^�=�.D��&��A*��[��=���@Fj�A�2l�}v��@e`���z Pj�G�\��>���J�^�]'�����^ɖz�z��4Z�}�a\fˍ�d����#��� �Mݵ%����L�/��o�%cm��H��$V�������EW�q	���;�h����R%f��u��+��iBH,ulL�|y�cae�j��n���I�҉���16�T�@����d_�N,�i!����2_��:%����}{ZWcYs��xk��\z}�`CvG��ez���t�kz�c��SΡs�ͩ�����R�2�>5�D�u����%0����!�,:���_��ť��<�?�#'�P׆�>�΍:�!���5к�r��^I��Tz�$��h���B���T�A}&xS���+��*��q�u��"[�buA
 �\���:�z���>��d4�ɠ�����l��"o�{x(ar�� ���� H8'0!�V*�����I��������X�D�&���ȔB^n��Ӷ���߹�:V��Y=�~�i{�kˑ��\�׃}ó�@1�ʙ��B߁�,�V"d�.+9�J��H��7��r�8��	%op����j� ;ĩ�V�%�NO����:�9����8�뺤�`��}S��P�����}�H+�c��ü����p�g��k�Z�{�[�A�\���2e<r�Q�ruEp�����O���r&W���8�ǘ�X�W�W���h ��=�ǁL���2%�W��7��B�����+S�J-l��5	 h0?��>��B�RfW�����\���j�{�j�h���В=��`2_�j��pxu�[?.to��_�Z���d� ��,&ؖ��wfٕ΍H�~�Z]�\���{䣏?���ߗ�ބ�ak���H�i��1�$<!���# /�� s1����^���C�ρ�6��Ze2�MA���% :A�~_ 2�t�?\!��Ɇ���>�^��%X �������~���=@�,������b�Ao� �?I������GW��'��i_`�Iu+y;s��j���Ssߵ�2]b���ڮ�!�94w�������ĺ^����w037o�ZbHR���5����%k&�G�8A�W�c�Zi4�3 9�6y�];[�
���+m�F��v�#�WM����f��7~.��Y����~�`[�aH�����Cs�ҵ�௾���?H.�(jRi�{{��:r,�]ٕ]ٕ]��.; dWveWveW~��/�.�s�cP��+=�䫥8G��Z~��ղ�
cAԞ3ax��7+J��i=�� ���j%Kf�/A�4�q��#$(p@E�h����?xG~px �}�my��f�}��g���c��O?���ރ�������ܺuB��b>��g���T���6��2���(�T��4G�f����%�x`v 2`)'P��d[���A�����gWWruy�u���=&��U��,ͫ�h�m��@�o�uaM���Z�B�P&�U-+���yp�l�؏i���k����A�-�x.0`�iC���_�`��@��3�	�మϏy����#`����rX�߇��jA����Ё��fsY�M�C[(�#S���6ecp�%A
|"FF��3��}�f�X���l�m����{?����cG���V��������̰�wl�V��MD�a�ݭ��"�F����oY�^Q����M����g��ߔm")��k������uS_�3Ȝ���-�m$.�0�k�D�����h�Y�eDP`����V
΍	�`�+�>���l�w@'>���!{�mt����N���P�f��f_�K�t���X��/5MWS�]��G4�8L�I2 )1�H,|ٔ`	��7�!���AU�^J�o�����#�Ŋ��x�"z�$���C@�NW��F�e��#o,��mV���Cg���x�����&���Y7S�������:��T��T��gSB��\kB�L���m3�Ϝ���߱�b!i��$\I�{�g���V�i�����ظQ�׋��W���#5vDN�2?��y��l����[rt�@�L�C��n��p_�^�󓶅��Z붆�D6�J/)�냡d3��,�\�ܻ#�#����ȁ��k�е�px"��)��F�u��`�L�a��6���=��0��֏'�G=]t���
I���k��R�8��r��=wGi -�lt�]K��g��/�.���1V@2H疜wM��Mc�	�
��D����΁��ϲdk�k#}��"kƢX�'�`��Eh��L��u�z�ky����<{� ��>Aĳ�Jvs�G���
��$Ҿjc��SX�=HXvѧ��=�U0@>���P�NX0�$�\�p��f�(@��h,LԵ����w��y�~g��|��G�d�<�T^�<�u��M�����z �\�g�Od���kX��&�Od�^�G��-K}�Ǐ�Ҧ��7���_$| �|��J.Χ:Ʈ�؅����x�,��
�F �>0k1���1��+$ m1�?z� �:$�ݠ��z��<�92���&�x���P�ݻ'����H��p�)){�km�A���eH�y���.[��(�����:6ؗ������XCC���'iQ�3L�h�{����%�|����|��a����Ů�e R��C �b�l��#���z\��gd��Z7��"q�to4����\�~����9�\{�'l�48C (W՘��7!�o��0L�jw#�^ݺm�\�9q�%�;ZD\}���w����SM��=�5�e���q��FyͶDR$L�
�Ό�����AI��]�زH����*�ڧ*8�@��?�4qu^9�x�����`�Rf.�|�D�ơ~ ������$�o�G��� ��+��+��� �+��+��+���CK��7z�.b�yЁ|�"�O��I%�=f�g���p���� p(cVw�0�]Fn�Ё�9��:��AX�(ɀ,�"+��oAhH#�s�2�XHbT^A&
\��Xnܺ-�'Grx�Dz��\\�ɧ��D>�ͿɋǏ)	��Z w}%i�G��/�ʳg�)���2�/	<@���8C:�,KZ�ÃA65�n���8�*A����?B�8�� py�f8Hz�S�	Xp=`�)���2j˖�uB�u��QR�&��Rk�� �`Z��.?�9�A_�b1�k;��YG� ��n �3�C��@�βK3�'�Ĥ�<ȓ1��o�V$N" i�j;�&��344-y��"t��h�4���g+��^!�N���f�vq�wd j�=�;lq�1Y'�K`]��7��Q9�Ȟ������`8��IRy-ۡ	������q������m�`{]���Iv\+@���'�'[M���',�H-�A�V��M�+O�A-��8�	l��k�L.�Q�<�}�(ɛ��EV_�Ft���-M�|A����V��w����u.yU9 ʂ�|�m'�4D��R�`,<��u��vc�u{2�I�70�K-4J6�3'�	�n��B���������Ȼ�:_H�z"Epُkz�0�JfG�Uӛ%f��7�Is��1���Wk�ٍ~�Ʋ�;�L�TkH��K�x,��γg:G�"it�"�~��ģ#�6���@@���V����PY2���Xn�1S��3���|&X#��Z�-�K'��&��B��k���:s��
���htK��/�ιE�u3��5�y���:��F�ޗW��]}�D"/ѷE�u�Zz���/W��d:���R�|&M�W:'f��%9>��ȅ��֍��VXo0��h[�gd(�X����l�������&��u���ڮ�\�s]�:����t�sU*��K��9��̵�Y���2��mR�t�)��T���2_�K0�gk�I$3����LיF��':W�+�>����B�'�uѰT:�6 �u>� �u���ð&�AR��Z�=̳n6�2�8��ڂ�Xu�Y�c ������m�� �Rx��` ��ܔ�ߖ��c�ח3f�#Al�Zl��s]s��'���>�`r����a�Y������s�"8��1c ��1��t��~c&��b��9`�M=x_T`
�� K`�ׇ4 ���P�NV����Hi޸}K.ί��N��{���J�l�O�BۂA��Fnܹ'k}<�$���y�K���._�ʏ�����G:�*�˩\� ���jA��%��}m݇ڦA�=Z���(�qOt"Z�h~1�/P^���鉲��}�� ��7o��q��[L�(�����ي�P�^���c���!/tr|�� S�� ����^��~2E`��͋Xc�?�C�d����u�;k��>HX�6&���d��qh�5d�竂�G�e�r�h��(��cs6�e|�Sxp`�5�$�:/�`1*_���,��{�V
�'���GK�H���ѡ�=zf�}�q��R�Sm�?�+������X�џ�%���>Q���J�V�K�%;k~މ�y�Q��YC�c=��g�{O�ao��� �	����C�v�ڒ���P�Β6�C��	}��nBi�9݀��ɭ�>*�G���"��rŭ�����
�ޕɁ�!b���=�x��B���098����o�yweWveWv右� �]ٕ]ٕ]������"��C�p��N�6X��R�(����~�\�$4N��9����Բ����o�m�2�i�;�1� �H�D��x8\#>`TU�P3�txt$��y@3R�7>��<{�X>��/����Rg��u���{���|�B¤#O���,�Fa��td��a�]\]2�����h�#�3NEP��8�,<I�:t�M��s2T�+��K(%�8r�Fc&�I����w��@n��P'��FJD%u��ICz~�e+��K�M�mFv���pY&�ח����SМ�ncl�E��T��D�	�/�y��^��30T��[���4�D�O#�<�C6��=��x>���V+��^.�2_,Y_�n8�6f�Y�! ���kW�k�k�[�3�=Ș-)�bL���mW�]���B�f�lB@L�)���V��"�뺸6�vbP��arO`�p|��������w\��JX}�A������,+[�p���k4~�����m�Hn�:��(lO�V���9Ý�kr}�'�겺\P�?(��jJ�x�A�V+��6&��{�6����NJ2�����c��Di,Grxx"G��2��	�P�%5�0����,ں�h�^.�'Wr|r A���RRb5}_�s��M�R��ZҞ~V�7�M ^1�$�erxG�>�d��MF�n�9>�B�t|�/�jz.��B���l�=�}�HǱ��p��4��K'�#�כT�H�/�)Ŕe +m��H�p�sžt�#�Qe6���kI:Ȏ_�Z�q�'2�2X�I��[d2����Y��B9��O��Џt�it<�^#Q��y��g�z�'M�<قd1ׁѾ>õ!���+�o�~*�5�� -��{:'d#I��x:>�K}V��p$��@�$=����+:�@�)_�P6:�� �;��d7t 1(c��L�$m���5�]H#%�!!�G����K�Grw=��b�����A"q-W+�(e�AC��No��ٓ��Ȇ����C�sT,�����Ӿ��9��^?е�c,C}B��� l@ �ڏB��N�3a;%�N��;}W�������!Y���؀���8Ɖy{-���Y����=^r�g�����CN�0���+"�qֈ/��>3��y�va��E^�<�թ�����`��q�{�,���HU�h/��ᦠ�X3��L&���Ƕ��^XC�s}��&%X��I�}�.����#��C�Dk�����F�=����� �F�d4� �s,�����13�� ���G7���ۜ��N_�Ç_���Z_��;=Y�4~�3�#�4+������S��@��c��rzz*�������-׃� Qȹ7rҁ�%$ِ�Z��c�I͌|�gЍ= �?��H� cc�d�4�20{����KJ�����U���`:�.�+V �gS�@��!�E�E]ғ)/&���M*K׃��'�\�IT�%d@> ,� l��l�:�\�\��A=`����0E���ږ�x���@E�enp����#�`=z4@�NLx�(R�� �#�E�-�1J��!3T�]��{[G/�tۘ�j�	:wmh^��b�!�(�CLki�s ��0�Z�Kkgb��9�>�^I���ra�E�{�<竢c%�y��h��y�� `�3ڪ�eRX��� ��^����mVk2̍{b̏G����oˮ�ʮ�ʮ�q� �+��+��+"o���ʲ.��D<=���# /��xq ���$CF��Fzмw�]J<}�\N���qAi!�\'��(� ���>�����En�b U�����~��Sdv���;���{�Ny��k����gO��Ç)m�2�e���:����t-��<}q�x�O	�M	9�H6��7$�7Jf��<H�!7N�e�; C�W�� 8����δى�Ei!؁�Mz����j�Q��tJ@�;�e<�@0
�0�����!�*3�h�!+y0�hu�p/�'d�n� �k,���d�`�Nd�"+ϑ�kYo�2��C�7M�a
Z� �1��JN��x1%_"�o�F>U�ŏ=��"���{|Qd4^Gv�l9c?@ 0C0|.�LC�ä-LO0�|�(m�-o�v�����C�����xP�ƒi֋�C{������ s&v!em>��h��ۀi,*
� 4��ٲ����o	���lk�p��X�!}AY�`\�> ~ 
��r��J�1�	3���I]m�/�����~$�F&��kx	��@���xA��[���O()��@�jq�?������ƌg��B�)줔1�/�|������;ߕw����й�y��@�B��罽	C6����x%������%d���C��}��z�&HV�k0#G�o®D:W�����;:��PYh� R�K��s{�x�*t�����oV�,.g2�i]��4��C�=�SȆ_0�n2� �e�߽�W:L�I�~�e=��ӋY���]��ɠsS��-�L�tL�����/tθ��t����RTx���N7�� ��	��Է4_P�T��9<�)YpG�ɁVM`1,x��.�.���Ϥ�}Y�K�tu� K �A}?���'����A�d���!P
 �Oq�#��X�Ro�-�S	=�n��;�/�:��Fש�/i�H���Gd$6z/�r-�b��(���($ϖ�W�xKM%#��<D ���GKI���K��Ɠ�ו�י�Z�f�� �h^?��>g�}���N�F8g7�f�ϡ
�n�[ �\�|"C �2%��������@`XZX"6�4�1F�Nt�dsx������/w�<�'o��h�2���1�
���=&(ܼyC��XU�`¸O��������с�@�A�� �� A���	��d�0ƴH���^��rF����- �.�u�)�����͍�<�@���5L-�V�	�F����I`|Jb�u��s�fЭ�,<w ��}Ͼ����@��g/���H�nݑ��\>?���N�-O�Z�ʚ��hC�G�������z ��.����R_���'r���ۆ��x6x"��@��/��|�O>�o��!�>��g:�.�	����?��<z���uNø����Z�f��ӗ�t�2�r`L0h�X�e�@��m�d���;�^0z`,���k���nߐ��=� \�KȄ�	F����!��߁��z���־_  �W �i����6��6�˖���O��oc�-S��D绛w�K�G�=�kV��п��q�����"�]H��7�ާ�cr�L(i�D<ș�~{׊�א���#�I-���,�Dh�n I��g0�!i.X�@b��I0  Ly��dM�4�5�nͭHA�H nO����?��k�g׹17�֣�g={L�	9W��b�MK�`R%C��T����:E�
%-�ǆ���2��ֶ��(�pN�L*Yi���RG�$t	CH�y���\����<|�PveWveWv叻� �]ٕ]ٕ]��*8l��lH)����_(�5_.�凃]�7%�z�}�c�����5�%�*�����~O�ܽ%�^��Ͽ�����SJ	�Zd�ΈA^��2=���@�z�-�*8Ğ_^��Ǐ勇_�����\�ma�o�l�X�K9���2�]j&�iܥ^9
��@>��ơ8pْ%� k�Cޫ����,�7�d��iM�</��="��{\�ZMcٰ4}�C3�d'z��)mഺ�����ٜ��o����\� B蛤�ȰD`����s��`Q��k 
�6�Cg[���Γ`@�S؜:��:�3���=2�i&[UN7Z��6x�>���4q��'�'[3H��::v`[g�;�ɬQ�}��P��갠y�_��d�Rj������L?j�y��ݔ����\���n�i�[P?�~ns8��!�)��N6��cڴ�j��y���I��GM�$�����tU�i~��¥dQ�d98I6d$Gl1��Q��z��U�8��cc� `���T.D�X&�ԅ��j��NR., �>�ܟ۞�f��>��K���~ym������W:��Ȟ�%�ALݷ�Cd���> Qd�����l��vz���"�ͳ��~]� �)�:	�|�t������5�H[�ŀ�sH��~W��'M����~=����_J���0�z�Ν�r�⹜�^�3T�x�O��#k6��C̥)ȖB]x���0�F?7��y�C���:�5r�j.��g��uu썵�z�6��iV�o.��{����3:c��4i�q������e����DdO:�T�λ����HBx$�0^k;TdWP"u�9���ӹP?����9�Nk�R�	�m�ѹ�I+�Ҭ\�@�Q�����	��<)f�G�ģ� ����I���qN��,�g�/t-ȋ��uG竁v㘆��,��:���O�?��D`r��߈�����/����A/��ӶK�$[�$��_!x��L�jHt](��n]���JR�TZ���>� 0���~
�y��3-c��5��0�>����	CD�HW�����8�"	`;<7�D���Y���8�ZW�뗗SY�Z��5�3�k ��Y�.}��g��5L���5�72��5%%�p�`��O�0$_�u�4���7�L�n�H�G2��h�̴��u-�b&3����E0�'N6	)�QO�&ڮ[6/7l̋Y(��6��N:�����lq)nձ9�I�E ���'���������?d�����hoo_�����;��/*_=�R^�<�G����_��|�������I9'��5��P�7o�Ҷ��8��ןH�q��������~�X��^3�M&���X ?���ZN�3�7d����)���CRN�+߬9��?�\F��'�Jʔr� �B�"��ndq`��D�2�����F�"���8�l��	E�m�~0d�$��9ظqd�`W!I������} }��2�;��a�
���Od�Ldk-r;0�	j8�#���j��3��zݫ�s��*g�n���--ę~§�f-��Uk���Q��c�.,I�#k�����m`B[c�y =r�X�p @^�G����c��k��zv!�sNf��Zb�'ǐ�,�T�϶������s��B�֮����a�Q`vCڴ�s[�|��Hhٕ]ٕ]ٕ?�@veWveWv��^b�96�l�^�34�~���v�.���+R��L�5Y��e�&�.#3���<���j�3�����ӗw�-�_�Z��]����y��/�UzȂ+���%2o����CZח�~���>�/^������O� NوA7eP!ZH�A��O����u��.������pxK;1m �L�AhcZ@���4�}��<�ڴ�q���q�E��Ud)�����z�F�I|��`> %�{�2�TF�A��xĠ�r��L��r5���'�m0���2�n#����\ƣ1��|OabLx.�sՁy�
��Ͷl�a�b��R3��7�TϙLo6�;ė�ü�4���zk��&�JE�>�ݐ�uCo:����I]�d!�4`u���V&!e��O�vHZ��{V�jx��I��jx��]o�lS�I!u��kA+[��N2M̌��]Ь5�<���h�>%^(�%�,��`
�SYd�"p��RJ����d�ǈ�kSck&^�Y��9��=��&���km�@�������{cz��7���4���Zy�s��)J��A_D�	��;}?�=\m�w����0���<SZI�:+�.	��@G�'w�����naƫ��Ǎ7�	]0�v�'z|���3d�
�6��>7L�i�Q�����)�Z7N �*�S4�I�y��M͠�|q�sѩDri�F��$���_������0`4��`����z��7S)6�B�s zɮ��H����>C�3���XR���/���B����I�#K��4��l��-�-��nG�g�I�g�G�r�*�q���;nW_އC���P����s�%�����R��km����BR����j^H�����x����C��Z�<��z_�F��n���\�X��)�=&��y1��]���ɋL��.B�+�`_�{�R������ʃ$`]@M��֗H��ɴ�*����13�1^Ms�a�{~���d#/^�z�\�z*��˃��W��t�̧��W��~��p��F"�}��h���#Y�{2 Q���V@����hl9�d`p A�B��̾cxMi�u�X��c9�w(����t,U4l���ӯ���ׯe:����s�ܾ}��-&����|�� �e�@NNN�҅I!� 8�� �g���G�:8�����dib.9�׾�kr�{�����k�F�뽼x���5�ߓ;��Y���F�L��)�����9XM�����'�!����Me2��C&�7�K�����{6�@q�,�)XS竩�W}�������J��g�X���;A#�~i�����폾#?��?��#c0� .h7ڇEo�z�u�X~���(����^$}�]���+���[���VB}û���f������!ܳׯ�ɣ��vNB�J,�\^,�/���|���ߙ��ۮ�� GX*�< ���1�D�肓`����<�R�*���"��`h"q��3��K2\�����z��c���P�����N�V�r��c(����b�O�� qݏ����79���5[�	|<O���{1��T���!�%��(꼽�vC�,h�� x���O��Mdخ�`q��.o�-���ּ-;�1J�tc�] X���X�u��(JM�V��T�N2s� �n��ȿq�ڤ'I��z_�}j������un	2m��s{=0_�O��1-D�E�-�O?5޿YZiV�A\�m?�T���W�"�?�]ٕ]ٕ]��.; dWveWveW��Jw4�C���~ă�W?�/�1[�8�����p�,�:LhxĭJ�c�;�-J�ܾsK�}�}����ݻ�T��?��_�V���1��W.�����@�|�)W��������ɓ� ���#�f<��8�r�1?��4�������Njʋx�1��ڵ�<`{|V�Ƽ>'�2H�0R3�@St�
f^3�0�M�A v�����A����<e6ْ��ѨG�`����⫭15��t���0����c>8[�Fu@��3x|0Q��=�h��P�|������/᡼�@��Y�>�����& ��=X����u� ���H��+}?2ੲ�s�e3�G��� _m��(ql�o3�<�6�|���jQQ�ΣN���x�~2�x��օ�z���P�m�	�xfZ:�$�B42)��V3���72�� ��X8_�l���L�Xql���!�+�ܦn[�e�o�y�6��@�0�)��6
�d�1��/2��>�@��x�����dA0�V"�)�m��"0i�it����7�~�\9h2��g�O�}�dPc�28A����:=����<{����i�c�d��L{��y�`<�\ �B�0 �VoM�0-w$�;yd�BB*�z)h��x,���ɔ����E"�vၣ�l5��g;_�#�ɢ	(����p�팺��}�f@ɽ$�u�@?��Oi�"��LdQ��sZ�t+O��/B���Y���
�:O��ˆ�v#UЃdm�1'�[���G�C�}$���4���vc�+��KI�\b��Z ���a��G)�HۛF.ruy*^��$D��֝��W�2�vY폥�q"�^�$����bSS�rI�Y�KY��A�*�K����v2:�B��:�뎘�\�0r.(K&�D��m]
f��K6��C9ݐ�@@
��� �Z�ߋ�T�2�x$ڕd�W��uZ�{�ށ^;�yy*c�+	�kx!iʚ���� �pM���y���u��sz�)0�ϕ�r $���=�� �!6'��Qz���+��[HiI2�ʇ�/�������\�h��Ye~�ӟ�x��9��x(����P���ՙ<|��\\���_�`����J׵�Lۯ��밀�7�"��s���r|r�{�2�]q� O�w���ߺ%{{:�J�K��Ǐ�/��_����������7��S�YWWWd�`\/�3y}qN��	�M����`BN���g�`~�I	��l�%�Û'r��]y��r� �YEc�38��d�곎��&��K��p��w�t?srt(�~�\��X�%�} �W.���g��c�x�u�P�qo�}�d�H�O����{bҁڦ��L$w`��G��� ����9�;܂� I*0=�#�U-g�O�~Rj($�d��lE�(�\0b�PO0NȘ� �%�3���'�������^P� �����E7$�C,"�v z~���]\�E�����n�NI��鳄���<Y�t�2��K7M���3y�[ߖA'���8ϰ����Q�]֍!ɖrcb�����]UZ"�8�"�C���[�!��V8o����R@�}�p�.�_��3U��3,(��2�"��Ê`Li�9�v��]u����歌��	z�D6u��E�d����K��>�4;��L 7�r/�=u��^�����^�8h��Y��%�������S]�b�v�Ϊ ��d�?����dغ�L���veWveWv只� �]ٕ]ٕ]���?����[�/�}����%�^�ЃJ��9@	�� �L��xBi)�Z��8����Mxx�w�<����W���Ba�@�=��ٛLd��pu5�g�^���93Bq����@nVz��ve��IMk=�"h��;d�A��͡iB�t�!���J�5�ѭR�*'?�4x��A'?�͗#aVbD.*�ڧ��2��#p��A��/�J����p8��L��"#+��d�P � ���j�:�	4;�iw%M#�j$�HPd�dB��X��W�B�ڂ�F5�x�$�`aͬpq�1���kf�9cЦ��A��*B��s��I�0#Ղ�B �$[gl^�`F ��������`��b�
Y�E�,Z��O�d���AVtݘ��0x��E �T S��`�Ʈ�J��nͷ�?@��J.��gi���*�?�[`b��@��&kD�C9��V��@%���TVi���@�Ƙ%N����mԁ9YM׽v�����LbH�y�x�� ����yM~�2�C��	�w�$�����vPCAb�ۚ�e��A�io۾��0�N
�W;I$[�>)�t
˄������|h�1~�cRj��:��_|.?��O嗿���#��ho�� v�u.����Xb�  ��IDAT���q)^����T��a}� ����~�Ҽ��g?��s�}+B]�K}����M�u�I��uEz	!��ֈ�mQi���a:��6�6�9����΃ ��Nh�y����@V:G��\��D�46�g9�Է-�{6��e ���+����*���	x	!��'}��M�D�C���Y�`�~!��B:�Z�$�8�@�F
�G4�~��G��r�E��\N���#�O_���h,!Xp�SY,[��M��p�i�XBR��'�^"k�.)�3�����UNj��cM@�7KW�L*?��BpY�]�s\7�\����u���C��ཀ�0������[Km�g�z)]m�"��D�	f#]W���j�R�s�=a&���tHBr�.ݸ�-A�Kݟ��a5�Y#X͞�߿��`al 8^�Xg6dRlV���iH����:ݣ�T�9��P>�����~+���������B���舲s}��g�+y���\�����u�fכ���|#�`~���N���Q/��:���'��x|�艬���X����>���/����������'�z�_�o�km��� � ^" � �L�3&��S��OE9�˫+�ϗZWJC����C�|1�}G&���nls�{RZ2�YW�����î�)a�F�4�Nݯe�?�����?�o}��< �	ػ0у�
�t�o������|,�GǺW�(Q��0b1��Wu��'O����R�4]��o����s)�� ��SN
�K&De^�< O��� �V����T�|G�rk�t�Q�>�z�A:�<�K��'4��󏹞]`�2[0i s/�(�GΕ�Vf2�5|�}��>��&��?��Kz:�t_�&��>�u!Ѻ����.�����R絬������(�ƀk+�W��7��n����7�,��-�S�v}5VhK���5���\a)e�vs_�tg�ب�lle3�;�5"�b�G�J��+x�.a^GI� �T��Bc��Ú����&cYco]����"$S���sZ�v/k26CqD��j,���,B9���!�>�?�~y[K�D�a�$�<#�&���m}����ɍ���#��_~,��+��+���]v Ȯ�ʮ�ʮ����pD��'�w|$#ȫ�A��[��@T���9�(Iܡ������C�K�,J�`��=�`07(�ty0�ZL����@�}W4y��]����pcd1�&4��Qt��J,k^�F�"�[D!�P�-�r�m�� �c 8��A^�f���w9�-
�д�H���x-�������D�8��q��'O�qR�'�y��xH.���!B�o����Y��44Y&�UjZ�fwGf�2��N�@�َ��l����hT���B!/Q�X�5�$k��='g� =�DP�J��:�����8�RF�kg�+���!=���4F���2���Narlۢb;{�	�7dM���R���6��Vҋ��b�fm�{l�h�Ҍ�M�6 ��6yْ�L�Z�=3��}�;������2,�k���6�+d�#��zm�c�c>M�r(�O��+!�v�=���%�@
u�I<�RƬΈ������ŉ�����)e����N��2`�s�'����d�8o������L��,~ɀ~�B�K�ʢ��3�!ޓ{�~T[Sy?��O�lRd��u��ܹs�������J����^~���!O�~,�Ւp�j=�1�c�9�:K
_�;��Q���/��p-W#���!P�y#4� �מ�� ��1�&��F�WӬi�.UbL�ȗt��`�:YeBC�˫S�ܚ�{:vS��f�z�Ǳ��7 �V�u��T咕fv܄�u�
eN+��$�.+��2�kc���BД�3����O �C���d�K�`�D]�;���=>�߅���|FC/-���Y}�b9���\��@j/! ����ރ��ť�Ξ��'�f�(����D�g�й=[^j_/���u���u|���Y������K �kQ'dh,|.��,u~�i "�w��������J�1�$����,��;����T�w��v�w��r�FG����?̖݁���g2��4hXfc�q�f�m�c����<���9�$�$̰�`�	 ��HZ�"�/�Z��nLP�A`kIp  ��} ���\���r����~�J�k�W��h߼8�Pz����������S�W�W�C �	~$%�g�$�~}��:޵�!�U��Ţ�Čw}�;���z�������?����?�D=|���"^p�;�_��g�-Bι9���b#!�s��y=���3�o���w�/�ט�����Fvy�x�6�ߘ�`躪�����.t<e|�"�����^�{�Tn�<���h�@<x@>�n������_�<F�c�<������y������7�>^��ǧ�~*��2bnݺ��1�fSYA�ͳ���xP�w�y*��Ն���Ї�xL��j�x���UEa����zRst�d����;�����-�����?�����R��#�_���8��f�{�z�<�M樝��4֕��mJH`^&x��7o�;ޗ��7�;t�����ɿ�ϟI
L���jM�L��4٦����g@	c2���eUm�&C�8�S[|ڄ��2YS  ��Lm���FxU����o�:���[`r��;��c�Z��썰��eH0$�l�9�wA���~������k%0�P��X���KJ���;&si�%�{-.�A�̙ɶ�1�p?���Q���>m��q�����0������b���Bn�&�f��ڕ]ٕ]ٕ?޲@veWveWv��t�#;��3#��gh�
�+4�4��F��eGɜ f0���&�C7�(��gÃ4�y�L����bN����}YFq��F��/��7�b��"�2�Z��\�8h0�>9�����,����򀏲ZYd���ހ�t���y"��3YѮ!0D�s�!ȊD�N��Ȩ�l���f�4to�)�e�M�W�� ><2���;�� ��}	��1�Z�ƲJW��T�g����1�pL1���I3�ٌ���e����~}�.Z='�d�� �eUn���,8��,�ᨧұ+8C���J�x��3��m����c Ts� �ځ�L��Ap���i=ABYh{��u{3�� )e<�yP��~`'�H@���}�����x��bF��k `��hb�.1_0vL��3v��o���i�?4 @�`5�kz��ϵ��YE����x2��	V`�{���L�g0n+'p�5Kg��",��\t�jQ
g.]R<��Ii�)�w�o���۟�&��Ƞ�GRSN�G��ٽ�� l���5e��0!8� �p�G���`�����7���ϟQS���>�ƂϞ�{����
c*�A���>������=�:����7 $?�1�;�	j�Y��y��@�� �ʬ*�#�|ԕ���ML��B�����K��K���XMo�>���3��D�=�gK)����b-�,��,~�2������wd4Zh�$����A�j�N�N8nД�mɋ���uHi�n� }����C�n�\<�	2��w1���f��KY]m�;m$
�w��Z7!����ZjeO%�t��u���������y%�t �t(��#�X\0�)��&O�j�(��� "Hu��$�l, ֍�+�΁�O��v�C��K�U~d���}V��K�>edƍ9wf�\KR��e	m[��^.�M(ˍ��9����?<�T�p� Y]n���	�rы�@w�UA)+ T���M1#�؉6�-fl�6�ᝄf6���\�/O���m�"J��u��<����ʸ�F���>�~��jo"9��t>�O��w�#{�����!��*3��p8��x@6��!݈�c3�2����	��0a�"�?y�T~����g�l��{�L�{G���S%�yN��t폆l��|E�����\�� �K�(1��HJ�Bø�I1}ںg�>��v}#0����3�'��Y.�iY��Hn�[S�+����|�Ay�;�Q���������ɳgOurS>��#��3tS����C�#�0���b�>j%�=�I.{���5`��Z�&4��W��ll���������!��G�cJ�<�֋輗��M� �?ٗ;w����_�����w�.�	�����ɗ�N�6H��K�hL^��إ����W��`�k&ڨ5*{�lH����ܺuS~��&����Gz���O�������)7�5�^$�Ot�������=ʨeNR��Ǿ�Vp}G2�ۇ9�ı.��L�s��\ν�����c9��צrf�B�]X5��C`��{�2c-C��톽"�g�(��:q�l���8ש�>�p�BHn|�V��3�>4��3��6�Dܾ��צH�((�A�v��u;po� �����/p�ǤX��e0�-�����+��+��+�e��ʮ�ʮ��D	{����Q �c���reA\�5 �ˌyq�b&��3k.e>�"�B��2㡯�Z0Q�ۛȍ��^��;/�ϩW��=��̄�|��� u��M���;�(�����`���%��o�L����̾|���|��GC��є��62�z-��à��}z�e��lN����33O;Fx��'÷�R��:�̠L��X�6�HQ��3���4$�����w;��ӂ�Vg%5�7L�5������`YƠ@��̎:�2Pj�A��8��-�T��:�� �;²�K����ܘ���t6F�|<ie���o����%}> ,9t�++,#�%��aԍ @	 -��CS�Ο��n%�jf��~e�(��ϵ�����m��L�#�#Ă�b�FVm�(��X��� ��.Hd�����ҷ�9<Jc��L��lP��i�Nb*�c�g�)!e�������sg�i�����4�X���3,˨D`jt��.h������<Ҳq-Hn�T�?�)�ą��X[��6�T׀�կ�+�6�I>�q&x%{P�`(m�7;d��f���G����>�R�$�C�ڐI'��R��!�d��Iwз��k��|���c�^���v�S*c{Y����C0��Ak86h{ռ� ���c������<D�b��D� 4Z�=y�G��y�����Q��O�ϞW�*Vr9=�htW�d�Œՙ�Fj=�#�%�dq�R^>��q�J���f��$�Cr|��Td�� Fj��'#/hl0h_� m�D�?��o�	8>�A�s��ё2�~������l�ZO�[�`'�gN"j�C�4_�r�ss/��2��?�M���������~���u-��I�-��uz�����m�G�RE}Y��REƴ�����)��i�� ��%�+�mlѤ���e�#�a v�ޞI����{Ŋ�ޛ�b����$l��C�G��Ѐ�$9���ΛթLm�D��@���ˬ��[G�M�{��{G�m�$4�Hai��l� ��F��?6-�\ڳ46�<+$�
�? �mK�]?�����w�Pn�{@�'�-�D��t����q�h��`\]���Dn߾+}�M��ӟ� u�{2ʇ�'�#Iu>�����Ͼ�!�s�����_�}�g ���L$�}������¼507k���X�jW
�$�&w�ޑ�w���_|������uO^�|)�|�k&@lֺ��>��eA�
�j�փ!A{����{�����!&��}|.�Zױ3������-�����	���q)�|���,���+g�r������y��d2�2ͳ�����Z�>�֭��7� ��S����:��`�ϯ �h?�3po\�!��G��@������A�������!��^��S�q�.ʵ��K��ɍ���~ �W#���C~O�s������W���Q��Zi-��?��u���?�3�u�M琷[^�X ؄Ć"c�LN����?������I2�R}	l7n`�H<��+��c��Wryu&��i�{}�5���Ǿ��DWw��5`Ējm��֒$����Jek��7$��v��)�:��Xw ?��<�����l����A�|� m��[�G��s��Ee��� _�{�����	�|K�����$���,N�uSK�T�/í|�%4��rk`��Q�� ٕ]ٕ]�c/; dWveWveW�`�z�I�M��  �A����8_LC`��8�z}gmf�0�D`�ιrR�@]��h� � �2�d<�û�qP-k�5ڸ�h�ۓ�dH]lhV�w���ܻw����s9?{mAw�G8��՜�# �_:�Y�v��_���Ӥ��(a�}��@p�z��ٞ0G�����ap����|�JE6#�q<v���]��u���A���,d2ٓ�p�����$S��u"_��O(>p��0e7VL��1�$���Ld������bA������i��ɶ�q�o��9���Qh K+%�@0����"��d�����$.P���ņA&�I���:^�@�W���@��<���� ����.x/XY�U�@ �Zy�%����j�=`{"20N�T,j1I@�@Z���d`2����N�3$Z rЀ��k�b�S�-vcӞ�X*�O�iP1(�g3�9���Q(�L�Qi=ҋ�g&s����x8�M���?��*�E47T�1�ARcs��p�_	'��(����Δ��}F�!��:��Z���x�Kcs@�äB���dA��@��a�G��J��>�q`,�����u8�0��X�3�N�����H�1�S�������y� x�����ij�`��t:G�-�!��KU�\�|�g���|,��X:�@�d q^:�-^ ���B^NE曅��������ytv1׷^j�]譼���_��g+��J簑�o�`�lt��:��%'�#!�y3�W��%�/���J��W��\K}yE?	���'�2�l���!a�P��	�gW�D���+99A�5$�2fb�B�_���%��(�������er �8�e��eg#A��x�'����Bp9�D�O��� P�`�W��<�I��[��]��)$�ZR�*��G���3�+6z=/�J'�!@@P`�d�+�?����6;���^�|]3�|=�ym��1�y��Iý}��e�(S��w��m�+H����?Le���l~�1M%��	��,n8�WZ�k�L� q�ؔ�<v���wbN����ڎ􌁆�K�~�J��Q-��>����y�-#��IzqJ$4��S��"��1|�e�X��ׯ�J����e�7#w�%�O/����������ҵ���X>�������]~���J�?���(���9�W0�PG��z1�H�0! �Ӷ�^�dL����t&]��C���䖼��G\�����ޠ�=]��}�#�ܓ��[����C��K]J�9�ҡ$ �H
nizb����>-��pŃ����t���w��0y���)*L�\�_�zMٶ:���$ �9p���/~�s���I.OO%�p�B��K���M��
��a'��6	'�W�dǇGr�}΀����w�<, 	u����*�X�9	4���׀A��@�Ș�Y�u�1�Z�kf�0���?M綾���zr��������/{o�%Iv]���3"���	���S��������^����(��\@�*�*3������>{�kYh�s��֊�����|�>{������_0P�i?��3��w	�3���p@�c�bQ6�h��X/�K�xq�=[��%��X'��)$Ǽ������'�7�?��$��Xq$��L��7qd`��ӹ�^W��o�������:�2��b��81�O���d�պK�	M�r<��\i�+ց�/�aB���]�s��e�<ca�������H�^���(Kc�v�[��ج��O�� ��~;�1E9G�m�����.~�u�ȝ%/|K�C�6�����ᑐ����4����M`ٱř��r�D�Ճ�Ky�:����-�m�ɡʡʡ�K( �P�P�P��¬�����T�`M�[K�Yd�BFb����k������,d#"X)���D�z�#�n��=���O�Dxc~dU�^�p0֯�����c��,C���0[�� $%V�_C��8���TG�5L.�3"��e�,@�6��y��@��th w4�"����>�n2�����U�����$���(�%3��a����x��H��S4�74��5�������[)]�;�T�:�}����f>
�@0C\&�ɂ
��i:`p�	�m��ܶ�V�Ӂ��J�e���`���s�7�tY�"��Ԗ���A7<[�\�)C���[��$�k�e8�l0l"f�; ���l_'��e�#>� "J~�m��\ ���\��A�@ȸ����ۢ����3����i@K���	P���yb�o5��2����u�t	����
CaЃY�K��錋��N���q�I�0X�YK\�^h���j�ɟY&4��gJ��Um�N��Ij���kJ���G��$B �h�$u 	�gȚ�m����s�� � !̢:w�'�yd���8}��|�,���j�Apm6��u
_�������h����5<3�-���i(o�6�QmI_SdZ���ui���8�t<���+ٕ��@���;�
�I#�V�ɉ/�O���s��)��9����H���I������z��$Ht�ɋ�3���v )Ⱥ�%J���{C��E@��L#�Mi9U�~� <�ڼ�Ŷ��	d׌%L.��]J��u���5�������^��˫#m3sj�;��V��Bf����}�˼"<��������Dґ��A)��k+c 8�X��[���] d1�
[̉�.Z/�)�a�w�=52߂!9����Pb��r���#]/����Y$�:3Cg 2��r��$���F���c�e~,aɳ%���HJH'n�P��B�K�$Y�uM����F2�����t>Q������:����Û�3���X�ƵL�������Y��_l^��R�t|j�5ڷO0�K��\���Rj�{b��ح�������:��r�^f��
�N���^����K�]�hL���A������_�����������ヶs!ã�4a0�����b�︖a@��\.>�\��97�8Ҝ�	��  +9_,u�����8^ �"Ե���5����X���k���|Kٴ~b��.�=x^ � ���J�X�IP%{� �̅l���e��q�@W0Z�Fb�����k����?��SZ�^m�6-���%��܂��@ȅa���6ޯw�ؙ��Wx�����RF{9Mt��4�m�uL�B�&{���ѱ��(r�%xf��?0J':n���g�W�W���?ʧ��L|2 � N�k���=tݱ�����|e�(�8ߍX.�_L&��5��`����ρ]�+�{.N/�{����ٟ����_�+9;=w%�7F��q_��$�D�:�*�gtσ:�Y���0�ւ�%Rp}��&�Ǖ��5���M�Ԗ7��;�7L o/�ؙ���ݦ   �g٫!�{W��gϱ�Dl� ��m�U\�~�mq��y���������r��|�L��آ�>c�����-`�:�/�Y�OCB�1pe߾������ =������P�P叮 �C9�C9�C�nK��
&�8��)���n�yp��[���/�?���~�&����-4�zb�)	���~o(�ј��0G�]�al>�I��h����(�^����ӌ�F ?F�1���O �~W����w�8����ײ�θz��|�i	)�3��3���}�&���¦7��PH{z��(%A�V���<��lNTUg�]�_�� �����c�ݱ/�9
 YJ2]Zc�8I�13�R�"2H
3�&����׆(֭d"p �p�.QGa,y�c��$�� �82��Uf�-n|��w�8�[���d4�O�l ;��A�#F
 ��|a��,�^"^���Tz�L�����e:�4�K g[V&k��Q!X�^�B��l����oW{��#�P V�u\�+	�����ғ{=|*�Ķp�4R̀2�57 1�e��6��}�}Z'��g	r�.P����)}SU���}~)۝Wa J������y�v8c^��#0����~d��q��^��^��'	�,P�{U'���8��4I�?�ο 0��fӱ��@c��3i2�:g�i� {��R��������o{ �i@�H��.yz�[3��%�P%i1o�d�ԍI_y��J]z/D�z+U��|��lt��ex���x(��k�G�%���}��4�{YN�ϥwzE��So.լ�����cf?�b�j-��l�_�w� ���k�x��/%�|�;���7����J�֔�F� �έ �e�l g�PD"�aW�O�L�m,�.A|�l��>�[������e����g2кp�@?���=&��WKx9߆�HR���L�^+����R.7���H$  ;Ԏ��~0Ԯ�J��KR�M�ŒA�z7�6�˨_��2Y�2y����G�u~�򵌡��s�O@x(�z��ß%��#��B�a��!��f��d��Rf����$`�J�3�6�<6���T���;d|�r��d��)�����O���t.�ߞ4:���(�n�t�N�'#�qڣ�O"@���� �ogV�L�K3H���� �S�y%�H��E�c*����nDWz����b���돸p�!nn�?��'�cm/�K ]t�up�i���B��ã��_�R~�_k]�>����W_�j�����~��yi0���q���єbs
F>�0K!o���ߙ����A��jE�� J:$+�i:�s"�>eo�P..6��\�!��$k�/`=�8O�� ~I��5��������x����w�
&�?��@�kE�sAL@&�,_��= r�����9��q�I$	`�}NN� �4Ȥ�9�3�!�\b����B|�g�����
x�aOB��wi�h\�{�K�9�!H��w0 C�>�J�=�/�>L�`�Ntvtt$�/^����.?��O���7�@�C�N���ky��;z��_��-N0��0#$� 0�]���x<�ёɀ�lky��y�@�J�x����{}��Ҧ�G�|�J�ӈ`b��o%Ow7�8��4�g������7�GZg`�D����ٗ��a+p ��m,H�1��K��38:&��t r��D4�n�=��4��U��e�K�y��N�Ҥ7d04�!���Q���H"�;g���o/�\���@����� @$pW;�k�k{'��=�VO�=`�=X��������-�Z��4�1){~�́oϳG`h���ƹ���\,v��y��)�P�P史 �C9�C9�C�Bge9 �LR�@���Z~������o~��կ~.�͆����A�`5[�b6Ӄ䚇(�	�@~t��S헫-eip��N��e[fo"��H�7�@���X�u���8+�T����!���j���f�l��0�3V��#��)�իRy�>���-�^!W`z�f�=�-���H�����ۚ�J�8�o�A\MA���܁��-��(��@ ���.���YE���m�ݡ{?cw��k��	΃�+�5���GYf��{y�)8�"�QQ¡u&�&UEfJi��=�BE A��_Л�Xx�d1Y�z�N�g��T��F4�M7���`�em�  ���Z���"�S��4��|M*J3u����Σ¤ ,���s�� ı"⎵���S�y��0�II��u���> ����f�1`P6�c�~pxGf:������j����3�o��'L��N�v����F4n�Z/�g�(RP?�C����~��K�����}������z��I<��CgF�X)�N����Bϐؐ�1�2��l!�6�_x~�<� X�Q&�g���+�-%K� ġO����]����0�>��b�#��F������A0�6ٚ�!��E9`���I��I@��;��]ɀ��"}.�3�B�l�}O�Z>�{"L����΁/�*�r)Y5�^��t��9q�?�\;J�r4к�H���)l<<at�b{'�嵬�7��\�8���7R�g��FH���	NE+~��/�����bSj��hn�o�`�8�D���8X�͒����$�W����#�[$��Ճ<�]Ӑ��8�,Њi���Xg����Σ�|�!� ��������Xr�u(�YF/�8H	9���h�O�7>�����9��H�y�N����2{�{6��ݻ/��ÓLN&������I?ѹF�h/�^{�4ͦN���me�鳑F���SɛL�2��h�I�	�4i�i_�'�R�<�]�nt���J�{��Lή���J�!b�@���sׅ���F���쟲5ߡn�������y�5_3��u�7�Q��%��C���0�3��E�5F�Bϓ����������H��c����ɧ������?�o��L&'rq�B��ǔ���@��j-__�l���od�}��gߓ���_���k��?�W�V�5gpv +	�=2��I��]�� �P���^>��32G���<�c��2���g�8��h<a?�psGf*�u��/�^��>}õ��?�g�O��?���A��L_���%b�i�O�;�d9,"���I��\�g���3�XP���Km{x��N�H�?�߯�3����7̚Nj�q�?� R4ޞM��9@���\Dn>Fp0�:VAHJ!������limF��Y��;�A��&Lh�ƺw:b��9^�zE���Syy�J.^����Z�>;�?����o�1�A�WH\�y��}Ǌ��*���z�"���{�u~y��a�M��J��ŋr�s7�����N�R����N���k�)
�����A[��"��Ұ�y:9`��ֵ2v�`H���}j[���d��i�̏�����~d�,I_ ���w	�'n=sQ`GZr������?�+�d�� ���Ƕ�tD`bJmRXx�0t2���?�1��<Q����5&v+�7�1�},U>*�~����)3�D#�t�:�C9�C��P ȡʡʡ|��T���$e&aړ��k��ŏo���vI�
�``���xD6!Xq��-��Cnc:ӋwJG��v���e[�|�ͦ�F?�ø��Ң��@�ʝ�1�;��\\^��>�����Ћ�yi���(yU�6��v�փ{_̧��j�B��2c��@�u��QyI�ӓSf��7kg�ʎ�ݍ1%�9�A� $���7�y��C��W��!���;³�vAf�C�.�`X�`	
��<#�@<�H��WK�/�q�f=0¼�)�;Z64��djZ��!�Ŷ�tT@6��6��~��� P���� u������?P0B��A5b ��fx=�d8��Ӏ;�ϐ&�)�X%$�R�����L��Yfc��u��-;�	P ��P��U�����Oɬ���ۺbp,
 "�>�]/w^3�@)
��� ��0~�����c;�̂��~<��}�'
^Ri����X�X9m�~lF�u'!� v��L�A�3W�r"�������}1n(�B�GX!c!&���[�[�K�����ѽQz�ұ}��X�2΁U��},�(
}#
�}З���x��7���TJ���1N�0kÚ �e�J���YJIrn� 7�M\��4�a�'����, \�[�0��ʇ���2��QUc�9!�ג��}����!�YA��=�wd
���y$��P�3�N����lW��j1���'�&`��g/z⧾�JdÎe8L)G/�����_�b�;٬ne��r~v.×��Z���ndW������F�|K�����y�ܘ���1P=h�ޗ*_s���Jx!�g����D����qX]/��sd&�`(Q?������Ƥ��	��FZ���1�d�`Z+t̷����Xg:�W��jF�//t���BJtq��P7���k ��V�@��J�r��}��=����% �
����II����'�qA0m�7�:������9��E �z��9׺��Vw�w�O��+٬Y<�ܪ�GZO��I��3m$�ACk��e�
����Ɉ��p�I��t��ϩ�ڕ�7z`{ YOz�yc!@�i�>exe��BJz�P� =D���rY>�~'��H�86��1Mch+:���w~zJx\��S�����~W����㑜��K̕���D�*�00/B���'�ɟ��G���'�W��'�����/y�θ��Y���5C����z�Os l�o r�]�ʀ�Zm�q:g�Rs`���?�:L��-�\.�d�>pvv"?��ˏ��G���k����\�)W	���	�vzh`>v^��DzQ*:�%	��%헜'|��A"�uL`"-$��e���A|���� ,��>��ۜ�z��1���c�+d#-���=	������{�m�dn8\�ػX~g����X����B��4���8??�K�g���x|D���:�F#��0f7��[qX�^�N�����������ޑ�����'T��t�w���#	��Q�&����4����L�F:��` \��s��U�}[Q����y������-�`H�h�gy���;���Ԙ�;�< ?�⾭i��s���A�k��'K��fK�Rh�aOb/t��L���~�1�c?F�>��d��X�!�'Nm�+�+ݳ@>*��W�7������5��a?�Ħ��_�݂j�%�&� ��I������}�p�7� F�$mj�U�������2j�O����C�e
�g���4��P�P只 �C9�C9�C����a���r�x1{2��������%�������0-{��BoAʭī��3��Al�8ev/��B޽{����6o65oq�� #�3�p����vA��L\��Yz����m����;�w}}�,WV���O�?�C�T"=��2���d9��6ό%�n���;�| ��0@p߲C}�}ǚ@���.��3���a ��"8H��Ph@�;��|�󁖁��� �rH� op����iѤ�J��>��Jg�ɌS�Ơ$C08M�/�5�tG��d��-e�,��LW�`��aٌ��;WN��  Y��Р���c��{Mnf�/����ܝRaaa���}�p��m�rWI^��cH��}B��4ɮjT@��0�w�S���i�����@��t�S>S8C�M�T#�m���x�8�U���dW�YPOxF�1�����P� 0�I�P
	}�6���a��X�o����ᵨf�0��.��Ǧ��@P�����g�V������q��� ��j�� ���9 E��$�k���>JI��gv��`��θ����?j_ �����C_.���O>�ˋ�(X.f�0ÈF��*���Ɨ�õ��� ֶ�˥�c�i+!O�؎�hm�c1��թ�AV���x�^����K�0���OR�'l��YK\'��)�Y�rq'���dv�Y�?�bw-�h`�[fRl�D��suD?� ]��h�/P�.���`0�e�>�ڍuN�#��
S�<�T^�29�D�x�,�T>�l�?���	�^҄�(j�%R��Ja�^�P��wCi˵d˩�o$��Η[٠-�&�����W2���"��< 
D�Hk�]/%_܋��k=��ke�ۊ����
�'ZEW��rq1�6�e�����>�&�u�\I���D�U)U��uv��;)�$h��>3��/t��^�	)��k,t?��?N�jp"/ sQ4��A��OR�3��;���Z�=X�gk�o,��r���$t��]s����0�j���h[��e�`%��1�0#1�-�!��}(��)$+I�c؀�H� �ߌs8����j��/@��I�PA��Oh�X��˗����\�t�[�u	��͒U��F?�GQ�L
(�$T�J�	��!���xO��w#�  ���uEPғ��D�j3���C�r���uvv!�����w���0��#ZO��8�B �����,P�k�K�ߔ	%0��'�m���6��� *poM^�>Pgd�Ėok�%v��>�=�+�)��$(��D����l4��q�M;m;�l���)?� ���6��Y>��ؠ��^J���sm; N @^�06K�$�IL�	F��Y<=ʯ�K�ۿ��������(�x� �(�s!I	���>b��q�	�Ľ��,���؍���Z�d����_�������q��l2��� 3���=�y�� �)m?������ˁd��z%�*��p�	�n]Ŕ%�K
�7�Q
��@Ƕm��Q�8����W���
�����;`ŀy&�h_ʲg�����3�=��N��I�>KU>?�o����w���7e���?�����X�{ �A��A��S���7��J�P�P�_V9  �r(�r(����B3������
�C?y���E���X�w�dѧ�!%��B��i�������$�sb�r@u�d�����B�t�Qz��e�Z�����=����w4��ٱ��u��f�3�`:��7o^�k��N8� 	̈�K��k�9	�S=��ݮ��� �^�@�2�vg]	��� �� F̀��QG�)� <B:��/����u�.�R�YͫC�%t�s�֛�d��i��j��޲����Խ�i��>Y�ue��w�<�h�d ��g�N��d���`}�p��������; �k��R:��>3{�I�� �Q��M1=�ИZXd"Z��C��x��II+��+�Ѱ����y�,3��iuA|��^C�.�Ѯ����&-T9�( �N��t-0˱(-8���,��IG����I��;��po���8���d���`�l8V�1�yR7�����b�V��h�^1��Y�e���8��X|5��suP�����_[���W�|�c?�7j�yX�(�D��\ӌٽ���L��*H�>��@���]��pŬOqF�{c�@�1Ι�A��W/�G?��\]]Q>,v �[��`�0rq~*o.��/��
-~�1TH����FC�%#f�0�-(���ّ_H�Y�s�|�b�(�X�������D�H+^2��8����T�YO��Xz�1���T��{�-�I���A�(�(�g�e���@�r�9�/��+ن���Ti�m�mX��o�r�0�N��Pܠ�Z{!�,8��O����Hz�Od���\[���?{#2C̱���%@(��l���D2ɬ0�Ѿ<Ҿ�&H>�F��V�t�)�T�'����#Н�%�$�#;y���,����+�=}!���������\�:o� �����z#�gzm��d��=�6�����)|��I��z��r��J��~���l���Z��\�v.��Zݰ��V$ fE��q��kl� LX�dv�{��?�&�R�k}��D^-�C d�*S�c���!5�Vk}�	��>����"��g�;Ġ!#��H:qk��%��3�����L��B�rgg�ru�LĚkAM�8����B>d�b3���m�.X�B/�SJR! N�! e�7�`^-�L��ɲ�%?�1���u\	�L����^;"{�V�l���״:�dm X����̱�������?��?s~;�����+�ϗ\���ꤍZJF��ވ��~2��H�hF�렾��1��X?Q_�uF����r-k�� |���`0�ٔ�7���mh�80um�  �a4I�s] �����& o2�؟4����M�$�|����
����c�t��8̝>��d��������O��_��_�J�O���yw�?��`�^Sn���X�D�3�e0�ԥ���������{�Ͷ�x�����lu�N������|���YO��?���DbH�dǊ���F���*�]JǸ��V'�i�����6��Vu�l
$}HaRN�򝌚�O��H�0y�9��$S�"v]z���C�3������M��Xs(�W?����gϐ��()uO��g9/.�nY�}���g���n����s�}~�����YB�5<[��q�c�v��%Ҡ��}!6}L0� u:�C9�C9�?�r @�P�P�;-�#�Ļ�N&i���WH$ ۂ�=�!�=+v�mg<	�����vhC�bKZ�z�]����:�[��4o|� �_�fUH��yz����{�Q���7/_ʨÀ�(���V˵<<<RV���+y���&��>Bk�w3;���6ӄ�]�q4��C�&̥�K�2̼�uf�ֻ����4�t�,-0�$��=z�� ����R;�dvvY���$1,8�e�Wd��`,tA e�n��C�oz��$�m��u�� ��� �F��#Bl��9IV@�7@G�!x��.���@�/x�0k3նX0 ��C�x� �_	�1Љ>)�l-�T����׻�5Ş����GS��(�`qtܾ�-V�3`m�s��Ҁ m'�$�X�@@[��Ken��~���ai> ?��1�O��f�� ��?�~��a��f��^��rm���9�U�^�s���@�96P�AC�0Ȋ�b�&��/��ʨ]� @���i�??
�>��1:�ɜ�:�|g�� ��ޚ�G���4�@(1���
�ɮ�G'���Z�*Sf�^��e;��~�A�#�m����@9�h��!s�-c�	��g)3}��Z�0[m���^�u&��D.�=9�x�sX&Ųf��Kq�z���ꢯ���]����H���a�m'��	[�Wx�d8	00�	������u�R�k�EϠj����K���1��	����[��Z泷���^�z���v};�:I2�������`Oke׀�O� ���ِ60���uRk��G�E-=�r"?�D��6v�Sq��2�-8	}�Ois�{c	ҔsE�[�zvC�g���?�K>�e;�?y�sH�;�K��vF�0UO����5��o����$��J^L������R�� @������x�J�L�L�R0k��:�����\��� #%s�E��ӹ'�y_e�@*���t�ǜˣp��˃�3O��>C�0�>�6�=丄w��'W�ٽ�����?���������G�ژ��}��L��o`�o�T�v@�dM�'�K����;�b@i"1}�>h˹_�($v@y��3�@Û�
X��hH���`�F��N_�]@)�X�|�{�`����|&�̻�{�x���q�|�Џ8���LH2��u���k�9�s����8�Sd��XB�.�A��Qll	$`>h��oo����F�#y��S��Ílt^�B��uh P������ǁ�q�zCIL<;�xg�{1�4�x�� ;�߿'#u�\��������K�7�_�-��G��{���Lڪ),@�K`�@?&�se�-�#%�r�N`��2�!�=&�cx� k�m����\��V�<�v����u;]��}��|���e:�rn���$�ʚ�kK]G�ʙ����[�w��|6�3�<�7����#p@�f����2{��_��� Y3$����3&� _���P5���G�<I��3���?�D�i�V�=�k}n��� ��D�bGvqL?� Rn�˥%�p��$�� /6� �ڽϕ��~�����~k�[�}�t=�
�#v��VԱN�]�ɭ��r�?����g�Ҁ] �h��)F��wk��At�s��nj�yλ�d-C��d}|����5�>J��}2IW��������)�r(�r(���[ ȡʡʡ|g�¢�6��N�b6�Q���─�r����G�-Vz@�Sb����˚R��������d�^;c�T� �Y�z�Z���<����<>M� �[r�á��}*��'����aYmДFAb�j�˻�od1}�=�FC=��ԕ�����\���k�͗R�vr}}�l�m���PpZ�z����/_��_}�5�h�/6i����OL #`�65����M�Yz-�-���P��+���Р�;$���l,Ȗ�Y,B��"���D � ?Ɇ��l�Cl�Ara�N&M+�9�!e}��� r�G#�KάȊّ8�C��n����Vf@�B�Y�8���S���N]~}^#x����4��`h�ߐ_�,������o���)�V�(�)ZX� >��(�g�{@�>f@[xj�!��?��CzgX &�5N�{�@Hi��h(�i/�S����,��� J�r�w�P�o
������CD򝑩�|ʩ5��_}�	�4]6&���k鞣gRP��H)V�f���G�`VX�(�� wF��\߫}l|� ��ݣ�Ӱ��ۙ��"�%P:���^�>�I�Є}�e���J���$�ĀJ���4����e�9�3jE;�b�D����3?�Wa��D�{e���=7M}��a��D39%k_������|>g�̷���3����姯��I ��#m��ݐ�9>Pl���e0^�zy���Չ~4�TO��l��$�dtDN�e����	��3�{Z���2��ZqǓ#���粺+ӛ�%l�ryHr%ն������|&:th0�6O +���z�\���d*rtD�`K��D�J���Y��+��� =��8Apt'ӧk��Nƃ�����,��@�V�d�B_�3i<L2�w��0n�c���i�݋�x��v2E����/$�ET�%g��n$���ԇ)��T�@j��5'��Z�����f��x%�0O:6Vzo��#&j� ��!���Hr�z���Ծ��d��:�/��![�����dө�`V.A� ~��>c�Ċ�ˀF͐lʭ<|��ܯ��\�f|��ZG�����[�����	���kE�Y���ky�����O����G����	�� f�0P���xOh��b$�rFרɼ�8��5y,]�u����=I<༂�u, ����_��� `iB _�ْ@t����Z�3�1�Q�H2�G�f+�	�G�@�y��~��m��y,���{���gV���A۬�rg�6֫V?A| �#�?`}Ce�R�ΆbWڷFrvr�שh&  �8�CI��e�@��g�Ð~Z;΋g/L�J?��#@���;��߼+?�៘�����i���&�r�€q���p��{��Rf��|x��l��Y�T���K�͋�Sn�W���|��[��9���!��߾{/�����$� ����A��%�?NN�>$���m��*O�~R^�R;���g]'zq�=J��R��6i�=Hܣ���n;�iNN�t�g�W�S�t(@_Ȯm"z`�Z�p����?��<�uLƾ$M��mV�|`Rl�N4��ZS�4ӱߙ��k��D�F��� � �m0�׾���)H��|x+���/u�7�8�0�d���O(5F��.gX<�uz]�u���<5�Iny&+�s>$X='A�8��= ��a)�۱�j���J����j���I�� �&�	�
[�t�g�,���U�>�L�*���.v��GId���眉&�C@rf?[m��R�ϑ�KYЋ����8l\���el��XN���$H����`!e4�	�6I��>�=X��]����nV�P�b�G��Ʀ��&%8��Cj{AnU7>~[���C9�C9�C��/ �P�P�P����7�����ʐ��'���C'wD���m������r�.����;]ir=8��u�43��Y7f8�L���qH.rH�1��(���`	Xp�׳��b���z��'�zHF��9�!(����2�2r��"�������G���\P���&痗�у�����(8��e�m�b�!՟�B"�I(5���ܡY��Kh�o�0�Cv��h�C&�[��R�N#٤v ��C�9�������[���-�����qrRC�J�*�mc��1]��(٠�Q�T����3��S���w^�f�1�`�� [*x� ����t��%���vC#`d�Z�%�x<@��L�|@|� #�d�������o���b;�[*%c����˴������	f0����^�ȁB_�3XU��{�=L��l� ��&��e-���Ϧ� �|g�ځ4PE�Y��[A@�v�#.S]�Y�alu���&BЋxE�n�;��x��~#�Jg���}�ƯϚ�vmρ!���}�=lP�k�:��; 4���#>���o?C&f<r�1��+�8�ނ�c�<B� N&�fY�;h���9|i���;g����'_����p"�㾌�:�z���XpE�9�� 7�n�>XH����i�{fȋe���.} ����r��$�Ń_�}�;�w��g4$�t��>]�vz��i#��P';wÑ�	��e�sX���2���L�r � ���k�ފ�C����yI_3�X���VSJxy�B�F� Y]�d5����[IF�R�5�E�@[�W�4�@�Y�e9�:�=�{ZQ4����(����Y*�Z�x�xk��I ��RK�W�ę/��{Y�������+����2K`���Nס\�Nu,��O��e�<ږ��(��/���d�p��}	`�����Rne�}��s�@v:�ӭ�e�[�>��=�z��[J_�ˍ<}���T�k��T�IJ��d�Fv뙮}���$����AVO�����g���h<�9�킣���%�m�&s��٣ԝ{����5<c��C�K�3(�m�e^7��Ǒ��1`P�n1����ߕ��w���Y�����σ�������Q�GG:���2�͍���{�G)<�J���:�0G. >���Q.1ѵ��'�A��{.!+�]bL���2�̨Y�[�<#z~'��p�ǔ ��C����}D���6�����7/�7������z�$`8����sd +��#K �`����O|�F��������b�5p#���o�_B������A��l��3���o�~/��� ���s��w_�g|��%����E�bM�zN�d��\ۮ���C���޽��K�}�ץ�t���eB=�uJ`ׅܟ �Ŷ���4Hea]B`�7iH��t�j�y���W_29�oX�H�XyA�Hn*sq+��zxU '���<�`u�~ �,��֠�jk��&L<<�ʻw_���d/�cߊ=�NׂT��
Ҥ��;C����<��M3�mõ����Ϩ�Vm�b�?a�h�g�t�g�Uh?3�	ls��+�a	��g`����������,Ÿ���}��B�����G:n�w.�}4��A/��{i���bm�Z����G�O��ā*�$�����^��������ރ `ζ�I����3tQ k�Y,��`WC�ܲu:�8HD6ɿ������r(�r(�r(|� �ʡʡ�wV<�k��k|ϧP ΄~۶q�c��NP�,�at_��N� ���z��Ԑ6�t"���-�f^��X�L��t����Ձ��ܱDD��b������M ;@���E0���1�=����(��3J_���2�4�t�R�,{~~���j���r!�ە���>�Vf�)��_�!{��K�ܤ*J����e���������Ρ|�E�����k�9��@>�j=�gԤ�(�F��|s�Eq�Q�E����#�n:��w�l���=������e5�`nr>�(u`��!��G��A 3n��!��/�Kc� @�<G�`�NQ{���2�s�yo�F6 � �g:�`}8g��Ӏ:D�a`&��1�$�/�WN���B���8#R����w��=�=K*'?�z��L��`�&���?��[B���Ih=�z�I�>2M5I2x����7ȼ5�[c� #�u`}]�Ҽ9�{��rݸe`�SM��8	�#C��@oZ�Вokj{d3 ��1��"�z��K��t�g�����d�T��5�`�o�"ȔE�̭��"�8��ˀ7Ę 5A4�}u���1�z�A^.@z�$wrf�3Lz��s!8�����^=軐;Bk"�v49���XF�Dz�J�(�?u�W�ZudH���T��	�9	��S>.�r�Z����A륕��ģ�S��(��N�@�R��-�E��
��ox0��^u� `��>t�z�q�d�e8)�x��$|/���m�sjQR�/S3>oV�VKkK��4�"�k�}!�٭�÷2<��`�Pl�(,��2�g�%��n����	=�z���хT9��я Mq#��:g�C�?-�O29��I2�5#}$�k3[�ݻ�̊���A(��+�{:GC�	�~Ŀv2��ʉl�G�IC�] �=���km'��:�7���;�6�[���Ò�~�X��y �H�f��������TY�[��f.��f�N"G�V�*#�J�؏%)Y� ߶�X�+������=�0.�dˠׁ{�����i�jj�б9\����<:seJ��hF0�����t_�{�2�|�;+���d�(����ڟ#�c{��d�kc��gj=�ᕀ�*����,[�,#�u`�-S�V|�|
��%}d�IP-��g�)��X�����H>h���� ���<�0��m�83@�5��W����y��!��vr������M���/Ю;���)��pK��$�3��'�_�H�N�d��9�_H��w���k���?���|��A�����������Hf��~��\�~������F^\^�~�N�q���V�;\�i<���_s0u��9:�1��D����Rj�d�[C���`�\���T���������ܣ���I�fO:��3��ħ9�K&@�������M�ϗ��l�֚4�!�������5�C<������_�<Sq=�L�$��s��1X�ߕ�[�������"0��g�YEϞS-��G��o 
��cw���׭���β�k��,Z�$٬2�GL����(JF����i��.��0Q`��n��Mנ$�	&N�=]&� �}�i6�ղ� �tTmF�=��4N�����D2�g?5�!E��y������z�c�¯��KB&+�;�)��/(�v�d�����!p�Gr(�r(�r(�2� 9�C9�C9�הּ�葠�sR�����^��ƽ�l�\ʹL)�"c����Yd�e��([΃ш��8@U���YbVug8izň�g�� �T6^#�Y0]0�a��^2
�O���'���>�a+���|n~�4�k�s�w���D��Y�9�d��zQh1�I@���p$�ɱ$~@Ce�Ty|x�EY��Ȫ�#j,���;SM 7�|�
��-K�f�A�.0�IE!�Ksj�"4>Ҏ���dH�黦�L	�ޠ�XhJ3@o���v��4|M�Q�K������@��BU1Ɉ�1(�P[]�a��c��T���Ȃ����*<)��o����$3ST��]���P�li�(�N)�+E���<�:X���V��c�����~���`�C}ǐ	(B ����̕.�O���e���#@C��T�]ˊM[��:#���s����X5c�������}T���q'tuAO����o��1;>V>��_w��[�����;���&�E`�����Mެq쏎�S9)���h�[�B�۵��0�$�M���2$p����XA`cc�����Fږ~e�32z��2o�R����x ���7h����9��4?�"�6�����w��#t���h٘�J�ɧRe$��VҠO������:�>m�i
?�3�x�F�A(��Q���h�is$�1ƛ馃�P�!%(rt���c&��\�m%�/i|.U��q���Da�c.���{k6z��$ 8u��&X=�=/�G�2Y�)[��wK26w�e���d|)��L��̴��m&e�cy{/^q-�d+W/�2H4�Ot>ѹ���\���?I6������FF��i}_z:��
���T��?���$R�X��:�Fp#3[F>d�z�ӍrfA.�I��H?k�)����P�	�Lq����<9��Q��~+�7�&���!�~�(������R�*��@l��e9�	�G9=*$��G?�����3����z����t��8�ۀ~7dlղge�E��G�1�q�0Il��/���������DomM� �B쇷�b��� ���h`�	�.��Q];|�U���{���Ã����,�N������9~���m�q,�/i8I��5�[0(6�C2���5PP#X	��3�d����pHh�`2�\@PX�ད��)���@�������d����w2>�u�/��V�k�6�lH����������٘?|�8�u��|H}��A�K��f�)�E��L�?�D�R�c,�5��������Dz���n��HBeщ ~��͙ow��n=�}c�r�v��~_��������d@@�jLR��xV�����
�\II-2!喘�L��;�i����Ȓ�: �$=���Zh@�Y~�ͽql@�F�`���5=I._\���%������vY�g�}C����A�VlO����5����f�g��v��n�dτt�����~�'��a�����b����C�J���7�r^3"*Sq\��dk\�π� �y�{��rȢ�ᨯ�����1�l�<�c�WW����Dc���3kd�#��]���ns/c�%�3�ް�k]V
�3����8���~�uI5�y5�x�؛5���s2�N�`O����߱��|��r(�r(�r(�� �ʡʡ�wV��Y4A���t]W�6
�B�
��п�vW��r��$=)�!5=|=�Vz����P����D2�&���hl  %����e�`$5*G��=��e�k�EE-\�z��_�.]^�����B� �eQ���Q�G��{����pr:�����i"�Wk�GzH�Oe5�1�r2�����y��Ϡ=M/�|�Bjƚb ��8̛wC�()a��>C�>�`�2&��5�f��@m���zH�������)�8��>����N���������uR�0�{)�~:�vp��$�M]��B|d�� | ����Af/�Էq����@@��2�.(/��(rL�Z=��Di�}�H�����+�����Ȍ���;����X��Ii$.��c� BA�L҈��X����m���m ������(4M*J�t�]Y�Irծ�!)�"�}��"-4��H6�Y>���p��>#��p����d�����vM��Bjca0�ق��)�~"d�V�hJ�ȳ�za����+�N�;�����ع�]f.�� L���>�Re��Ƹk���#���K��ڌp�	H�����W �	���a_af���"��#; rf��L�&`�|U�ܔ׮$h��D�� 1�7�f#�|-��夦�+)����x#�_J_��iB�f�!�A[r��Zh�_ï\��@�+��~棬f��@���^(?B/��x��j����F|H��8L(���$i�KV:�����$�r��G�5��L��F}�(����U�IR.�M���)�V��^jo��OiC B�qm��|[��6���z_m,�C}+-�AR��h�z}G$�h����Z�:��fP� lUJ����2��W��16�P��T�m �ǜ�N�h��"Z/;�ˍ���c`�����lW�f]���B6+�u����yz��=���3	���.2�e��=h%����$�k�sU�5  tk�Ch��56dg2L�<0�|cI�{@ā٭I�1��8�\�z'E(���[�@(�q"�ɑ#���{�5,�T��L��5-�I����5��$�qsp0Ӑ ���t*��)��s�����$�l=�?qmp�R7?1 ��⡁c�@"�k�1�>���j�WL� ���!������j�@�zߛ�Jb]�Q�0�h?;;����R�:�'W���H^K@@�>
\�׺µ��5l���<5�hxXY�����mv�Խ�t�����2���3�5�9WE������B�ͦ✏q�pw�s�qx -癶_�����+7�R�P+�l?�1*���M��݇{駎���G�<���&9f�X>�qZ����E;�\��{ 3�^��\��DB�N��&�8)���� ���w|:"#	�x�^D�\����O�rӿ�m�ɓf���1���3��{3���&E�m�P�\�l�zE�O]�}��	��-[����,*�E�:n�>����kJE�$���ul�%����j��|�taz�۠�sJ����Ĥ)}c�b[f	��ya��V�F)���&cY�6:Gnd>_�S�Y���=���$0��!ӣc�
� k�s��M�9���٩�ǽ%�e�	л6a�)�vڬ�����$��P�P�� r(�r(�r(�Y)�6��fU6���Ve�˽8��*��^?��f�`$�_c��2{z2��:�Ho4"���qd�z�돆���}:CV���ԍ˶�k'FM? `�=β"�E�Yԝ�kŌKHqm7+j���:$��������/d����H����Rί^H2��u�&�����Q~��_��q.G�Ԥ��g�oj��ctn��L}4��RJ#R��*�u�X
&! fV�d������	8SR�,����2���� �lL�!��c�@��ϝ�B��;�����<��N��	;|�ބl��z�v�_��șq�o&G�l�S��V�˾�l��F�6촤��Ueπv*w3{�yk07x1�~f�݁�Y�=�/�A��ߎ5c���A�,˵?�:?�G�r+N��A<'b>ƨ��6�P9�L `�&�suN�%'O室�c�M�90��*g�c��� HJ��T T���6bp��B>���������xc�Ƈt�V�2ynJ�9�u 9R��4DE���A�vc�}�����f�]�y~Ա�HC� ����>c�|,; �Z]@��� ��]�1p��g�5s�c��{ ���ҩ+�Q�;�.� ���al'�Z@��I�#�����Kd�}����́e��ة�a����3�[< �kf��ŒL�][y}{2<�����d���Ӈ{�кx�B^����h����(y;��BbY뛶�Ҏe8I$�g����1���B��G�Q�����xh�[s)�L�È H[�hJ�x1e�hF@��h�6���D}�9{��ޣQ-����2��kvZ}��a_����5��f-���y6���� h�u>{�����[�ϳZ&�����_� _pM����42HaN���N3��$��*�	��kJ��l�k}�[9�^
S��D6�Z��?	0��I����ˡ��.$�� ��x���Tdz�	HH�D��B����v&e���"��Ѷߍ����L���v�}cm���0���'@Q����n��9YI�U����O�$��<ǘ�R�/�<��c��_��ˁԸ>�p��Z��q�AR���"������dQ �&����M�ڧI� 2��0
��� �`}�z�X-�����k"�Jm]O0�5h~SXı�|���G��w+u_qtrL�#��h4��3�NCF�!��2�O�)��O?����Y^z����3Dl�KX;���F��h8�|1�ٮd.�|`fϨ��r��_h��r����j߄���n���''�b�{{:��g�k�{�^P�^dY2�!�sa�5N(��y�x<��r�1�J%5�\l�RL��MlhR���h��!�=I����OtnLu�,��O�9_;��ρ�%Xz��@!�]�9��u@?�� ��{���z���Ix���]�-���6��)�A�(Ju^���XA�����RcP���Ji�4e� �%�{-�h`"�W��D6K]y��{�E���PL�
��:��K�G`[�%;@�>뷨�M���*��0�}�y�l͓����%N>s�kl��M��ٜ�2$���
�$���\>��o��suy%��R�������`��i>m^K���tdcY��v&�1}�P��A�s
�W�����Q� ��aP�|g�܏c�Cwѯ3ݫL�}����n�s(�r(�r(�� �ʡʡ�wV~��o���/_��޺.6�(L�zHz�:>�pM�xȘJ�Z�~D�GG�\�ՋKf�/�K��/���A���Ymײ\�\���!�ev�@�0ٳpb��5-\!{1$2�nL9�����e�w6�j-d?KC[��K^5��<�v'#=x��T^)[�y�4����k�o����3���(A����z����y х .O��Nf��CX@�r�����d�|~��@d06�p���d�h���@ZW������3����s�5=���eUR�A�`ܔ��,��)���)��0n웮�����9�/�
L����g�`�?p��,���5�?� 	��}A�ɱJ�	{N��c}N����vY���C�3�5�����S�f��}oa�3wz�ẗ.ձl��^�>�뿔m��@�1����Qe�g�G���<4?i�ZK�3�(���2�p�l����[����e��I�p\@��)�AaRN��\J-h�?�0��ρ��,
� ����}h�褫��Q/]}�:�svt7v�Q~08��;&N���|Z�>���H��a��wrnx���5\��K�E,���겝[��Xj�R�`ړ��fs�q�Xm`+��(h�%�u�"��@w^ Z �3si�}�>��j��Z�'��BUp�LYi7��MR!�;�����!�4���S���1Z��$�+� ��u����ҿ����%�����F�L���]�87�-dɞ����5�y��_���w�� H��6^H,%������(��'ڶ�����X?:����1Q2��0�y�$5a���o �f���t�݊�ꀙ���{y|�@���ѕuΝ�%�8@��X��@0�8|��7B�$�d�oe�6���O��f2�_��1/hD':��Od��AK��2@�93ԵB | Ӯ�����| 8w+�~�eV����|,gG)��^w��=F,?֪ø�<�� ��ff��A@��  �^��M^�5�^�:����	�sM���y	 Щ���`���	)��h ��1G����䕼��� r�2#�m��_�Ȫ�?�a�̷gO��������<==�/~�2��g�{o�+Kv]��s����W3�X$E�� �a�����_0��F�,زZ6HI$U�*�����sFdd�k�yo���%�y
��{y3#O�8�^{���ɹw��z�����<�A�ձ$�|H��;rtph�W���` Z���2��w���9���hC)ʳ�y��}�dk�����c�f@�C�m]�C����z����c�_�I�{��VJm�꼜�2�cɌ�g7ݷHB���zv�Y!�K �AD� i���C���M3�b0Q�6�i�ݢA{K��O��[����s�rL�����Z9��II0���(Hra>P0���bC�׍t��g:����������'�锾E��K �*'���q�>�;�*�X/��C����ho?�d�|�;f|<�����ѣG�?[����j�-����.oX����~���k,�&1���%�D�dR8�0t=��d�]z��vo�~H٬���g��o�<� ��U������tCp˼�7�ȹ�3}([��0���KL���7��4A	K:*��o�]�odrs%�d)����A��VO�v��S��t�&ΔyZz-x���z��M�A8�-q�,�v���d�@H�{bH����`C�5� �rz�����+�'�'o�s�ݕ]ٕ]ٕ?�@veWveWv�-������/�V7�U�hV��>�)���%�(a��e�����/��/�/��/	|�ŗ������3�փ9��	����7��l�`nۤk�P:�rH7o�Ibܕ^�ϬM�^�C������V̴���� ��h4d@�*�0(F!��C�Au��Wc9}�Fn.�id-e/�/� y-��PV�r|t,��ݓ�N���\�?{f8z8m�k�b�? ym�0����ܙf#@�e�ˎ/X��b�@TD�vY�u��J�),x�`F�,e6K�.�V�ۂ%��r����;=G|Iҵ�Y� ���qAfR�Xj~�D���	XV����h83�(b�Q�d��+��0o�4_�M`���C��g��A�~�:��R3��^ r��� ��֟Bpݗ�AM 25�0_բS0W.C3sϜ�I�&��k'�h��P�	��xX��� �Q�-&k"YX���5�����lI�z!C��6��o����%ɭ��6���I���l���ñ.�%��1�Ϯ`̋�G�W����{Z .�O@d�=����Ay�鑗�n��m��/��0Nl<���v� ��s�Ҭ�6̤����H
)! c���Ӌ �-yȌm�O���A�m�r{Ș��{1 ]��C����y),@Z'�Lv�*qAp�׹K
�m�W!�G&)H�c���mh��R=I2����:7��A����Kk0��ݳչw�3c"��Q���e�LN&MJ�N2�)Kt����H�b������:���1��]��3��S��D>$�:���@�8d	α�1ӿ��T��r�Y"�k��DIO�fζ��� j���Z@4�6i���������H�����ѽ=�%n!��_��V�`�/_,�\�/�OZ�0�����J�XW�:O��D���t:MI�R:U"��-���m��u�����It�7����~�䑾���,3��,��B����B��9� �y��u��c	�����/L:3R��M�*���@�Iր=٬L��4�� ����b��ͩk�R" [�=d7���Ȱו��>���c�g�!��@�L�-m��א
�<�DZ���c`�bOt0Ն��T.�/��K�)	I#4fe�2���+���MFþ<~��^\ ;� hݧF[���uZ�.A�~,����=#�W���/S�a}��	־n�ìv߱��p�k��Q�@F3 �d�����I��x�3�+�He9�n��z~��pӥ�����5f�{,��b��Zl�I��K�I�K�I�{��4���9}-k�_s��00$�D
�Z ��^@:���	��]�?{.�o�P�y||,= ��G/���m�ϣ7�qO��c?ts}#���d�`~�++���֟:�!�2h��>��|"�g�ħ!��>���1L�u��(���2�L����S2���K�Kf2�N��<�N�y�e>xL Y�W{W��&�}��^��`$�
k�im<^{`UۿL���?n�Bd	��
�q��x}�sv�ĉ��Z͘LI�xƪ�d�������`�t:-����,M�`���sY�R鶱�8�a��(�ػ������ͅ~�}4�j��`�\���Ⱦ�n�*hd^�����X'����>��<y����p�y�����	T�o�JLjL�=o1�}���l�]veWveWv�O�� �]ٕ]ٕ]�AK���E�5��5��r�G{zȽf��`p��6%}�z����?�~�����;z��Pxquɬ�gϾ��^��{2���ρ��b:�?22��d^�L#��R�<$2�w���F��yI�OL¦�4�Q�4ɛԂG�y������5�B�J� :doo��Q����P�~G�[{2���l<���Xݔz �>�,�����O���2G7���mW��"� �\f��A�䵱*J�k-%˚<|Bf�AP̃tFK�g`D�q�� "\ 
Yy��(��y�6�c?P˛>�U��'~�,���P����;�L��mh���J� 7��(v�%��Ŋ�MP=~����e_°������uΠ*'��/0�&�C�}Q��� �X�j+�5?w@�%3��5
(O �^Ԡ�� �#-�l��(`^�I�� ô����ܷ-�I
g�]_�t�ﾶe�8��]G���O^23�$z?��.�-�c�8�j��-���*GN&w"w|������b��ΏÂt�}_&���5����\ݾef�`��tm2?�,�Y�v}RI��s� ��f2�l<Ȅ��W��[m퓥���i��3���� 2T!�7�m�D-�3�3��bd�C��f���g^�+q�%���f%�>2�7���r$D�|��M��0g�;@�ғ������f�m����,o.�+��G\r�Me:%�6Re��.+2��zz.��?���7�.�<h@����R�t,^������O��ˋs)}�]KV�u>Dp5�/8p��|)���> ���]�T�|I��A´�y� �0�N�5�9
�,���?�νN��<�`6�DUK�.���{*}Q��'n�I ��O�۔`(ru���r*��T���ۓ��4Z���I ����M�^*�a_��x���Ͼ�>�"��|�6F�}�s��d"�d*��]9~p�Y�M%��C�֕G����%�HMu��w��4�狩�&�Z�^"���uxh �X��@]-��R��G����2��±��Ԝ @?���ڧw�Ȝ�)�I��i�n x���!�a� d���� #R�	�)-�^�}%��e����$�L?9�������9J��C�l4��P"�����^�-�N�F�`�;�+�y|��I�(d����:��_gdoY�c Yf���0���5=|��~�-��gru=&k��`Ou���9F��[�v]�$�����'Sq�*���6�:���}&7W��O�ޡ`�5�S-����:';��}��` �6�����¼y�4�l�̱��[��kP�m�n�1�y����)L�@0�ϖ+�t����7�V`�G��e�������P��z�q�$u>]�5}��b��/^�3���}�kt�? @�[�'?���h�=�y���Jt�.6��Z�z���}f�W�Ѻ4�Ll��{xtdf۾�ǋ3�N����ãcz��Of2�ʽ����=��(`�\]]�G���͛�{��{(ayC�(�~I7��ľ��,jH,��%�C��	k��8��8�8���#�4�?C���a�`�G&%���(/E^�po[3/�ؗ��ᴿwh��6�!�����m�$Κ-c�@���?���� 0M��b����ח��k��p$O�>$�3ձ���sI���Nk�O�4���In�h7����������?����p��#ؗ�w�AO��ʺ|
�������x���M����w��veWveWv�O�� �]ٕ]ٕ]�AK���#��ծ !ɋ#=�I���( ���=�o��T�z`���=�|��{�B�3���O,�N�T��L~���"��N.���+�0�^--��cy��<|p���Wx����d�M�����!;Qb�������2�߀4�[-�"�������6��p.���x|�`����_�D���;?}-� ca��Y���e9p��.���CFmH	'����<g~Y���@� m��;��ДO�0;���s�Mm"�D>�Z� Q�B<�̰��-k�%��TY�is�?����@<��%��d�
zEX@ ���4�� ��_3�m#�Ȍ�P�3���k��1�T0A��Ϟ���k!��v�s��7X6h7d|�߱��I+1�hPA�h�ZhRww������%r����@��D�E�V�]������x����å�f|�Jz��(wuE��g�:`rW�J�8���nq�3�����ۿ���Ulf�B�"�u���M���Z�r���4���֙����n?_3?���Wi
���0�4jMfĒ�Tn�1��`#2�	fx��!�DMf/3�F��I�U��?b��Q�(���4[P�=��ٍ�Sl�~)O%�i�)�!aG�q�1��W�O��,��1�#���E.W�+9^�e8:�A��2Y��|��D���v_?�<��W�c�P�L�]r�9CG�j���٘�[� h[~Y��8�[ �>���!)ײֺ����^���Bj+���� �q3T�e�v7)���^��l_��f��mܐ�	��Dfc�WyB����]?�ܚ�5���5�:�f�a%f�()�$�A7�'�\�p���� ����*�9�4i�V�D�Ҽ*�9L_�N��Gm�K�=>f�~�� aԮӒ�0�J�m;�Fk�d�)d��J��#�"�g�^$R���N���@*���@F�Ld@Y�;$`YMq������a���% ��P��M��2��V(����`�m�M�K���n�rIQ��Y��hT�@�jcD4o����������Z`n�:�Hv�>�\Ll���� ��f�S�	^�����`�;�Q��F�ñNSf�����'�uG����{�����������(!0		)����C0�l,1�$܋G�L&��T���b��Ě���o,1��Yb����}:;�ao_SU� i@t��Y]?�j 7��T��~&�:u���:�w�]�HG�� `l���C2 ���g�ޜ�߉���<]�L��^f:]l��V�t~u)ד��~�J^�x.$�,W��m��s;�� �씱HQo0uW�A��+�����!�a�X ,�煜_���_-_~���{�~$�A��WW�r~v��Bʫ�{> w�c����<�:H��A��㶸�A�;��J�ѧ˿%.�{�B�U��xR�-m�]�,5��fB�j�ڶݷ4<�;$�qxx�������� �:<����i��H ������g}�����ټ|�����ұ�G�_6��٧����s@/�Ii��k��/}�3�޲��Xh6{r�c�g?����翔��yW�{#z�!���kuD��,!�I���mCic.��V.���c���+��+��+2e��ʮ�ʮ��^�{vE�̨ġ�������o'8h���0��A�g4Y]�i(z��=%�V�����j��w�ӗ��kѣ��z��\���n6dv<dٗ�#��O����!���A�zZ?L0�F���EF"��N�I$K� 1�@-z=oH�I���r���<z*�wޓ�W+=h_]�>���~����8@R3=���'rrr"��BNO+29Jߤvp��d�P�*ߘ�������%h�^��}ֽ�<IW�eB:�dD�p�F�W�Q�<�%�Z��7�$<3ބ4�;����C<�u2��5�}�8 �!5M���i% �f���V�X�Rh�m����8�LW�6I�~���վ�sL�shao(��%�zԝ��fa���){���8D���AJ�J��\r>&�>���EYf߉A�bOE`&�"w��u�_P��It�8��".$pV��Ϲ�d��^�o��?�#j 㻯�J�����}O�|��5��۪5ڿ޸���UuoA"��N����B��s��$�-i��L^�a1���c�cYt���sĞw�6�H��SLc^��I3�0��AJ b���=0�Z2�G�NW2_-xa����@BF���@A��e����KGa�~E@QtJ�۟^h&��M��נ�q�9��-���ӱ���h.�J� ���"���K)o.��:�)�u��lұ�&�Z����{*�I�Z/�t��g��#��.h�+#K[x�tMn�J��DdS�?���Z��H��g's�s����g=G"ȇa���bK2K$�/*=}_Dɬ���~t���-0��Z����T@�k4�2��d1�W�RL���q��z�Ǻnc�T��=%k����y`��Y�`��qS��t-Kt�N�� ���?!�Dd<+�B�̠�؜RQ�F�_'�Ó�T��@ǂ���~��D`)������^K�Ӥz:����gu.���i�  eR�2�I|��0vf�d�5��;
�-3ۧ�Qm~�so-�C�+�C� aEI$󬨜,��V���Џk!��h6F���t)���7��#�X��o���$֋̌�ky�~�����^�܎J;����^y5:of�Ȝ�b �Ι (9�ٸy$ѵ~(��G�</s��G�1��@t�:Bҫ�nRr	k��?��������5d�oQ�	s�y�xƒ \���P���V���e�LI71����]f=��̱.��v�����[&^���?E� (|O��
�RD����v`�G=3���^	m��a^XЇt�>��H��TQ�R�凮.���Ҽ�]�b�f����Pڽ�Bg�2ӽ$��.�t�v�~�p�gτ�f�L8�f�h���t�s
d>�����>�[��6����'�y3���奼xyʺ�	��7�+^�u�7�G����C�W=m����þ�4u[{MB
�>��X���'oU����i_ǳ(ܘ,J���cu��c� ����І{(JQ�/�XP���ir/�x�{�c��G�/��ឰ��b$t��-�	v�B2��g8���D�?~K�e����o��������3��|kt�|�m����F�{l���2��:N��=]/+��t�pp |�����B>������S:�| ȀX���u��,߱7�В��8 K�vGveWveWv�O�� �]ٕ]ٕ]�AS�l#jP���Һ0 =:���$�J�"��k�	+���z�߰��
?��#��>�0G�����&�8�C��Ϟ��@��u)��L�UB}v�r!��bм��ހY��Qqi�[�3EƁ���zxKˀ]�W<���Ph6��`f���T>��C�����?��%�`::����S���g�LTH��yӠ��,N1 B�e�,j�)�a@A����?!�9�T�P����y�8��Z�]��Ox`�����OP����~WQ���R��e��VR#h�i8����y�/M3~�2��A�a�|<<2y�w ����$/��%e0u���ho�����u�l����1� 5���;2=4��Oa}*�����Z�
�^� �e�
M��*�,*K�������_P�<��XQ�;��.��U�&#T�S{||�,aɿ�4pWr��.��,�_�p�׃�{���==+�'v�ߗƪ��cY0�\��l "i�o�S��In-þS���b&����H,C��Ԥ��������d+��{��jb������n�.��TD�Z�>�����g`���Q�	}m�`(�i(�bm�|�bC����Nv��F{���xȸ��Y �k�cNY��S$.^#�x&K��}��f$�AC^W�p&�4��K(+���qy*�͘�~9+d0�ȓ��uɾ�&c�-	*�U�Et<� @B�F���O~d	�'R����M�̂nA����ԕ�� �^�%��{�" ���{M �t�_��Z0�1���=�֦$ �g3�$	�L���S]���T�UL߾�ٓ�\n���8�u�D�Nb9<���F��T����)�������!��7��Jc�-��A���Z..A�o
2H���A>���c�<�p>f���î�녜��|�%��ځ>�XF���r#77�8�kOD�' `;���Ø�X���&G՜��Tt4�(3n6�������l����b��k�`a��s�4�b�w���k0$ ����|/��T���Ua(���c��<�7��Ǹ��O�?�N� �q�0 �o�S�@�:	Y�ҙ�ۚUn%���/�,��%⑮�A�g;AZA�,[�B�k�:�>LE���L'S6��`({}�AV��Ʉ�:�d�A�����ݗM��u����-��{��d:�=�b+X8d�.��f����Vs��D�\�T\��N%��A� �a&��L�s�},��/���}��70$�:��%B�@�����X�w�����lk0^t�����@綱�gs7�j�_鼒Qf�s�[q�1����>�:P ����sJXa�����^��2����Cb�>Y.�R\^��8���X1)�0�b����'����ѳ%ÃCۋT5�ڂ��#�{R2��s���<�w!�h� �Kl��29N�-۷�r�>�@�޷�k�������=��}0�	~p��h�~ #�O���I�d�uӴ�m�\Yb��V�Ͷ��C9�wO��=��>���|Ͽ�R���+�_�o^韸n�Di��������
l���w�b�99:���P����>�=�7?�	���>1�v2t T!�e�\�L�u�d�+�rx���������7��+��+��+e��ʮ�ʮ��Z���rG�Y��:�@�f���uN�>��ya�jH�\<�,�F�ɍi4) �p���7���+f;����C8H!�0҃z��BN���f�p��O����0�n1�����	kֹٲ���bi� 
U�. "���l��Y.Y�@�������Ǐ� <�}��������_��ʁ��<y"'Ǉ��ȳ�%fZoHSA�:r�T"�9t؃��/Mxසu��X0��ʐ�A�B�&�?dѭ�Z�G)���Q!�'8=���H~�>��q�^�i��5�Vӫ�0 ��V����G���8'� ����֋��\R�!��EԦ�8�f��'y�Sf�W ��>ԛ@�>x���7k��d�G��3�C0y2�Bg�~�T|C=�C��[�w���B�����mL���	��(^����o,�0����]fP���������3;gk�w�mW����.�^�I�8�����wd�-C���&�7�FQɠd�̿�r�/T�)�:��L�%?����v:�ʪ��-(�fD ̜�c������JƤJV���3`%4sY�g2F*2{��K~?�&��dЗO���u�E��|�^E���erz�#�V�T�X���h��Z�r���nk��2�RP�JNM>��+2�9of��+��y�����ud���3�w&�2�9 �u� �"��@�#��c+�d2�im,���i?h�Owamx�0R�Q2ʫ2�_����q�����N��t�Rh����0�)�&�VmmO$��-}����R����Γ��f��h��J�=}.�=�}�S�ʎV#�pm�0Z�J�{����-�ǁ<x<�����}.����0@D]֫�$���'���6ފ�y�h�h0�K�j� �fdLwz:�62z��㖒/��`.�*�
�P���Vd0m��n��Ȋ޳�n���˞��E�Y)}�Bߌ�ml�h }s�Nx[��Ӕ{Ϋb�!�A�
~6�0zn�2�
k���80	���
@$�h��d]���&���I ��y���֛���7��f���lJ�%�%pPR�z��t�I����`���)�˄s�Q�״�zǊ�� ���uc��O
�0���ﺼ��Y6ؒ�N�����Av>ت�;�����$�V�5%� \_\P��I�Ҙ#LRX�mt���~LY,�J����%�̝h��?F�L��Q�1����Aߤ-���z��Ԍ7!�� ���L,��p{0�i�۾�rq������3�{����]���C5���P��}�$��;�`��鷬���X��t@t�]WJ��<. u�&]�`ƈ<|��-��GK�ߣt՗_|ξ����/�:��^%�f�Ŝ�|�n<?��@\�0�k{$��K�'v�4u��4k{r��}>����ޱr�|� 7�P� �4�� �?�U�l��zn���ZB�`��D�8/�z��|#�B�L��y򶱇��PK?�t-��k ����c��Nf6p���9Þ�iҎ�K�[���X���_~�O|�/�@�
�{�S^�~�?�pP�=�.%7&a�ki�� v
�`Dl�OV:���B7<��t���܁y�麍16�����E����8iy��G�+��+��+e��ʮ�ʮ��^��`aن��VϞ����8H᠆ F43ԃw&a8&�J��N�n^�x�������}������n�{���|������c�Z�� �����9<�g  L������(,s-1FJ{m�|wm
�י�`.�~�j����@��D�2��1C"3�����O^˫/�p}I]��+��/yM %�@���������`h���^���Q:�����f�̘kj�p�ơ�L[~!ȼ��TB3ed&v����=`C0[l�V�����d�b̌u�`<�IS3*MZ��TlX�1� .Jl�@ԧ	��8}N�q�l�%�gf���o���1S�5���R �������t�aD���	��J�@8���� ���Vί��K�m0��r�#���c�� ���7�ӹ�����*M�	���F�ץ��Z��jA�0��y R����<�+���
<W�m�zm�˲'��[�����;�Bƅ�/�̠����|6t������l�8����Y��H�NB�)�@��kzk�F#4�uܣ�O��%�}Hr� ��в�a45<>Gn8>+[�����;�9H����'���8�xn�`��6��H�d�xLW�g:���sԹ#�v+n�,t��.�7��uފ��"���C�s$�:�d9�by#�Ή�_2�Gi���7�"�D�p����F�K���|b]�������f2�����C�'��h?��o#I��%�V����M��趛93`�q��A�|��� �* �<Serl^�T��z�X�ff��R�:����Ф}p�c��a��l[{>��~_�NS�$��"a���{�"�p������H�ξ%Ά҆DK�R�ʌ� ����)��0'�/:MH+!����=�9؃�<�K�1���?a&�Z�ؚ���m�����?�F����� � 4����saAY�����6ј�@��t�\*�|��6Eဧ�X����0_�?k�]�̏��cJ�k�ʡ�G6+p� ��`����ȸh�M����Ս����_/-m�s�v��a�6%|Ot-�w��{��v�O����S��u jQ���R�]o'��0zq�8m���]�:P|6�0��J���H�:�gӱ��1�))���k��F�ms|t_��9}�R�Ӓ��T��{�=�������N�F���X�={.�����^꼌5��d`7[�E_��W�Nk�\8b	&6�y�yF�yʽ����� ��[N���~ v�Η:���f柑��!�^��>��s���*��l2�$4�b 	H0n#��~�{M�-3����k&09�(w� c����މ��2 �Nߜ���9%��][:/Ï��꒿��H��~��K�w���%��p2��7kn���=A<�u��dk�NjH���!���ʭon/�C���- ��t(�v`�e�"�g�/��K�g൰7�	ܠo�)t�c����d\ �ǀ����wc����~��A#2|��
��	�#*	NnS�5���!=Fȃ'���h�%���*�g�ϭ�w=}�6Q<��d�7�1GK�r՝�C�	������7_�7_I�T��
z��+K4"�K����6V�L�3�w��:�����O~�{ѹ.a=ٕ]ٕ]ٕ?��@veWveWv�/QԔ���/���}28p0+��ޡ��y�D��pH�B������3����/��\./���h�e��l��/?�R.�ϑO)�����M;`9�#|��\�����6>?��e�a�D���7�2\.�fӅi<��參_27	; 5���eQ�3 �@�Œ��x�t2f�F�}��Ï����d��D����ܿ�P�>~(k�y%k��g¬҂���d�˰n����"Y�bK\��"@̓oa�����B�#����Z��!��9��A�+���N0���P��� |aA��0��6�a�s��Z}�8��Ƞ������43��HLsA�y��^4��:**�'��6�k��sJ'�� �@��f�0{��,x�����Am��4�|Ԇc���y��;�� ���1��EQ9y{���}Ʀʊ���5�S�)w������߻�����Uߢ�[�'2yy�;���#U���I��Kk����v�1��d$�l(��>�&�����	'?�[�d�<(Cf��"����~H `J�,j�y�{r�Ufb��[	�bQ��6~v�V8y��؜�R��O| ���[�%�~js��T�//e��z����(a�^�eY�4�˳��o�G�Dl�tF4�پ�޳���Յ~�#�^[��D���1�{ș�enA8�]�~KZ%��7z?5�Uw$�h'���Y�_e:7��:���<� +�|��EG�Z��]h�Ϥ�x�h�l���s����H����
��8�� Gg�C�DS�	�]lV} 2��L� �"h���<��2���/y ˚"-�~v P�2l݆(��8��D�;��]OL�ƀ�'m}Ӧh�X�y���)V�W3�(��!�u%Ե���e׷��AWl��Nk��DI�r�'�>a���=�Ȱ��X%�b���\���w`&�h7NO����L���Y톱����%/��8�-1������_:G��9�ja�`�uVzI�B��h���%�0b��<ؗ����`����S�ҵ~W_}��Jt���j-󥶱F'?UT�x�q�#]�Y��I`��$��n&�y����1��{�mV?�Yy�xd��]�ٛ7d�����dL,t���J!��#���W����䝷ޗ��#�7���ɷ��z/ǇL��N���@X�ශǄ�H8�`_.gd����$sq0)��-���[��
��#�6\��کJ�r�?ү�!8 Q����6�R[c��c��&u �a \�B�10kjit��rR]��9��w}�j�����ς^ �J�W'�	ڜ�7ʖ����R�PZ��"y@:�B(Ū�DR�t1��|�y�ϲ�>Ev!%�&윝�����Y�l�P�J��u�Y�����E �//�Z��(#S�t���:��[�k�[C��kc���(�H�3$��>���Ƀ���o���!�j�&��|�j��+s�������]h?\Q^
�w�M�����$�J�
�EH�.
�/e2�q����n��y��[��簟��{|�o���d|}#��k�G���Yl�]�=Ɠk�������O��!mn�XQ��%l����K���>�����϶�b��^ʣww,�]ٕ]ٕ?��@veWveWv�-8�ޕ7�>�.�}�A����-E�u��`֌LVS��XN�~淿�����O�I�m!����Jf����%��9u�g4�l�&��"���RI8���C��?n��4�a~�� �>�R)'��fm�� ۀ<����ǬB
q	% ��V�6��z�\���L�����G����W����yݑ�߳�+ADmPK	��͍\\��%�Ɇ�����d��Mq ��q9��z� ����4�a�:�#cY�$����g� �  ~ �C��H��6*�@ }������:d D!(�  ��lŁ:F?h�(��6F�0w��`������?�6�����pGeh�CnŮQZ6mfF�0����߷��r&52� '�#�5΅��\G�($�|�IC2 x���;X5��G�l���ɝ���L���ek�`: ��P~{�~Ჹ�uZ�L~�jŬ����ӹ�ݒ��}3]w�N�Z��1]���o�� �#���e�5m�[�0d��!2�C�v���ݕ�r�A�k���5��cc3���6)Cn�;X1xOL�&��`c�� ����O��|ٯ��cB�/��h��~��D��2|�5[:��� ��7�2��.�<�Q���|"�o�H7N���>�Џ����wzY�D&��٘�c�L�\ObP�1x�ʧ2�\�|q-�?�vFm��ó�|��&�����xd��1L1�u����%�M�鵻���?�R�z�:V+dC.&�i�mV�=�(�Ո�̖�N�c�U^f,<[^N�ɵ��2^45.$E@<�P5��@�@}�P`���<9��� ^�f�k�B˒c4#A�s2|�!���b*xm ���� ������K �aK��mX5��=���m+'��M%_]�������7*Ym�!����T�p��~m|T��0J�,��#���z��}0�6��9p�cL�`�(d1����G��?�q�sj"��	�/��n[��g�"���M��<= ��o�y���;0Tڜ���=m!�~M��n���D�Gdy�׹G��vW��Rˌ�ًŊV_|����7�L	t��T�NAp�����KK��zSr�ƚfU� ���W�1�L�g�^�t������Ɍ������i�1�p������
��c��Tiu�\��oַ���� &d`L.���uz2�ʥ�ux n����
}-�w=�6�D\��R��M0#�RAݾ4;-�t��p͂<ص~O��?�Ժ��C㥀�g`���L ̩8�T�_������n�$���`Do�2Vb���x���{��X8Y�5|�3�7/l��-Աf[Ɗ�-A(���ם��ӿ�� �*��L`On���s&�|��O�ٳo�Пe9L$ y��u� �t�����iuz:
�!��1��������`\�א���VZ����2�3ct��)p�4���Ar�s	��;I[����$B6e���W����1�Բ���:�ǒ螳�qp��}���wH��0,E�))�	 @�T �*�d2T�iSם�I���z�h`�@:�~A��3�����:�<y�-z��Z��n��j>�}�X��%��:����e�p�^3�i�zd��˯Q�m<щ�ۯ��/u����$�`�O
�gl����X�i��uS���B��|�!��������(e:# �+��+��+�e��ʮ�ʮ��Z,�h;P#�pu~%��+)�����z�}9<> ���z��F�";� �8;=���^J�2=��ђY��Kh�/x�-�L�QWQ��\r�,-%C�^��D�ӈt_,��3����R�ML3�^dCB���H���a��M����<�:�F3p��?N��>��H�L�=f�Ј`�����W��<z�T���_�q:��:@���f��zʃ ��6��$(W���0 �Z,l�ԁ�	2�� n�p��6��χ��lG�S���dL
]vo�����,�)u���a�z� ��w���Y��!8���za��c��WY�d	?=��<xH�HV�m��X6r��oS����F"�v�h�� 2t���1{A��r"���4����#�68Q�$0�t˘m5]�XxAPY�d�o
��S� Kݷ�x|A#�v�Jf��e`>���(%��-��Y:"C���)�TZQ�)����t1��Z���AF����_�I\�c�<������sg6���뀠^Y8�������/|�/C�q�t��y�� )����̹,!I�ںݠC�i�C:K��6IMfnA[ In�C,�rc-F�}^�ق�G_�4l��T�� p�>S��#�lh*`���sNV�ȤMi��`KAp���O-u�a\1�5K�����?�A��|���siF'���@� J��qK�X��˩,Ǣ�\�	*�0���W����Y�AT�N���W/Ɏ�?
����X6KI���:�u�}D��O����3���%��"����M&���Sygݔ'� ��'�2��6V��-��Cf����l1`�D�E)���9��t�k��� �����!�Q�98�nm7G�5��I�+�d�$���ʂ��ӛ�<��	�B�?��JL�s�)�FS��	b�fE�	h������6Ow��I��xc {�@��)��1١f���d��-�	��*����aF;W8:4t�*�	�`j�k�gr�s��"K]�d���](�������C���L�q�������a����8Nk����-ji_�f��\�X�6���񠟄�A���mRi�`��\�u=H�K��Ɖ8����j��;F��J 1��d� ��<=�,�ٳ3��-]GO���M�17������ǵ{I�ӥ���ۭ���e,���a2�:�̖[�
���d| �P����� 9������{dJ���b�Z3����9��}�O�C�uDp�jz�1	:�+!jIf<L�4�.�#������I����S�x�h���D~�ӟJ���Yd7$��z��|���($�2��e�p��c?"x���B���,�����Z��)���7g�i��#���|��@�������{�L�9�.���w-V��8�w�	��N~n�gZ���WZ�%�D��`�N�
Ϻ��h�i<���Q�<�堈��c� ٲC{_�^���%��/>�d5g�����;ʢ���yo�H��+��ks�ʖhǅ�n���̈́L�@�C�H��B�����F�ؕ�~�J��@�F�m����G銬%șQ� +�L���O�y�i��O�|0Q�X�y΄�H�IK�8� ѽ�fmLX����;o˓Ǐ	Z�=�ϿD��O�\�0Y�F�ƳԽY�Z�D��VJZ�"�<�{� �vh�3 �k��˰na���1�$����m�;�'��?���L���5�3b��k�z�ȵ�ǐ4fn��m����%��pVH�| �S$�,�+���28p�.��e��3s�(&Qxdp�.�ᵞ>x$��+��+���]v Ȯ�ʮ�ʮ��+�
����P��/�r��#98>��`$q��l8ZL�AAtH�z�JrهƱ��ߔv�i��Ƞ��)� �:^�0��у<D���?��с���q�U�C�����t���#s&����D�ɶY����3/����@�����3H `��S��������Ф���'���#����|�����+9����_�����l|n0�S���N��t�"Q#���I!u�Kf��NVmH5��&C*M��A�%38�� �P�o��iT:)*��P\0�@��<�=U葑3@&<:ОAh � Np�6��a�|p��<7"g�ꤓ�s�;Sk=l�4�,��ӆzӾ���s�0�#���s�k��d������a��!B��ָ;t@ ?�:n;���]M����6�?�
���*����H
/��i!܌Ǎ��{����������B���CϘ@��)���_�k���g;z�L���˒�[j6Yn�Y9�3�5�sdd��*�N��l������+�`PU�ꨃa�٤�.br]̯v,�ڟ��ݛPxb���k�z��v|��6�NuL.	�u�-�Gt��Ht��t,��R�/0Iϙ��� F�l����o��F.ޜ�KH����^]˓c�N�錘k�2-��J�m1LG� � �G?@|�����X�y!٢#���*�Ѷ���H��s��,%3 �f�OE�WB`��2�!õ��|���̺}��S���t�o��x�虀g�@��)6�h�e�;�` "������v,�
0�3y��2v�d&ryV轌�DZ�߫��rO�L��rt|@6_�s2�� ������f_﷖f����iY�b*��Ki�����	��Z��0`��li���a�\����-���g��^�B�$b�4O�VK���y&�ٕ���`VC��z��o`ncvz�1��^����@��dn��+X�D&�����}�WK^9��s�C��k��"�B]&I�򕭅��ٓ;�;�n`��9�3����ϕ�k�u=�|�k�t����й���J+�rL�d^Fn��A�rua.��0����c�Z¨�2�e�*Η�|;=��X�#Ȣ�� X&:75N*�7����}�t������,@�^ �!E�~�y�,�s!n�\�4)����S��gH���<��.6�?x��	�.�}�=y����m�A���o��}�=����V^?��� �����9��o�������/��ߓ-�L0і:X>��O���\r�[�N[�?x ��{�O���'O孷ߖ��JG�\�t�> �&ج�)H���T�C���|�3� �0��'�#7�8&,]B
g�o���w=�u0Luz����w���}�)����?d)K2^
)0�Ot�Ól1_��G�Zϒ{$ k��t�t�����Ώ
���H��}m{2 u ឱgD���қ{$��z��~�߮�5�f:�����
��c	d̡�5CS����C}~`��u�d�J�]Y[
������:%p�u�6���XsX�u\�9i�!�V׃�tu<������d����o�f~g�}d�H�<}[޼~I�LP�h#Ȃ�?c>�ф!L����K�Y�3	�<y�DN_�0)X̉:6}���V 3|�J\�N���z`eAI�ң������F�������ײ+��+��+�e��ʮ�ʮ�ʿ�Ҏ<�Y�6N&W�M����\�����O���'2:<�!��̠�o���?H����0����7�9IA���3�
��$5� �>��@NNH�?���܂��=������H�z����ۭ�t:-=l��j��w�g�Ȧk��	�Z�<�1��yMh+��}�M*j���f�=��09�-���}��/~)�~W�����?���A�Ϟ?��I���a������hŬ�&p��3[�eXZ��nP�&2�N�����O����+eb��P8���Z�N��,Nc�0L��&IJ9|tj2pӬ݂e`դ��!�+ʧ�e=�8BPG�S8�Pq�eAgԙ�^Ij���7"f��>0IG�.3��ȉ��سiԔ�b�f@	@<�-�-�uJ�i�i2����~J�c�!�A �2���#��4A���E��5��9^����D����8Nf���N�t�o�?�N �<.Q��4�k�Z�l՜Y� ��w�#@<GJ��֎�.6�����{�D���5�Tg_��%%�*I'5����\>[~�"�f��M����:����!���2�o+�c���o�!P�3coCz��E�>��'-����^�av0�3� � �Y�����$�gx�`� ��7�����\��$%+��ʜDLƬjf���k-���E��r�!Qd�`^�Hx'h��+c�-f3�O���`����s��;x��H�rɀ�沈���q�0��&ҙ�s��Z����f2<J����慶����){�})����%K;Cgt�	����{�}Ѝ ~d�n���J�]�a�1}>�K��^&���Q��������NWr�J�'�US	�DF�R�eH��vg`^����ו��:_�}&�L�^|��GXS`\O$&2�#��rq&Ur�_�́�NT�#�e�
'��漐�&Q��M�x��Yh�m�&�t��ږ��Q�əuc7
���P8c�0�s�*M�*��ǧ�'�D��-'��{u�\Qf2�31i�2k�b�&� 2v����؊� ��R� 3�:0/R�Gג� k,S���KK�W�7�n�rR�K���@C���d�(�Yƹ�>�ġ�dم��C��e�f��~���N���}������{4R�U>��^���譎��П蜤c��/�mᏀ��ᆾ7�7�� �Q0Mr�xqR&��1i�x�I��e9:8���!��{��q�s=<ڿ|>g$P��ݷߒ���WB��Ԏ���cy�����T~�����ӧh���/������M��_����������}����>��G���6m<���лL׾�3��lN���d��ya�C��ltj0��:6����L����9M5��q`��@���9@ 	��Ͼ����_�\}4�����c�����{���f��=���!��!�G:����KzM���܃Ĳ��1�������8�ײR�O��o�[��ɮ�.�+*۫`��b���`1d�r��V����F�e 3|�o��>	.��:<ܧ��	. "ŭ��ɔ�9��9ec!u
���9�#}�.&����5i�z�qo�r��V"���{��h����6t?yS�i/�=�/^���_�z�����ɸ���i[co��83�慃���'/>�uuv�6�at�Y�y��=�������H�e?���[iţ�#ٕ]ٕ]ٕ?�@veWveWv��T��,�rr�O_��-2L���5��m=�&zB�d��^��Ս%���:����"y<@J�t�Ut}y���v��~#�O��=��h('�an��~��)�Ì����b��!�����@�&8BJ��܋mP�G�Պ�`Jp�C�@ X� H��i5W2���p:��h ���%���G��H����o���k9�C:Lˡ����@v
�F���Aϙ�C'%�-�LD��)�`:����F8ø�~?��n�]� �0(^�}����5����j�������w 2x)3E�*�%f`0�)&�6�&�A3�܂�x�(��@G�"����~k��D|V��A!����dIh0Z�[&����T��3A�g��q�Z�f��@��]��6(�BP�A�h�;H���V/H���V�	u�z��V�-��7������-H�����=��5��o��;����.����d>j��(��j�]&�f���*V� ޡXd˄�V#��A�?$�Lk�R|���Nn<S��#���B�Ł&�C����;�Σ���qB��Ew�m�E�Y�+��ך���xXߑ�|�b����K��g��C�Ab��؅,	�ڨI�
�Їځd�k(zT��`�_���4F&��cY��Gg�L7S��k����v��%����軰��/̤��cIu^�M
�L.Jd9˷_|*ݳ.�hd�"��Ѯ�w����o�R����.��IZ���mn���%�������oeD̡|^��� PTk%+*��`��'m��2��乬�S�f&����-g��ܼe�ta*�`���3�9+d1]țg_�V���Pg���OOe>~%Q��1�����0�N��B�!�@�f)�r&~cA�d6�g�!)[D�x�6�E�-7��R��I_�9���[%�0�6�j_I�u��B�ri�K���X4����O_K|x���>Ů]Y�%�9��I恖���n����Ҋci�
(%���l��p�Wؿ9�C
H��6�/�$�ߗ�'��c���"c� Ն�6o���Y1U�� lb���[�Ls��2[���"Џ0X��� �Eo,�%�}�u`���~ x���k�G :���^����7������|68Ox��g���<(A6����Q>��O�wޱ�.��k����y�?��#��D��g ����F���|��O�?���F���2�ߗҷ9�ᣇNc�1�����U�m	��O�Ho8`���c�'�%@��2�<2��ZF&�r��#�e�9Hn��L��瓵�hJ����	{H�f%Yo�tDr�YFqN�X%Q�������ƭU�8r�,u߆�6ht��da����������s)=����!� �����o�R�\kۀY���נ���`AJl�C{!��:|.�Vl�D�މ�A��IÕ�D�} �C�	K��AۢE��DͦK�p�qφ��ېU�1�rgX�釢?�=�rſ���Ϣ0���ol��1������c6�l��4e��w�_��=3? WP�s���G2��P��Q���=�0�ZM>�N�Mi�q>%['w�B$1���O��gd�F���W_�L�^�����zF ��'�u��^`�S�.��_���ʮ�ʮ�ʟF� ��+��+���	C���!�3�2O�݌�
���țW/e��I�.Ry��	i8�!��:h��1���|x9�!4���mD̐C s|3e �o���^/�a����
��� ��;}tqФ�� q0D ���1�0$�'%��@���oԭ,��qyy�C3�6����}��c��A�܂$�fW�ݑ�zC9�ߗ�GG��7�|�������T�88|`�zX}uz&�|-�eJm���y�<:����^�?��r��A9�9xv!�g�ЀRIU��~��ڲ!�d@b	AOd]�ij��t���]?����峠=@	��Z<;�-4[m	��tMo��~�����#8�� �f88اO���� p�ղ����[��`1"h����d-(��݀ �F!ӱ����י�(`E�l�\����pA��֬q�GP��-���HU|���7��2n�4���?�]�ϳ`(��A�)lXp+}���J-�af���A2��s�~"�&��;�{2����3:dp,;Ьp@�LԌLx��p��91�'H�軽g������X!yf�z�F`����b��� �ud��G(����{폀$�i��t��&)�~��M2g�ʤ���[ï��(��qm�	��pm<Fo 8�ó 5�='���F�]�0�J�e�c,��72Y�,8>����F�P���t�\#�L�b)�,���f	�8}�9�X��.�"��&a�Q�49<�����@$���s"�y���-a0��Ӯ" 	p'o��I,�GR��e�[D�?����0@ʏR�ʂ�Ь�T��f�u�$� \�9��� �, �k/h?����*c��޵\�'{�o~'W����t���5�K��ߥ7��S:�!)}�\�`�']T�@o�3*��>{�ǫ/2�f/m�ϵ��/��1v���UF��e�}��iv���g6:�G:_u*]�Z�I¶C{�	A�� iy�lz�:� ��Y�D���K��ˀ�lx�POe�,L���?�%{ 5I@�6����|{��U��lr�JBu�����.5���
f�7��5��O���XzUU���I3��ό�=�3֒�_Y,�rT� �ɭ1��;�Y�h[,Ɣ_,K
���̀���~���u�\�(=T���OU�yU���3�1 D^ɽ��!�����L�?zLf��Ɯ��4*���{������#��GJK�KO� ���<x�XN�?�N�'��X�R�'��wx������9�������u�$J�����`��ip�C�>�lo�y6Wk�\�W-�9<Y��yل�y�}P�)�v��o�(B�{a�x��=���� ���QO拙��_���<s���@��g�a�
�}0?�t�h6�y����t������Wӱ:ob�o��^p�J�æ��ͅ��X����?f?��)�^�؟$��}ʙ�:l[���{�&I��J����*Ku�=�.�4�k��ƿ�4.Ib!K� ���uwUee�
�.yϹ�#���>c�xmٙ��������s�����N)I�O�1='E39[kU�ya�A�qJ��ҏN�QǞ�x ��壏>bMR�@FE�cM���f��lS��H*�n���	fZ��W�Z 2�������s���3�Ѫ�x�L��}}����翔�vM)ӬZr>;�d	t=���+$.��z���F� ��L����X~�Gh�|��9�� ��k�A���{�ˋWd��&���~�l۝��Bb9�C9�C9�v9  �r(�r(��S��#�lc���L�G���2��������n�?�7r<9��J�.�2����.�D�ZB��L����\�B�3�g�R��`P�l
j#[r|tL�ql�,=dv)�CP��nް�D�����CX�!h��#��6fԇ������R���̼�����Ƶ4��2*�)�΍�>=4��n�����\���Ʀ��Ņ��|ͽ���57}8�� �|G�w��ʉ��UsC�L��o�!`rJ����psPa8�َ�HS;��8Gm�7�� 8��+��d��B	#ˊ���,��3�hA���}��iS7���G�5B�q�Z�p�2�Hd0��;M�}g�n������zXX ��'0���������Ay����3x���iK�x�ܖ�6g̡{������[�;�G@9
fs����\�e�,AP~|�%M��r����	��4��g��� �!p�������yUW{�*�5U-�JP�1�­̗�~�8	�ҁ}(i���p/��p� +@�"�tm��Y����kg0�;��]c{+���x�j��$��f�s0���z�9�ǋ_��]�F�h���@��͂��V�2=�U��m��|����1b����}Q%�)�y9��ڌq�,x�₱��8󺉌{����y�k3=;���F�}�2XM���x�Hr�W���&v������dF�R������J�~ �a ����!��qRQze.au+�&�0��!ⴗ��?���������_#���L��i"i��ؚ\�g�W�>2������ϛ������;��~��h.�]�h��+�62��S���KKsY�2}Oߑ9�|� ���>���
dy�2��i�sO2H�����W�2:-e�ױ�Y��&��	��0ܡNG�X��T�N����)�&d��輖��k����R����K\��������	"���S��g>1&A��v^ ��X��ðKK�|�Z��t��d�CJ��oP�(F��m���"��c��� 2�z�q���`��A1x24�2^��j�N������^Քmā���DǩZV��1���e�:�@,�qY���D`��P� 2}����WE��{� ����-Xl�S`m	�l2HB�8fC�}���EN�>��EN��8֒:��0;h� 8+nΘɯ��Ly=~����Ys�<�H����+b��v�I����k�B���]���=�u��O���m�/x�&YXJ��
���iX���ѵ$r�k�鳗:ޠ��b�FB�j}� +��x��\�\���J�~�� �9� ���U3%#�T\�ɓ����󟝞��}�c��݌L��6�0~i2����׀��ט�i]�j�:ެ9����@cn&3�fܬ�\��8/P~��D̙`9�-�q��]Sp]��q��l{f*A��m�;�y9�N�����7��:�`���dRY;��6z- �S-��<��˶-��X�:�M3O3�׺f�9�� 	6K��d߶[����H>��G��?��
���i昪��#�Vk�Y��W���o��RNOO�N�Z7+}{O��������u���^����}7���C`cd�8������𿹙ƗH��ʡʡ�� �C9�C9�C���(�[AˠSV ��fPf�,lc�ok�^@��k����A{��7����e�W (3t�=�M���(e���N$�a�ޮ���Y~j �>=��4d�`N�ID�z���^I]o|Y�[�A�.�T�|�M�r>cp ٓ��~�������AJ?$]��nu��J���[�ņ�2��-�n�T�NA鬨��rF�J��Q~����?�c����X�\��HG7��`��,�NƳ	7�ؘ���G��_�'�|"��¤�.:ԧ���3�<��YiR3���}��A�1)��ل(��s�u�[��A�0�l�#�H��D`�a�3kA�6�q>%M����5��8�0�=C�57� Ö�/0�t E�C�w���Iy�N��aV!b��7�t 2���M=i��P�$pU����yk��]�/��+����*�ʂ�3���$�Ƶ��{6e�~�D����T�j��	3���v|x_q�X �*�H�3�;A�C���R3�oM��~�\��{cw�/���L,`��N�:�k{>�o��!}@	9J�����)�``���
�)yP��8 �W����=��6�1[9߿��?��/���v���2��%��&o�X6y]�g+�� PU[��v�����PR�Ό�	D����O`��j�!e�$kF�fܘ Tm��V����� *��@�8�F�`%e�g:^�=I$ձ�̱�	uJ	���;K=]Nq�ŝU<,���vc����F6+=�P���^2C��:0c77��1}����0��sm���������t��t��n�[@�2�1?䭞�����,���X����V�B��x:��S����F�1Mz7҇���� ��0�B��3c=��Q����`W���|+7�L?;�:ձq7?L��ց����(��w�s�J�0����`�Uuz�!�`�T�\V��:�K�|ၽX%G�����KE���k��%�� ��V�N!������ ��|B�*�gx��rc��T�����grZl��x2*�{	�A�w 7[t�Nb�>#!X|1�d���8`FE�8�zJ:F>A]̅~�����9`�} �=x��ס���ܽ����\XR6	c#��r�6֟c<���� �0ǰ���t ���J��?�$HxLC9 gxր5�lu���֫ip����	�?G�kH-(�����~ �3<w=��j��n��HF�=�6��Ľx�V���k2�>}*�n�u��{��fHMFc�r�k��Xoiv�Ly}'`)�?y�{ ss(������&f�ԣ����6iuF���3y	i�ٕ�{�Qt�����ǔ\mVL�v�4�h�q�5G�q_��B����>�{1_9���rQ�N���6C	b0f{6�����IǶ��k��������<y�uw��\?ח��;9�|C��ƍg�]�sc����]�f��m���oJ�o� ���ҙ��9 IE���b��t�u~j�h�wաߚ��|�4*��xf���B��800��N�&rzz�y�w`�R�	-%��[�x�X`�p>�(�ʄ�����?���$(�vh�3/;�w ���h9%�jG�j�X4�����sy��7\�A�k*�Czo��Y3�����k������,�H�ј��c��O��9% M����}��{��8{�������g�����eo�r`�ʡʡ��� 9�C9�C9�?�]c�Q��` ��0�E�~ПRv��;����Q��������PN%/`�y$� e`�(t�%�r�j�\v��b��p��F���2#z0�$��+�/W̊��4\F[�4�M�>A?`� �X `� P��5r��E��A�ȗ����g�� \�Q���1 �Fm�?�>\h�/��1�gs}�Á��G?���g���|��+��&/I���!o�>^�q,��#y��)7��}���"8�%�-X� .0(x��Q�Ƴǀ�̏��<s����р�v�" W����'�����O鳎���B��`�j�dV!
�9j�Gp�,K�y?BcQ��� <�&�Lp@'MMw��r����r����qƹ��2bȀŹ�o�s ��ϖ�֘d�����*%�.��Mcԭ�^�HcY���e�"2)/ ������ȷ��}��p�ˠ��|����ϵ�	��ϼ~��k������h�y�ׇ�PN@��Ϝ�
���y]���{q��6�g�ޕ�W�<���+c�}�#�c���6c����ځe��a�"~P��(\C���;L�5���
RkƧ�= �/�%�q�1��LU�L�!a��o��&����i��P7� ��3�q|�f]!��L�t���Q8�8Y�x�āClK-C���9(�"۾��1#>�w[j��ɺ�JC��X�����k̟��t��P�rìe >��-�X)x0#N*=gO�4�q6��v΀Z�cB�X���	�p2]P�j*'�T���m��PD<{m`�d�g�k�N�8�X���-Ų��$1(%�=֯�T�=�3,6���f2�a�3��`����E�곁�s_}��$���t�R�`�c�0%���8�g[ӷrs��\���Z�R�<��:vt��I�74�G�y/C��J:�J��T��x�l���c��>�ⵈNyzN��Y�-����u��a��w�6
�G��<>7b�h,����ze�:�$_u?�5��� ��@j�.W+���������H믩;���ڦ�4q��$V�Ďe�m� ��r��#S�I:t�( ˓�&v��R�M]�1�L��r�����66�%e��qUT<�yFU�{jAX$'Tھ���+�s%aGb��r�Z����m�o�|��l�o�� ���� s�h0���~�7�s���s�;2%*�Q�05���{���LVk%� ����S�����km�G��Z�Έ>f&���,7�K���9vN ����5I+'�qp}��cM��`3�:�u�K�>�8�y�F���ū��Q�� �
$� �*����3��7_,tM�ӮW���?���ɟ��L�N��������w���cB� ����wh (�`'����A"j<����\>��]}�kˉ���c�C�ޚ�'��q��Km׷����'��٨�^#k�	XO -�_�K� �FI+�x�c�L�:�V�97V/h?Enr�捖;o8cX�1�jѿ��SɌ�c<�z�Lh��rM?: p�/h�`�o�[�k��k��`d�VS�'S���d8�q,��t�9,c0��N�R�8�{��jc*NB�C�0�gp���'����@�V�P2z�,���{(�Zm�o����|��=����&��\C@fOҜ�vF�ǚ���J�p�G�o���h��������������{n�s͡ʡʡ��� 9�C9�C9��{��,�
��|�0sR� �D����ҧF�f��F���;�����z�4��� �WB�G7����RUȒg^)�v0�MU��g�%�]�Ȩ��Y���X��yB��&[Y&+���}^�$e`���A���0`Gp�`ƫ��.B9FZ2��J7�����F�g2�P�ۂ��`�iꊌK�g۵d#G�44d�wt���{_1�0�9p2N;j��nV�u��A��݋�u�jg���h4�T6�z`��u��U�2��v�noM(7�a�6����2I�G�L�� 
���v�`��.�">7˺A�D�����܌�d%����~n��>�Rz0��ýv6- Ѳ4 ��E��͈�I�l�E#�戇��C(��3�%뭾�������}�'~��<�~��̀����5�W<pY�F�p�ǃ�<>U�-c �gH�l���>�r����A���s "���˰D��,�v�@��� M��4��<�@*�[���@	��+c�@�ڀ�����q�rkf	��1�U���P2�&�(��??�-����0Z�4II)2����|J!9�'�v�Le�	,
M���o��jd� ���||"�(�~��C�3�ҋ ���Wm�N�tF�C	U�Ї<ct$I�cw,�Y�`��+��}!p,�aL��xp;_H	o�\zH�h�ʵ��E�Q6�Ӟ�&���	0�i��S�i�c(hr�=0�p.�H�B֕|UH?,�~<��F���ωz�ɄA�!8�c��G1�{ɬ�I=!�|w��d��INes�1����~_�z�)�/�A}�q�//���N���� N)q#��5�G ��1��uC�}���ԾB[J:`H�Zdr��번�cJ�T���$4y�D�)�����~�19�2�U��
��<:��,�|�m&��3����o��_Ir2�<B:;2X�X�<=��xs^������`���7ߔ�ҀT���|>t��!�r%Ni�Ǳc����#������1{
�/۬��[�l���� ����8^h�42�Pq�mr^��GJo)dlGJ�`�Nu�@���i�����(�Cƍ�	z���>:�z8��խ�\���p�o��
�*=������t������c��BzI��T�cx�\�x�,��(V���d�t>dҀ6Ύv��MO����K<&x�� ������Q�5��3���S��O��&#��r�� �
����w�7��������ɓ'O�g?��d ��� ��o�������^~'~���~%���/�#"�����p�{�Ȑ���cONNt��!K��g� ��3S��O�����<���۫K��R�b�k$� p}rt�y{�X���S]ϼ#/^��>rD����3���Wd9���Q�����x�`�cuI.K���/X�WWWr20)Na�? ��9���Kc	��M�T��|����~_�[6K�1��;m�j�T��Ӷ��,�D�L.̧F׉ �1�% �]Ц��!�vk2X�o���"$�!G��T���ѹ���]>�WTsk�����L�'X/�^M@���	s
ֲ�'�����w�1���\�=G���I��dW�' �� ���W_���L�����"kuȄ �ɷ�N�:HB�k��g�e���2�>̕�lIi���,���� v{u#�����k����O���Rp�ϥ=c4�`���֤��{w�{�0@ �����H�����{.��ʡʡ�P� 9�C9�C9��k�#�d�n\�,Y�'G����:_��Ɨ��F=�t#���r��k����l���n� }�0>��d$��J�5��j�����m��$%S Abd�����4Y����̔��0scl�Lr��*ı�T�,C5I��e�z.���i=fK�t3 g� u�2�:Vĝ��pd�#�6c�:���1+�Vw0}m  ��G�8�'zF@r�6�[�!���f ��>�d=�1y�f��58	�ZA_,s��1z� $(��6��n��l؜cS
����燙��R5ͪ��	|���= r�d�]�Nb��G�"��e([�02A#��z�x�v��5�c�(#���V������{�E�nW�W��]�n� Q��ɢ4t�YM���.����Ul�X�6K����c�2؂n�X�R�,!%�G��S`R]<.7PC�y�S�1
@q�� �*��c�/�MQIp�Q����d���A��!#®����[f>�	�V��1�"���W����%=8�����Q�d�P� ���8��{V�q��Z�(y �� ��o�:'��$JxB`�l�_Vf M���	��	̷2R!���Y��zM �Ղ��&�9���!+I�4��wo޴ף!q.���� %�ݳ�dT��e/�KD0!f ��v%7s=փ�D*�$e`�#��`A*Q�X���Ӂ��N�NE�E�0�_-sY�*`2=G`ۀ�Z�_{�b�n�m��hm�g�p��@mL����X�[�EE�[Q��|���i
�d81y���t��$�zX��|�˫ vz�#��O%_�x��Z��TbP-��>Sm4��S	^	jk�=�p#:^W=�r�yk�S��tN�s/�K���2�G�C;+����ވ��!�=g���Ƕ��L���J�N|ك�}.��w��,��RN�L���)�ʄY���;I=��A��e|��C�����X8�����h�����F�,*	�x�厾��s��z)՜�(��s��$�f6�f�u�Y5e�0�a�B��<[�}/
�����	�sA2Uzm���'���ҁl�[>3d�0�"���� �g҉���l,@���Z��V��^���<�����'��e�������oA_���H������
%����\Υ��.[=tD�1X[�2���D�Bϟ>���?��W�ƿ�z��z�#�n���S&���>��\�yM�	u���O�2@������:�	�5�)��z'q��'(��9�J� &�>&V0E_�zc�~��ΰ#��0J���u����x꘦��.ۊ��n��Kb�l�d�1�8�uo�v`� �?�C�4��?Ykj7��2/ (#�o(�9hv_rlB��]p��_�0Zи ������ƴ{�,�e��
�`�v Ǝ��� b�)�����f̱g��e�ޒ8��p$�G��	<�:7 r� ݬ�=8����Y <����_�}u8ԟGS]������r~�D�s�㚾��d.1��������Qo1�b� 彜��3����3��*���]���x��+�������N��x+��T��������tn��뷯��o��~� ؃�[[��k��7���]�3��N�Nl�@9�C9�C��� r(�r(�r(���=�,o��N�ovBi`H�W�I#�����)u�݋�xt*7o�2h��(	)�s���u �l+�{���?6Qf�F�A>O6.�����f�a��b`��-��7�2�D �,Bd�u���*'a�e}���F�,���M3���iZ���q\�q vh��\J 30�Aoȿ���Ʀ�H`|fUã$������^��ЅG���m����%Xgr}}M`A`lF��`2ǋj'���F&/U;/	l���j[�l��T��� +"i}8���� =�����x�_���f��X(4ȥ���F	  ��IDATS��n3�x*�[�-M�*4�+JN��l�`Fޚ�Kl:����eQ�6= ���5����}��Z	T���2
ZI'�
�3v���L���٭�����Z���/Ln%�/D�;�pX}���gH]�ap��#P��j�C.�L	��鰕��͵�X�� 
,� H��{�ԍ�]���8�՟�|@K����3C� L����A����^�]�:������ㄶ�����X߃.�=��%���A��� �� �e�ڊ@X[���E�ƨ��{/_�T$g��_=�$�KU^3?�]J�����N�;H&!��8�y��w�ٸG��� 	�A������s�
�����zW�|Q�ե�|f�H��D�^hmm$B6,�r;/��"���2 %50%�����|�z%K=_w�,����Z���,��3~�"m~k�K<'O�K2Ƀg�j�]rV�����`��WJ�%�t|����C��4�l��\�|��K``��V�իW�ڽ���~JQ����V#8T���p��*��ˋ���Vd�y�%	�Re:IF�c� ��d��ws�8#d�'��
*�<�m :%��eE@��'�<��]&���/��r+��\��zp�1 ց]A����̿���o�W:�Y[���{�����|�ڳ��={����Xq��D�E��4H����=�ف?��hLY&�:,?>�2{s'���+�"���mA������w��PH��$��.�d*��*��f����[�[,y��|g DA@6��U�X�3��9)���l3&Kp���ھ�&(J�eE �}���p()u|t*K$|�ǉB�*��:����z0/Rb����?![S~�4S��^x��������s�v�n��7�o���bݳ�
��z+�ٍ6;$#l��o��w�\�,Ṯ���Ϸ�|0
��2�0lj���u�x^�����}����[}�4�׹�RG��d:�r͒�+��X���T�6a��.$��C^����
r��JU��k��踱�q�YӱF �����暒ZO�>����k�}v���� �0w�I�~3���g��LH`�?�H����2��F�]���_Bc��.��u�G�Hh�Og�n�����g���I�q.0�U$x�ۦ`�j��F�!#?4	�D� T�.t>;BV_���� S6��;?L2�' ?����D�=���������]꺯��j���(p�0AK�R��<�r��?�~��}rT�V�{i���F��ZIѐmJ׏�ƭne�c@�h��εm���'�0Q޼|#��� �
&���L�r��;�)�r�����������'M���P�P~�� �ʡʡ�� `��M/�Mb�H<�����lh����'"P�
�a'�S�U�X16�	$\
	~lv� ��$�H��9RbG7F��UC^Yi����9�h�%|g�I��Z�kJV!0��!6Z /tA�R��`8����Ov�\ͩ�M�}���ݽ�)3�{]��e�2���:$)l���+K�E��$�u� @@)$D7Fáy��|�A(�,�F�@�1����PJ��M̠�Ջhn�kj�c�`q�f���uf�L���!>Y#�|��U���\���?��ŔP	MM<�(����R��# �m2>ͨ�b � ��{"�G���0���Kj�ӏ�e_�5����`����S��-߹;�b�&%�"m�����B6�����Y˚q���@27[���j-�HI����ߡA����#��U�6���m�j?�B02�V��e��+��G������{���c�n��e�j����Ž9��(�d��~<xN�����z՚���g��Akj�=�OH�{~��,M*����Fo�?5��*�/��\f< �µo���em#��0�cY�嶒�"m#����F���ېq4���dA�W8��r��07pό��1�с��c����]�A���C����d~k�S�\fo^Jw��HI/L��A������$M�2	��e�R�K���խ|���&==qW
�7�y|��jϰc�}������ϻ���>P"�v�l�²U��N v�=3��B#�Vי�����B��%C�?�j����W���\����7o�ًG:��:N_��D�(�W��)��t��嫯2}~�yy�w�ؔ2_\�x�c@?�PǤۛR�K�s�G;�j M�^�5Ӷ,~�w�=��s|�@��>��K}��KY?M�h���ճ�����*��Fh>����|_l�k�����8ﵿo�����}�*`�ĝ!� JԴ���X� z'�3�+J��e��7����ŉ<~�X��D��ǒ�lY�!���[�'7�O���^]�Γg�g�Z�@���?c���˾Vj� sg��� ��x�`�	B���z}H&Nu�O|G��e�6�i���R� �p�2=6v�(�����dB��% �����zC��W�u ��\� ��I� ��b���oexf��#y���1Ǵ�!�t�D��kt;���f�Z�b~G����c2`��8�u�%������µ�}�JS}�������?��o_�6�Ȱ?${�f�gan�y=Ic&l��:'����z��כ���ӿ#Q�bY�;�b���|��  �OƠp0��zN�&$�0�E�[�bWݷw�1|��ޮȜ��bd�~�Gۄ��s�m�#���������Fۍ��Xp5�(-�w�6��������:40"⻱�m�)c��D��%%ȥ={����x�L�XRx/̲�!ߦ��%XcI�������T�Gp��&��kB$��mp�0b�:�i������O�ڟ�}�cy�m�����l��'�%{�������$�s��<���/?o���s��W=9{̗^�@�P�P~�� �ʡʡ�ﵬ�w�l�lK��-܈ ���@����%P�'I�����$�͍nH�Q�&ҟ��7��1鏢��0���'#2.u�K�~/����C� MG'c�/�,��l�(���H�[жvo ?�A+u����jA�MP��x�>�7a���A6"�y�����=�&5�{����d��H9!Q5pF�ؐC�)|I!���.ے9фV�������/��'�r~�HҮ>箔�o����*��wA��6���R2&�:�3-E�g�&eaR�ê�L��Ix�7D���#��b�&p`�z��ۂp�U������eֳ>�D����qY.���@Z���X�M��f�����I�D�$����)�!N��>K�$��b �m�RHƀc�m�b�B�f�_�2&��x}& h��RNս,�ؙd����u��=(�ף��qo������q�	*����u ��^���0��k{�=h�%ՆZխ�1\Z�+ �j�V�)h��A���b���{��W{�zH��A8�=�2hd��e�����i}K��|�0�&Ő�-�;�g<����V���w!����UQ��4=�q���G���������?�8��Rk~�43d��u�T�̏��XL�Q��`�V�T�ݘ��ݍ�jf���XY��~�Kg�T>>>�XF [�e��$��]A����u��l^�bfd�l���wkY똘g���8A0�w�����5n'ᣱ ���;k���=ӥe ��޳���!��х�~?�S��;�m.}-��E�!����VǞb%���k}���72��q���Ü,0x
�AJ`�L�+��{O�F��4[l��Fù����>�㠦�L��x�|��[O�ݷz� Q��n*�p��xpc��n���A'�Ų���}�I	〞S|B�DD�v�:D;6�0�Kz]������Xf~.�*��Dv* ��^sL�c |L6��>��u�1� 3�_�IJBr76 �g$
���=��O*��1����#9{4�\�՗vyy��p+�l��	�LFc�;|����;��|})����Vw�_��S6r�u�}k`��S��~v����Sy��3 )X���~7I&$,��q�ڲ>��"�^�	Y%�шk	�;��}���q���o+�W��Heh�ɇ�w�k����B�P8X.@���e��,��v}}˺ � ��w�y�b�vk������V� �:�!��Ѻ"���I�����o����	u����v��L���0a��Z��� |2
��w�ѱ2��ﻂI �Jb�C�L���rl��h0��@�RH�K4�u}׿��B��Tb��>||
>�Ԇw��G#���A�^�W�O r���Xo`���������h��y19U�û1�݌���	k K	�٣�6�Z/5}/d���yK�O�h��Y4�����:�3�s����O�ϯ���%L���$���d\݉�M���T��N���ǧd�#�"c��	RW�TX	9� 9[ˢ.��֣�gg ?���Bc#�	�I.�>�u
�a4s_���z�drt*?��/��������G��ݗAĽ �O�d�q}�t(Cٮ���9����o����I���yP?��8�C9�C9�d9  �r(�r(��S򢖛��n�6��`(
�(����%�ۻ��݌���]���Y��e!!R��H��5Y��B����Sy�䙜�=����V����B���l2�!)�ؘ���6�X�O�Iݿ�����I��o2n� 3��Q�xő��+�(w�l+JKT=..^�˗�R*�ߗ�?�Pt(�/���	�²8�t�љ;	#�B��L\렧�Ŧ���N�B(e~ߥ�( Ӡ�����+��'�G�&�<���c[ɔ� ��4N\�>=��p-�,Y� � c��0� s�����\S��z4���X7�ۨƔ���O�h�3�
d�B�
�X��V�c b�+w��j��!k��5``[���(�ql��� ����d �E��,h��i�#:�`$� �m�M�����:��z�X$�	)yA��17�{0QܵQ��^bjo"���D��%� �Z��U�s�#w�}��>t������t�y[e8�����%�#�0x
3';�eS�1��c��|w� UX�������:%:��,�m�fس퉽[|�jr�jc+1x���+���g۳"� ��U0@�<�"*���J� �%2VN:�a�m+w�A�T����DǉX�˥�(�Z@����Q���ܘA�`gN��M�G<�L܀;d4A8b �1J �T�LB�O�X��ӱ���[z3�=��R{+�`��g�ւ1�pS<�|���`t�.f����wc'?�!۰��3V����e���1���3�� I��	���|�a��8\������%p:I���X$���]X�o��c�Ob^�R�`���z�%#��	T������n��%��>0T�f���9�%���>%�	?F&V)+=o�)�v#�W}�`�5N�̫��^L���*J^!~9Ɣ�������3+�q�H�� �#}���c;�������B`�n���y�Ș^E���p,��1���Ft�93�{1~�L�VN��ߜlȺle�D���)��)��HH8;;�����:M�U�M��b��܇6��9��s.����H������������a���Y�c 4�.��3�.�W�Oώ壏>��)<*�D�ׄ�H��s� � 4�$���hH���ͷ��ruuMo-d���s4�կb�����/�` :"��|����_R�	�F��v؟ȀԎ�ڬ͋k�q,=9;g<�����P���M���`�I��	��L�R:��tڬ��}�~��}� �Z��2	,�r����{�gXAO�g]��߆&��X��?�U�</�� �`r�kV�
���c��Q1d�"S����I�yQ;)Ja=c}�`�!QJ1����>i՞ufc��g�]��6�,�aO�R�y��R������8��-孱y]$�[02�O�yZyl���k|ǖk��jt��� ��O�S����}X3�Lc��Z�Wx�᝙ǙO� xH A�
<�no�ɬ�ϗ��Fv:Џ&C�iԎ�i�Ҏ ,ֹ�K�6�eR�Z�&`�y��X�2�5����<dZ;CƓ���׿�����{��O~N��=vv[>S���p��D%x&��q�1�������
�u���Z�ܷ��AVšʡʡ�� 9�C9�C9�?��,P�B��v���&�˝��J�fȢt����nF���\��xn��1	�͌�s���鳧����O�s�N��o����/����{���YѤ�;#o�=3F���)eSJ��}��1��"�e�F��'��@���d@�L��n8�JU��,�ru�F~��?��Յ|��O� ���|��a[9�l���S����j���ˬ����IT @ߥvy]��2���4��%M�����@(��B���o��7v]j��zq�(��B�����f�
�{��Jm
��~�z���|A�˜���I'�^��;��5�7��	����6k�  ���1F����A��dw�dY���j�յ3b�_��]DY������849/���i��i8l��T��@��i *w&���&r,��" �%f}�gA}J!PR��7u��%����qm����r��4���vho��=ӦoA$��
��%��H��H|�>߉��uit�@K�d�g�n5�����S�J��CFW�;�ؼ�,u����_0��:���w @��d�ek�(���y`m�"2��M��m\��̘�i�P	D?9�jF��USW��ms�z�Q\�w����$}�G�NW����ə���h&�0x�6#�m=�2l>� ���1@�@23�n�����{0��a��z9;	�"��	e��NaY �U���e&�^&���;f�'�X�� P�ԁV"�b�B�G>�`�eel��%�}����[BC���%�,�������y�����4�b��R��>_Уã��SbP���{��cڊ�	ex�c�їs���f,=�-�1��u4ү�����OȚ`�Y���+�tr�;K����dֆ�[�<�j1�.�d2d��w�24� �}9L@1�Rϙ7��������{Pk�[��⊒�+��6��bRe0�_c�4����[Y�\���`'����Ѷ3�Ka`̣�Z�+=+�1s� m�#����{�`X��#��<"�O�EL�s#���Q04�� '������0Hd�ژ�=b�i^qL�LGڧ�z�/���#�mv��K����-���~iA҆cm�����0?�:�ь�;L���p4aP��O��UY�?d+1���������2@���
s��'�՚Ab̝6�4�]��#V:?_�~�{x��&�	�)�%H��叠���2����3�,qc;�L�������t�\,|'d��4�^;&����'�����c��l���>��� ����g������X��hc�~8 ���AC�2A������g2��b�{��Ya�W8��v�%��L;n�lA�1Ax\��j��R��Y�;��-��˝�z`�����=ڍ�!;�*`��ݔsЎ@�μ�<���=�O&`�x6?4H7�&���Gc��x�'�XL� c~�!1���g�KH����>��(��D[[�Zx0l=r��a��*K"�6}L�k�>0ڿ�!iW�sϘ�Ɔ1h��.��n[�=``K�9uh�C���r�v����?���w�?��~�KM���͜�I��L�1��q�|�ˢ ���Oc������>�/w��������x��g�ɡʡʡ��� 9�C9�C9�?���3����=M��C0�Ym�G�̢l�	i����r��Ǻ)2�<��޼��������'?�?�P7ة|��<z�X~�O�H�²��6A@�ƕ�|B��e�[�]��>lE`�4Ix�^� H��oCCTfP��	�̃����bv'�o��Ͽ�9{򋄁�mnF��	*�[}�<��Qu�c�hD�,H�4f`��lY�d3!�� �����f�g�v��x�`�h��x�q|�o����ْ�>7Ӑ� ����+�Y̸��~�����?��f��U�O���=}�Nh�Y��H�`H�,[dP�W+�� a�:�	| �{n������E��"���!C1�]��K�/h�7&)�f���H�rc�E��Lr�1�$��ҿ�&oA �_.�ـ��m���g ��#p_��33T��M�A+�7޿���a���~P��z/�]jf\7�8k��d/K�W�%��㉫4%�����P�w('�{��=@�b$ -�ȼqA��f�Zw��(Wӂ�ny�
�%�A����!�����x 2hO0��0�&Ơ	j�3amI�z�v$�c���=���qr*Q@���F_6�أL�_�!�c��#�w��UK���a��#>e0ZI��N�W.#:� a��c��G]  �����H»�����7 �<^�<ڄa݇�P���,��$t��\�&��G|,2�e0J�L�����̤�,�v���x.���zeT�BHfa�,*�2h�����fm��д��<��V�ɋ����ӫǁ+�7��4k-օt����#���5��O�}f�__@��y��-�ń����:N�4!o�Ա�ұR�'�;���?��j�2=�q���z!7o*}��`��8�S�� hC��5��iY%���I�H:�zN$��I����u> ��Y�²��/u��N92�W� ߗ-�w�\�*9z\�`���hL����mR�y���_���N�� �?��i�0y9  (+U�C�C1ic�4�<�e�k�&��7o(3�p_p��X�e$E�s�>l�s
.��[��;�3�ƺ���V��tv&��>�I�m9�/>�\�o��sy[����e��b�.!s�����jǪR�<:���,4�� 3�>�{��4�H�|]\\���M�X����o��KY/��S��	F��v�!��� AR{U�x}�).�Y��,�&���V��, \���H�'��Jj{M� �y��z��^]�}��^�^I��F��ҹ炯��8v�<�!��O�bi�*��d�_��������6M�g�X0���蟢}�j�|'��m�[v�?c������<W�����@�(p��Eo�T<��l77���۳[[�� ����&����L�=Jw|�H�h�i ��ڷ1��?m��Aw��{�᳢O�z��7��� A�v��+���?�ccxd�tX�:� ѫ��e�anR� �}�R�Lx�+���У%�3Mw]c_�z�������8L6�>' ����x�6�9�^�`퐀}��ٴЉi6����cʻ={��>\�ie.o�(=�u7�O/�Ñ!;���d���n!�5б����G��~�m���~����W��?���r(�r(�r(?�r @�P�P�� �@ɷ�<}�����~��،�� M�02�0À�dL�m*�O�\-��jM�'��Z7h��L���윁h\�gP�t��b`:ƞ�7Nƽ�Z�4�FpHw����ã㑱O�����K��)yB����a_sc����nv�/�.�r}�V�8��Œ��[�>�g�}l��I�lll,�iE�,L��+ݘ^˝n�����F	�C������,ݫd�YK�ڣ�c�f@.�G0-�n�2����rA�Go�g�)�no�ˣ6�)��l��ک=��4ꯛ����2۬P�N:E�I9�V{�]�jP��߳T��	�潡�- L�����3���lr�7�%& ��$H�� ���4ƅ��r�`@!ۥZ;����1���DثJYW��]�U�e�~S�\��Ҷ��Id�M�ΐ�L�(�9i�R��H �T9I}�Ů�l`ޠ�7�Y0���1	������]��A0��x�Ta�@z�����{�p���_>C�������jύ !�0D�s�Cc�TUf~d{�bG����ƴ�H��g�ﲝ��g#�#`�|��çE�B7�3>�~�7F@&�U��V����x>�=���$�O����`�GC]_z����lC��2��8�����"˨U?���PC=�N���%�2I�9Y>�_�J��|o<M��Hy���)��I%!�@f��Ũ]p_����V�NJN�3zKdS�}��ҟ��Yd4��;����X��$tG������]�r��d�_`) �$�0�n��&�ؽC 6q@o��lǌ�L���3�FP~-f�ú��D�R%�&4����ds��5�ݙ<�W��u\�&����6��f����@��JnoV�ݑ}�QڃQ����@��Rcڠ��m&�m�犵6���T��V�w�.�~���sh�]��gY�,^��T�oX�hH�[�M������Z�����>�X?�/>8���d���m����D��{y�+����w|t��(`��K_��V�������LN7��{�E�.�zok=o.���Ūe��2���BR^�x�IF���w��\$	��DҺ�O�ص\�`Ô�?���`��Z:�F}��>�3FX�s#��H^�h{ɶ���n�� 0=:�>��ر�� |���L ,��7:��-e��~v4��g/�7�������O��B6Z��ۇ��՝̗K����S�qp�/����L%��R����Bݔ��	e��ρ9�^:��7 �{ �^�yIo����W_|&���!�t�o� `�ZR�s����'O8w�`���2X�1��� l���D}o#A`@3��-|@�ɿ3�+�����W�K�f�2���\yrvF�L����Պc	|:J$P ɠ������K�<��Ĩ��O\�>d�Ě�J �R
���~#[��k�ޅ/�]}�ӓ#����wߚ�e7d;�(�X;��#��g�@ȹ�}����^�cl\�hgXS� �b�������ҟ�R�ll�6�<�Lm���=��}ws�a$W$�K�� 0����@�)JJgUb2�6J��q-lD���h����>=̩-�_�W�IS��X9���$������j�`!#�4�[@�k6 > @���0xGaڑ��B�I���ki�]c��{}�~1����W�ָ`.s�ܶ;0;��X�~���%�(s�*��u�u]����#y��s&C��!�,͵�������R�y�������-�� t�ָ ����P>��Ǻ^��N5Ƒ���?�%*� u(�r(����r @�P�P��^ EpCKO7Ո�|��䣏~$�ф�Rc#�@;5�����dv  ����G4��{xD1�P�mΠ�z��!g��$����l�̠��:q`���)�����>7�4 �9m����q��I�1w!��Z��RR� �q�5d"_]��-��T'���\���?�T�3goY
m�&�p_�G�9�Qҗ~O7�����dˀ��i�37�fa�<
��.�^g���Y_�o�� [�I��:���Y��<��)]�0[��|�|�F��)�D���T-Z��0%����V��Df&6��6�y[�ປ�Z7�[��Wl@V/�g��բ�w-�8����:�G�)y`o@�m�(�z��[8&�Ȑ�b�ܤ��7�����̛��-�Q���w@�(����2Qqo%́��:X;4=/MO{�ߤB(oB��{�����o���{�5�1��������K�$xs���dfr�8@_�c\ - Q��z��e�m���!�����RK^}��hT�5�á�ꖽ���`����J�d-�V/ݾ���!��z���:&�gb�����/A�������N��^N�[ ϛmv�f�iZ3p�9
�q��0;�	��%�D���1��$��Ưw4����]z���v�=P!L��o����{����օ���ieJӱ�-Xe�v�/ӳ�t���9�l�w����Ǳ�t��u|Y�z]�5�w<��3�'����w��RoWz��d˜ׯ��	;�[ZI��[�����+��P;#����6i��|W�%Ǘ�z`���^�d ������$}}O��Y�������D����(���"��{\��o�sYoENk���c�$��'^y#��c�i7�mq'K=^����#m{^�qt�/?��;�f���.��f28��{M�����[z�$C_=�e��	�òYِ���Kn��rUQ�_ٲ���F�(�9{�@'ڪ��$@Vy����j/���}�ڻ��$�휲V�e|��v5<G��ܶ�c�޳��
�B�>༚H҉ ��4���F�;��Q���EA�4�	:Ʈ��4b,��v�(�����Œ��dr*��۷�r}}��K7VY_���k���
>X)�!au7���b�:A0~�C�k��+����C�
�?�� �e6��9jŹi0�f�:����`u�7c��X������R[�no���g�O���f��0?P
]{`���	��\s����M�Nǒ&	���z%���-w �cn�w��v��I	�%�;r|��'>��#y��;ΰ�?���v�v�d�#!��_�D�!�X�F�#=ad�A͞��ol>ϙ�@�Y�`�H4���b��[8�z�y�.ٚN�ZA�Q&����{�����K�c�@�e�l��� |@�úl����R5�{���l�c��;x���(Ώ���,�#��R�񙌵�&ٴ2���y�Ɓ:�j�O�O�N
u�ʹ��e��v�}~��%�Pj�)����S�I#s��e���i��]i�'�E"�/��A̱6�dl+XOc��6�q��Q|Ed��H�[��,[0? 1j��[	�kH(=�9����˼r>t���ַ��kI.3��g�����?���7��w����-�Cϛ�������M���CI㾮�vM�yM��y�Ъzh=(�r(�r(?�r @�P�P��^�k�&�Aj��N�,��E����"�Ago~\! �)�Ȓ��4ED`DyB���؆/Gc� ب"kl��̴�zcs���{?d��f���Zs%sf�Wa����+���$�+n`׺!�/	X,��{J0 o�!��$6h`_|��g�홤��Ǽ'dVZD��b� �.��}�;�ȦĦ8t��z���s��hl��A��`ӰAgD� �� W�䊐�Hc�$[2c8����.������Z�;	�1���v>�;dg�q?�.�|��@
���R�i��y��l�!P�^e�7&7�X���r��-�-�f&[e,�;�EH���N��*��6�
��}{�{;��_~h�CP:���d3�)^�&�d����k�A��I�jL�Ej0�a�F�N�+p�SN���``�C��C[��8�����h<��Kl��9V�`Gy�Fb�Gq����!9
�k�������rr!�����<d�m�R����3�%3_�yz���|���gu��ݯ#Q,�4�3�Q��H"���˨b0'���ڧ	~����ЮLgނ3�gu�Ox�D
���k�<E ZA}��; 4��,��<�Le�<E<���.�� �BS-p�"C�!��IQK Sp��H�� �]��،�!SSh;I�^���^�vB�@����l���)73�~���nN����3}n�����z0�E�r��u���פҕ��M
�m��|(h�^���TRz|؛T"���b�^��gʝ7�,���Jו,��8תm_�]��%Т��l	�@��~_�~6ʡ�F�e<�t��(����Y�:�����s}5�䢴�@V��/ ��N�p-��:W�r|6�6=�M����]4:�.g[�����/��%���+�߾�J+v29Ej��]-��+�?�NdZ������@ʕ�Gw�W�����b���7ɵ��%�{��č���r�9����ܕ���PZo�vx`[���cD�<Uv軔�s�pR������� JB���{�Fů_��Gd�����`%,٧�7� <� fZ��\^]��奼��e�t��	�F�����公����L:��[��#��(�q���o�ޒ¤��ֵ�!m�$:n�)��UĠ���N..^�<�w�>��{O��#�����F�39g�>�( V����]~w!�|򉜞=�����1� ܡI!	���Y����?����>�X��`����7�_�r5���R�>�o2g�K�����������������G4q���2�7��;�^����B��ƪ1Y��` e'"���$:t]������	 �B��-���=v���NW߃�K�3�d�m��zCSu�C�yƄu�b�M�v �qRS5�-P�XϠ}�zCzw5ނK���z�t!�*�qrr$��D޾\Y2��}$��*`������~8�6c}8�(vDg�Ny��P~��4��#�ak��0M�/�bR��])Cnofd� �2�1���8�xܧ���ﳮ�' cX��h��$�L欧�#b;�W������>Y�h'`��ٱ�LҎ{~��^Z�Y�Z�8�&̝���lX���/R^+�(y���f2�t�ꛯ��O�m���Ð�|62�n���f��J����D�޻��Sm�^�C�NDM���ޡʡʡ��� 9�C9�C9�?�R6�����h:" ��8�5l�N�
�N�o�D`Y��^�c63�����Ǎ�yX��l��e�Ccx6����v�j�F�@����glب)�ۦ�����3�G�̔�26x(Ϟ=���f�\�_��W��  8_-�^�e<)%��������ذwh���F�Oij�o7d�f7� A����1���e�Z0���b����|0�NJ6���~��ER4�o`H�4�]�Afr�A/�'�7��ɲ�����Y!�$�Z�a�Y������v �dˌ��r�n� 
7�A@���a`��L�L�v�@*3	���s�D OU��ӈ@U��Й��}�ފ��U N�o
eP�>$�a,�<�aE*�՚>��e!��PT�#�-+��w�fF|k8<��j����Y5�[m`��A�>=�)t��.��'�L�fڹ���3 ��Ƶ���q������@��E{ͪ
�r%�v-���i���^�ɍ{���y��$z,��b��w�'f�D#$Cvhj2\�v�8���sh�.-S煬\�m3���L��t�j�W�?Kإ�;���	"Ʈ ����e)��V�t{��w���e��l�ޘT�����w��Y$�E!?���~�L̶{w2}����Հ �F�����&�B����Ħ[$fJ���*P;�]~'M��F���0��!MY�u9�Ȭ��VP�Ct�(�s��o��3��H�]���C7��c�M�$��c�k�K��F�{�F�Ѽ��l��I�1�/|��	n �F�}�}�=2c��~ndh�ϔAy�buUeFF��?�&����� ����r#�n+4?_���� �����x%O��XhF^Ꚑ/�+10
rI��)�WaB�c��[`n5
>[��@P��r&秅��L�����L���^�'dh*�+���)�J溦t��^k@Њ׫t�(C� ~�2�4)�f�0"�GPt��^ ;wv�H��ۑ�|)�����Fn:�L�L�S}��Lx�dA�l��b$rϤ�t��π����d$�2�&�����|�q��k��̆-��f�k����&*"�SF��F6�C��f`��`���/7�s5�O8��r_�:�9:���\�d�ǔ�"c��3c���yyz� ��9�ӛ����C9>>����|��a�i:�%F�:�?�=]S�2�oL������õ�#��ͭ�΅��c?
�M'rzz*��z/;�/�S���l�}�'1��t-<N��_0� u9���?�\�-����\����|U��`%@X	�ϣ/��_��r��=�u�磫�Ky�����Gd�p>�lnX�}A:��ѡlm���o����o�-�-�;����@���㜆�Ϗ:��%��	�VN���%e�z�l�)���I��� �1@����`>������zEd�B�
�V�� ^�� 6��4�',yi�$���}V[�����_D0
����s�<�`�����>��g����}瞜�y�{�����5N��3O�Q�z�0)�fbTnL�W'47�(�I������� =���3�A�-@s �sm+�����G��o�������ͤa1� d5u�!��V�.ۻ�%	���hy�v�'s��t9�J���,���cW���(�J��eJ��v� D$���9����군�E_�xC2��2�H��	�nޜcf㉎�}ޱ�A%�~~9Z���a9M�|c�k����J�W#&Ѵ�~�qG ��C}Æ �)��)��l �MٔMٔM����U\C�s;�SR
~+=�!�#cRX��L'#9�/��[�����@��Xߟ-y�>�rKZ�5���6��6F=8�4��1���L6Lqo�+*�@��ʽ ��@�h2� �&��>�����>���<~���|��c�~Ĭ�!\l��F����3f^� ��4�!C1�uh�:A`s6���WrtxDk�s�D�%"걠- ���\������vs�ǎo��Ρ!92��P�,bh�S�Zh|^%�$SA�����<4�3��?AÂ�sڅ�fݧDn�Th���  N J����=�ڑ-=�����^%+��ło�#�z�������e��3�ϕ��gx�,� H�9 %硼�w���g�z�? ��>�kvIUY��P���l�Ҍ�AX�B��80`KM	��/��J��g�)��&͆���!���,J�`��.l�� �5�3{���WyƾϿ@����������d-)5��:�j>4��:�H�dq.��� X��2_��B�w��!��~8�es`f������ p�=�k ����tA_33��{)� W�\�&��b�NF��5��;MvdNӔ����87�k���5��>����f� $@�n�)akK2�Ȭ2�P���}3�����=��*��	��İ���y�bd9|���9��U�t�����o�{)=�#�^��JU�2��Os�R�muY�]Y���c�[Ci��	��e�׿-]��bݐ�<�g)Lڍ"��ףrzL�wl_��54x�m*��K�s�̌=� ���n�B��r&�˱,���� �?�j=i_�)zj`
���=�9�r���K6��Ng%��S�u<��C��[�74��tj�ϕH� �0.�"��ŕ�_�@���o���y��B�S�`yOn��gI�e�p-�֡����h�~�s	��z��/��#������O���2?�|��hg0�j�4'�i`ZxC�F���ZR0��@#���0��0`�d��m�X�)	�D��d�š�je��p||�k3���lmϵ����#�����d� �]��cL���e{8ທ.����9���"�,fʋ��ǩʜkb��^|	�`K�����K�&`���%@����52ҹ�}K��/��)�������깯y�����s���X"�?��$l����^�x��=<�P��\�p�-gl>���0������~�ky��k2:�?�'�N����}*_|�9;;��$�X琾�~�?=�y3#����{���7��\�9�}f�����t2˓gO<��:���@�F�K��m}�(�:�0�eb�/�+���4����2  I�r����� P�{���_ȟb������/�((hq�u�@��)���p�d�kd>�~բ��o��WZ�H`A�������k$��k���hqɵ�w���t`�X��ZƓk@1�k�j��]�2q���ﰞ{5;��sH��N\��BB�V�C��L��$�Zڟ��j-'����f�{!���bƱ?���Pڽ��O��9��m����C�@�u:&Ph  |O0��=�>ÜZ1�쨘}�j Q�gN��K (�>$��TS��������Vb����G@�|�|�r.wY�i ���4#c|��?�S�x.��)��)���/ dS6eS6eS��%Փ�@G�ȳg/����d�u�4͆��ћ�zX��,��)H��`=�p�A�ј��v�M�����Y�%�\��7��(SSTk�-f�:�p�[�`>��ԃ|��mH3�$7�ld=z�1O���>�a����y��5�8���)(M_[l[�g�t�qO4+e�T\@��1�ؾI��?{�L�W/���!����'y�`�1)|����Z�W<l�4�q8'kV�EL��|J������	�d�R��L���S�l�.�`�,�%�Q,s�I���@����s�M.���|�W0ڮL	���ҍ�A~IC�%�W�C[�d�������6����=��4r�������U��$�PT9�U ����n����{B��R��R�f���I��y� � ��fz�:��{�� �K_�A���f��p�B}����Wd�h����?�#�k��̋&\K�����Km�����o`~��z#hBP̧�YU�@"��`��������KJ�ENZ�uW�����	B��~�C�Rg�b�e��-�{��-�I#t?4 #p�!�s�'Nn}��t}!��䰐-�5�+��k��t�!�N#jC+�ٹ��Iw���Ͳ@����c^I��
�mP�����L6.L�V:פm�wn�P��Ǝjr��T��H�촐ٴ�nAپ,�R.Nϥ�����t�nC3��b%��
����l5�i-�R�����T��+t���������|�
<b7���c�7L�+���L..d��y��.<8"������ v�� A A��ݙN�k"��0_8��v�U��,��'wr�ֻ��ۗez�s�k�s�D{�j5#�!���%��=L��1dvL�/�^W�$W��X��$��Ȳ�� ���īV�eT#�;���։L�Vo-������ޯ���N�0��ly�ܨd�S�������WϳlzρM�>c=�*�n#B�	�"��dvj �`/�7 ��]ӗ~�/�a�2T�;�z�ZH��+ Ϻ�d"� ��c��m"e���䙮-( 0xb0qY�[��Q���1>9��L(���/��5��Z�J����X�q���缧��~`>��;"xv �XOΎ�������; �dz%��O��.�2���0g��"v�t�u���|��+����!?��]߃D$L`��ɣ?}��B
�����S9~&�B�<�V�UϵoϘ@ϫ������ū�\_�|C�-����O��a� ��TZ.�oO�<!h��'�0�F��Ox�}����Ϟ�b2a ?��; %����� 
�.9a���Z��� ���}��#>�|�g#º�@^ kK�EƵ사A)� H��''g�w�YW�	���d&_<z,G�f����恦�
 ����S&����y'����Qz�5h�����'&���)<���c�4b�XW��ѫ$7ٷ��Y�� ��,`�Z�
�t���������@�`]�m>_N�N�2m)kFvMLY&%��-���7%�v��ΐ�2�=�) ]`�`��f2c��g:??����` �U��A=�X1f��ۄY1������X�6h�L��TkA��o��`zc�b�������ߑ��6�r�?yE&��)��)��l �MٔMٔM����<]g�HhxM=���ٷOx�!8���;�z�����xh�Då���i7�pLM�(�A�f�g��j�Ng�c&���/��$�?%Afq��x:�C�-'��|(&?e��)L�3�Ȅ����\��FW0�0�˯���9m�̲Q[���`䕴��8܃i�{���W҈_|X6|�3C_���&r�����?�/���L��ԉ,C.�#�0��W��@6nfA � I�p�fdAvd�ҧ@߻���#13T�3�0�o1s>s N�qd��8��:��yc��3���Y�����AR�cx2@��f��r�w�J�|��p���D��t��#��d�j���#k4�KĂ��u(�����0� �?K��8�����A_;*����4�E�}�> HU�9�~���N8�G�vP�O�AD�c�$>���>RZP2w{K��,Ȉh@?���]a�d�>3��zzNn+r,{��_�1��V\��Da��-ꁯ�3WO��؛����5$3$t�o�3>m|g���5k�(oH�U7�'�,��x���)M�F��x�Z.�rc��(/k��t�8�G����גW0­��`~ 8�����1��8q�:�z4c_ԧ�@x������/���S�y�S�I����H���W��#�[����*E�g�̏�?�C� ��S,*�@
'K�m�\�)����q~��ՙ�����ע#[n%��7�D����x���D�ij�/ ���7 7���� gd�/��2��,��k�&'�O6兪�ϋ�	�V � �2:k賌D��:�t���-\�W�t�O��Àui����R�~JdD}m�9"�Rs���P�G�r���J�p,��G�v�����2k*�e�g��>+t���2��EF�c]����@�.�����B*&�:-��DL٬ݡ���:�ZK�L��� ��Jg0_��d�U�ru��_z�#��x��>z7p[�SK�'��C���6� t����RX��#��|��0�����XO�%j�7���J�![�[�,�Q<����?����[���+@!o�S�ʗ�?ܾuK�.Θ=�����$�����T@6ri~c��l�h��r쭒�K�̨Ƽ�2c�!���AK�é�9$���+V=��;���/n��tO��gry%���᫗Rx5\Q
��~�`��jʤxr]�g:ާ���	�O�Ѡ�0�?�3��4�/����ۯ%x���ru5�]��Ư¥|�sX,�鴛\��pq~ƽ������\��7�ܖ����F`
I-�g'��,	�t:�6A�d�U����SM���B_�+�P_�S�������="X.�3/Gc����@�̇��]��fzo0˞O'��x��L�J�6�輐�oAr�����Lu��Ki6���ruarXc}�L���K�+��y:這8����򸯬g�z�0`/����t�P�X�"��0ύE�!�$�q����ji������ þ8t��P��	�<���}��ض�>���[�S�V�a�5)p�lEjd�K"��%1�`�����nk�x�Y!֍�/��G��G���n^EQ&�7�4����:� ��3'�\�	@'���bN�@���t�f3b����fC�S��������ށ���M�i{���(��)��)��}+ dS6eS6eS���G~"O�>�V��! �L�gϞ�h|I#�{��H��SB���<�A�z<�Z��-w�ޑ���ONNyx;׃���o\F~@_ho<ؙ�4 ��bf�e=
]�Cy��&��L\�e_��U8��� I���i�6W&7����$*��H\/]��1���0���PZN�t��d6s�01�d��c`qq!���J~��˯��r��j�#)S���=��8��/3 ����,�>��J�&y�X&���g��̧C(�z-23�%�B0D��4u�����,(ga�G -h����7
�.V�s�$��{C�gp���`���x��/�,���� �����4�%�#`�+�|�g�0�C�v�Y�u���M�*Xk�{�8�!{�~�`|��2Y��|e��g`�H�! �zB&�,zo�N����b�ެ�²5����N���&�<*�_�5S�i�&�Ǚ�Z1�a.3�	F���*�	ԀP���h��kfH��Yx�'��82@�ZV���Jfm������V�d�|ب尲���G���Z���1y�� ���v*���m�p�7�!^�����s���=�L��&�$bF�5�G��v��$�0FVnn1`.�[���;���,Xf��^�1��J!$�
��<q�5Q* άb��oy
��T�އ��r��%2�%���[�1瓆�_N���tz�����'��E"�֛�x�I"o_<�Er�s�O�+���� Q+%�"n���E_�w�,�u��M�6�
�7��^����:H����@F���\փ����;$��_�du�
���ՠH�]H�m��M��)T�3�9�p��$4Aǽ ��m�tmJ��활�IKt�0���@>VQ�u����H	#t���.+r�0wR^�X��f�g��m�n�Ec���
��Y��N��/`Se(��uo����G����)��^`�[���t�����6)Kg�d�u{)��t-	�`��?g��p:˜OT��@�7j!S��04��	ǝ 1���솜�� ���7Q3Ҿ����V�
�αaP���~�����n_Φ&��y�}�Ŝ�X��>0��X��ِ�kw�NN�c����*�a����WfsC�*����e֛Y"��X ��ܑ��znC"��d`�����WT��,�x�.�3�h��^�&��;���B+�Āe��<ר�b'�OUۺ������A�Y�p������Xǽ�Y�,-���Y��u�3��<M0�1� 5F'���T`�f���������K��o���A���d0���N�5A{x�ppk��\�)�L^�zk�4A�����t�$�Un��;����}��~@ɥ�Sʇa�5�-tϐ��I���oJ����R������
2x�@"�`�@�	L�C��,��h��X��m�v��Ub<������w f�e�?�z.�d-�F�08�	 �:�Ʊy���� ���=�t��w����뵫6����|����VE@�ۺ?A{YbDI���;O�@�fS�e��!�X:>%�v��m��1��!�W a{5��+�G���a������(Ê~ؗdXV.)�fx�dJ������ߺE���������0u:��^{���my����?�	YUHj
uL�E�vص�FR��)��)��}. dS6eS6eS�C�N���!��PX���ċ�3=�^��!�^�Ƅ�h��׃}������|�<�A�{4s�F�dˌZ�й�AF�%�$˄ 
�/^�!�2W`tu���H��ǃ8�1(A @�FF������%�A�h顲��x��i-R�( A8Hv�]=\Ɩɟ�zX�(3��8 �����_����?��|��K�K@��wA��2�4�Cm���	v{�	�X̗zx�k�j˨t�;��0�&o�Y(��L&���ӵd
$#pϕ.�1��)��|�Ӵm��o��a��ʂ�3��B�eȀX���T�O��B'[��@ :�����ދ�A�!]h�~?f,]�ɏ�	NX` ``i�CR+����r05L�ʂ��X�s'��>Sg΋B��<�3b�,yk��[�W`
��<�穙���Pf�]%$v���P:	���Q�u���2%k	ٿ-��,� �Y�Q�Ȍ"��>/]��ք�K�X&˵�@��[~�c3-�G��VH��rҤ���9��,�ZJ���{�"�hc�L�˯jO���kP����nH־	� ����Ռ� �t6e ;&�P�3��bVwjr`�3�-����p.����s\��^����#MFZ�l�)V�?Z� z�i�{�16���8�#J0p��Q�uAu"��0��c	�HV5xD��T�$�O�����dۉ���[���)�%�g��l��ڣ�3�(X��4`o����d,��X�u�Ւ "�������8ں��~!]�H���g`@�����&�6 P�y�^!�Yl �=]�R�MFM����$�����=:������ځ���I�����F�Q.��m&:��|��|a��k��Xk���&Sl �BX�T-�i��b����Z�(��x��	,�
�Щ����n ]��^ 9�
��| �^���n�3��m�N ټ�d�0����?��C����Y �uI2ׯB���`;�ص�l@`-?&KYK
b}�T�f[�-]o*������,n3�F�|woO��>�^W״���;�c��fԢ6|?��@X�����ߕF^�zq�����d1���]���+�$
NF�;X#`_�3 k���m9?9e����w�H�e�G]��9�k,� �b�9�b�'�F�qt���2�9���vy�=b�Ȍ��`:}L�����|`	  J�E��������ج-�k�O�صSBj�� Z ��u���`[{�L=3��,��/)R6j����"�Ys��K�W�s��1�����)mHs/�{�)[ڶ��'�/��z$��+	��*[r�F����-a��L���aN "����� 0/��j<��w�{�6���裏�g�Ɨ��u�ѷ�>��2���Y,�4 B�y � ��H�X�$�<���5���
�����v�c;��i
v!@1$1 ��39I�K�g ԂGK���ɮ��{����rC�x�%�`OS���%n�X�S�/���C�G���=��\��E��=�?�wm�+�V����є�?80����C�{� D��w�O��1�:]��m��ػc0��1�3��4u߳���/���`�`����i��^���{=�1$��ܿ/;����歝m�i��g�w�]&C�W�Lȷ!a����Ϸ�o���6��W�ziQz�d��!|hnʦlʦl���l �MٔMٔM����|��7��8��$$���T�X��4))Ѱ-w����MJT@���8�" ��3<-$�͈4+*J���D7i�p8CNA���dh��r|z �Pb &p8Cp��.c=�97�4J6?�<'{CVB��`C�ݓ^��򮖩I� �>��|�;N�|Fqx��+1�m	���H�ϟ�L���s���W2�)���Aa0"(��1�Z�}VX������x� �����#L��pĽ(�PX&"
������� 1���?�jf4=w��z؅���Yv>4�3�-k�Bh��4�/�19����,`�^�&�u�C?�A)�Wܓ�q�$��#f26s #�$�H�m����5�@r ��nv��Re����,�gf� �9P�e�;�C�uR���A�@@9���ꐛ�a�+�U�H-�k�� yU�`^�צ�<�LV*��G�;fI���~����6�X�8|ϱ,�����l�����\��B��}�X�m�~:�`?�A���4D�s�{~=�s�4wL�J�A耺� []��q�莵�y�"c+������q��LE �^<�O��#��C�= $^z��=˞�{��y��3S�F#��yYب�o�3�L  {[M���K1t�s
l<y���se����Y��Q���
Ǟ��B���BEP��/�(�;��+���3�M�:���4��D͂�h.:������!s��,��f��}'nK�ٓ*4�A���m�l!�?3���1�&r>���L[�|@:���6#V/�ʳ�CV\�Ɉ�� ��9u��\�_ԍ>C[�c�2Z����m���
�_�Ϫ���w	�L�������X��tl�!��"K8g�>����pX�p+��%���%�������=J�鼘�*x� �y)>�ɰ�`�kA��0�
/���B�V� $�R~,�DqX��I$��:W���u���	�W�Ƈ���q�.����1Ъks�Zbm-��(�;T�[˦�8+����Ӛ�e��J����;ea���`ni۴�]]34-�k�]w*]�8 (��q.-VZ_�I5&s�^���of��<~���z��d�@������3��� 8�C�t-!#���M�2X���Xx��z!v��³k�Ly ����n���}:N���\�՝�mI�zݼ6e�z�~����\�Ŝ�c`<6&��-�̃�󍥆��)���.?6�+p�y`�J�l?x-ed `Ò���;�*ꮴ���ȁ]&�g�'���vC��Gn����鑁�����]_*p���>C� ,�É�A ���x�^X:wv{��[���'w��%��g����X��Rb�!K�z`�w����ا̤f\�O�0���B&�AF�<���Ԙj;��hڏ��cߠ���X eƵ���w�)Ǳ�N:�KR���o0�<�늂c�6؞`�@��:����c���{�U!'Ev,�3܍A��6o��|�9�~dҡ��/{T�C�=|���Ξ�C�S�����]���ډy���D_���t��3�"�k���9�d�·%�F��`xl�����G�y�{<g�4�9�C��cK?,`0> ��eh��>u��$ ���Ku���8
�O1B^YƲ)��)��)���@6eS6eS6�?\AF$૱��+��r��-�o�]���zd�2��a ����T��3Rn�P
���?�\^�~eRX�A�@`A��j2eF*$��ݾ�+�Lg�pk7[<�גJ���Y <P.뜬���8t�g]��r��rQ�8��N�m� p!`�і �N�џ�<�V~�/������gIN���!�GqP���iK�y��T�����@[�	�Cj��Y΃7�-�����&����-�� $�HO'���Ӡ	}��Q>a&lE��.����~@��T ?�7 `��  ٦7
� �<YP�[B߱	j�b�`��3�xR��6���	Y���G6.�x��^bW�d�(s��#Ә/��I����gD��\� �L���= �Q�^>��)����`�������֋z�"&���V�e�.|�Ư��*�d�NJ�Xʴd�vAf�8�R�@@ ?0)膀J�� �.Jܸ�[��_�{�ydƀ=�@~.�� d
��qJ9�~��x�)�a���Lp��]+c��Nb�� ����3��{F���W%N�^o��f��K�ߌ�ݳ���,�X����
E!�
&��^0�� 2��ӟ///�����$�f����DC�l��2�:i�0 m���e ��e�{�	(�d��Ԗal@�! �k�0�5R��aI?�n��TS+��gD��/�}�֮�';ҍw��I3:�dt%�Ҙx�hT���B�Bz�XÁ�[:뵠�kM��N ���Э	�8f;�t>Du 	��<�D���O05�Ͻ/4&�}NJ�T��}���U/��Cd��צּ19`�>ӹ1���nQW*l%Үt^�g��E�V��~^����˻�����cm4N��R�v���������<h`��?������^Z�B��"�A��&�,穜\�g`&w�]�޾M��8H8~��x�yE�,�࣫Ϻ�v�d���
qt-77�5���y��t��� J:�{�1<
Y�	�Dǝ��(Z'��Z�e��f:�qe���6�Y���s���� ����V���^�a��/2�߾���#����G����>e'���k�LN ��RV�R�ŗ��$��nY`U�~p^�,Od����������[4��^]�{�/o^��|�IR��ʘ�F	��
�r�B�;�ؘ�P�΂�<�s�XPc��N�d�ZðC���,! P"@���Q齬n�&�C��s a�8�
A�u��_�L9�阌��I1b._c�3&_��c����L�\k��/Q�P�D��$��5�RC3�# 70��'�3�����,��ki��#��������������666l���X)=��p/�d6�����) Go������(���󚓏4�#\�%lm3�dUڞ���_���>�x$N��0%_,�oX�>/��ep�sq���h����Us?�����f����6F)��H<iD�����'E�G?��z���{�>�N����|�1�%%Tu5���\Nu<�z�}+Y�e�|sR�����_���W��շ�~K@m��g����&�<�ec�V���cc�)t�F���312ݏV�yquy|����z�m��үڿ��/������CٔMٔMٔ�m�  ��)��)��������=y����>���]�������� �nǲ���1%(�Z����w�y��d���7o�Gp1BfC&k��GL2k�k"�.�C��޾t�<U-�Tg�#�N�7��;z0���*[�D.��/j&Adz��`���u��n�t�FBP�����2��~����_�_��������a����W�P������� 8z��nz��ڐٲ�`��DF	�L�Ȏk��Yt͌q�(����Py�7�����#�i�o�F�J�>���'�w\*Lr�� P���m���M�^�\ל�d���1�ɬ0ȯ�FI?d;�0:_˪,����Z�/��mFI'� 2!:��3� �%}M,J�� ��U4�N	f�`�M6�Eyۣ�<c���Gn�Z��E�s��C�4.��͏~��r�$��y�Śq�,������|��t�+��Ԟ�e��Nɜ���.>֨��ȯe�zr@TZ�Ur����� �Vn����a�}͂�d�T��̷'���g@��@&��# ��뙭+� �֞(��ܞ��^h@	�-���%��?�Ψ
�8�q ��Cx�;u��5�����!c`:%��z�8[%)�=nm��;�gv��3�J�|�2~�������nįl-#������{!X9oO��O�,d �-m����-�����YSZ�	z�4�į"��t!���]���-�8�@�X�����t���10)(x�����o����δۂ��w�&S�w�s~a��v�9<��t��[���G_�{O�q7�Ǉ�L&�\�R)����a���������hm�h@�]��;ۆ���:�'s\�K����:Ǵ���2?�k&��2�n�˓��Ɩ���}����1���ė��T�}i��W�w��C_��\z^F��r6Ҿ�l�����Ȃ�)��9U����
�kK���#߳��r���s���e�Szp�[���d������@ȵ�2�!W�5 ���=i���M�1jI%�� ��<�y:0F�:���6%���峧������JN���br���*Mn��Q�}�|gB��}f�7�}��a��"�yH��Y�Q��Ku���xk[�:��}���?��������y��^^# P�y���N�`XNt�$��~~�� ������-�b�[�|� ��k:�o&C�(��b���&�X���W$OtJ21��B�2���|c�p-rx��x����h^�u��L )�xǾi6����)��B����lV����n��^)��w]����������� ��/O�<�Ͽ��Q{Z�Hf!K��ha�����"&i<�G`����`^� <@ȹ�I�X�~��:S0�K�C2ocʵ��m��U���ҁ[u3�[����0�=�����M�{x�tt�k�v��2YJ[ۅ}9�=VLo�� <J��n5��m1��:P�@�P�U�������'��]��U	Ls�s�޼~)������K&�$+�'[e��A���̞�'x6H�"�^,�}����@�}�A��  DA�E���ӆC4�)�'�οz�o�i����tg*��~���>w/��lʦlʦl���l �MٔMٔM�����3@ ~�@�wwW>�������<��Q��L��đx#��>��4�A�?�!��'�����0�T �M�%�v�7-�L�	�I�`s���Cb�=$.L�7�I2�𲀟�����pF���5��J&���C��Ζ�qC4��=z}��g>~����?�����S��Θ��,�8l���b���9���lf��>�1*fv������ PYr0�z|&0" �#P��x��yy�e|"s����hh�|�oR'��
J2V�)M���}|Z�Zp/"AO�.}=H�--��^)L����X�,���E����F�<䃵��n��<�pV` �>�Ə]_����J��	_�:dH�ޖe���m=��dQLޤ�RϿ#SeL��ع��ujh�f�k�!3���k򳢐����(7P c�pF��%��u��&��T�>�aI�����$Fq:% Ӛ��!�m90�<j�#Ȧ/Mf�%��7���	L�<��Q,u��5_�2�Ho0E< ��8�<���kp�b��ZR���s�A�0_�}�p�ϱ�G�#�����ݒ� I0�<dN2�&�)a��7D�M�'e���3�(;�S��֝���~=��ؗ[ݹD4�19:�Wu��Q��*�Q93�k��o�9̂h�:�����b}����*��<�Y>�`�糵����DՒ��I�M�*�p��� ��(�v�)���V��cY,ǒ�;�c�)� �Vlf�P�f TΠ���34/\�8��M��v��g��WV��]�[  ��- 3���i� 4Bk[Ë̊�6�ۇ���6�3��Z:oC6.]�5�ҧ����FA�]}/����2�ٴ���׌�\-a�<��Ξh%�ul�c��R�����3&���	�=@ >��й>�7�D�ߚ���4�[�S	�-���[�5(e�-Z.�d|�c����+�dU�_6��[l�׬:�k6@���}��|P�D�6��F�@k��>��X�%�p�PBfacn<==��b%�~W:�>J��!$��w�e<����HƗ#@Jc��-��5t4�j?K�G��>�������Ľ���Nh���mzh��q��;�h�m�ɍ��x� ������޿ߧ�W�ѡ�������.c,�X�����>��KW�_G?�|����X.t�1սC7��st-h����7X ﷶ�)��6K2�䊐|�fD���d��;�}�/�KR��R�.0/�.k�A]'�	X�A�d�,��`=Vm���i P�=�)_r=��C#��y~z"O����G[��I�0hOt�*������Z�M��J�gh���ky���k����T�|���ԇ_�ٜOY�� H�-�S���BE%�|x�:�MK_-�IS����V�I穭	0dǊ���V�*8!c���_��e2/
����0 ɾ
������_��S	�J�LMǺ��Hq����Tw�w9�!x�H><�dB�U�q֏"ߘ������s x	L��V���Mz�`�[����ĺ��1bt.{�m���'�>��`L�G�+c�6u��ϤI<�^zM0�P�`���׏��씠�����{�CpǏ _�!p'�I�e2׮h�)�{��*�(I����_]���� �}��ﷵld�6eS6eS��e�lʦlʦl�_� ��<���]� �)\�����o ��������dK'wd��LU�e���I�|�	���T����F��H�qQ��! �Ђ�%�4Zz # ��:]=OM���,!� $�d����C-�lX<'�w��7��#�C^�����)�����J~������1�D����و���Ȅ�,�ʤ6�ܴ��@�L�p-�T���� ������2�M�L�Qe��O��$��̅��Lh$m�"8�#`�;	�c�|Y��9���UU0�v�^E����ĕ���.\ N\0�dF<X8�f�$�p���K��"�c�ωv�Y����'7����l���~l&�̲�Q���z�)�9-j���<^k��0��K���.�!K�]��:���b�:�]��H�H&��dHz�IgA�)���r2�� �8=8�/�ZELv�E�<�Y���|�v�0�efG ��y͆���0)#PD,����,^�@�Wj`������t��A*�v��Tf��yX�u�"({#�V��
|�SL��m���lR§U�m��3�Kq+f^��A��2K�X��u)���۷o�Çu>����\.�_J1/�7���9� N��8l@|&�S�9VN��p��`k{����;3��X!�>����e����J�֖FgUn�M�'�a.��%it��yi8qeA�����R%��D� �Z�����L��D���{\���px��>%R�e�O���Whc �yP �W:@ώɻr�Hr��1׵$�O�+�m�=(ز/J�<K��T����H�)�$迁2��B�`!yr��i�"�`&����5d&Cf�s�X��ҬT�
 ��3����λzc=]���ː���[���X03�.Ȅc���NS99-����9�+�	��'�ͣg�����:G�[��d^"�}�k���yLv
�����}���ڏ�;��UL�^L�	��4 Ō���O���9�O0� xP�I�c���{����K:_��d8F��j��{ !	+��X�r�E��vȂ�k �s��]�����K�k;g��%�!s�i�������{�]�˹�"U��'�,gK9><����epu���!���~D����2�zV��$G���I�Z2� �$̮��3�����7�;<�D�?��<��6����#�v�B#6�l�Y������z�0?r��&ݹ[���`�`����=ʈ����8�d�����IZg�\�C:W�Z�������o-O�}�{����G�l�3�/�jr%Em�<l�]�ǟ�k;��9y�����<{��{��G����b"[���Ӽn<��CL�L�s =&P@K�&`�D�Zs�W"̧�t�����t}��R�$�� ��ʢpu�Zx�z?	JHQ�,qL{hT������[҉�L���D @tn�>��9,ֹ |��^¸���}��z�+�L��ɚŖ���2�M�L����S�K�Ȋ16c�aI_"���Y%g'������գGr~x�u��L�(ahv��[�����O�L@h)��o�6����H^��r�D������	�^q�к�����~���&#�/��ch<���ř�o�ĺ����MٔMٔM�^� �)��)��)�!
��q�C�`:�0��x@�
���y���yIxt��3ݫZ2��H�9��Hl�B����˳���ų'r9��p� ��Il���@�|6'� _��dA�>�v��Θư��Tղ\� v��f`�����|��B`��|@m�`B�-��!���S=<��g?�_��_hv��*� xx�Q�d��1 mjxU��*����q�����>(.��`@���q9^G�p�D��:�ǚ�&�,�;*�'���md���I�2R���<�Z��[�f���~�̓�2�����fl����l�:&u�:Lĺ6�j�f�+�%�|�-�'f����$�,���F0mxz/yA�"�*P�7)f� J���\��r13��5>�.v�� E�2v�o�����\j����T`�k٫�T�;�L�.�e���uq-��h
��L����:�VԠL�/�R�-{��>s�Ȓr`!�r��Ѻ-M�ǥ�1
D��;z�5bR�!�,L�7{(��xJU�5�����F����g�N���.)\��H�c��׷�\v9f�C�/�EϠ�v�M ��o-��L^_�jw���;������>nY�������L&W�l7e��x��Lݷk ����D�ژs��ͯ+&c[���E��sƞ�S9yS�x*2؋e���g�L�J헭}}^�`x%��i[�:p�-x�bi��G�\^ �V���uY,��s��l�i����h\r�_����wMGw������x��B����rUj�_:�ĝ�D�#+^�Lc9?]�˧c�M-hXh?��O�a�߂a}%~S/�D�=P.3o�1Yw��}�B0|&�|���eƎM�ou�F�2��v���7`0=��<`��*�P�\-�:/t́鼐qR�O:)�0{#YP�ly �����E����A��`��C�q|��*t>)��K�� A�{�^�}	�J�%S�v���5�d���n��;z��~ӂ��L�1F���J#Yd���ky@M��]���U�y��������A�}c��2�NY���H_���T�R�����ߓ$�l�u�֭{4JN郡���W��������,����ru5��b�$��k,��W����]�fD�P�%e$��Xgvoɛ�/��o��899��/^ʒ�'��:=�}������F�5bv~���.����G�XE�ĺ~n�`�'���6��f�?������'�Ic�bB��3bL�̽߇�S�0`������0���:.��'@�.��Q�5��
Y�f������eG !t���KG�����G[چs>]nb���9X��Zȟ��Y�������P������z�@��y�9�9���0ǀ�9��Ubrz�<��ֱ�Yz���ut��ܳ��I�Q��7����zĜo��X�kĞ�	 �BǊ��bn�ӵ�?[�-�`�I��\�� �f��=���aC�s��`k�{�z��}; 	�U>�I`2�I����#+6j��A�f�{�8�8f��~�uKYq�G<�����/�������)�I_"��H�c� �(*�~��w߻/��@��.��[}˷t�?$XW���`MF��d�_������{��ߗ��~��>�Z,;��MٔMٔM��S6 Ȧlʦlʦ�E�����߫�3��no�ޭ�rzr��C��O��W_}iYb��t����V��a:@>��4_l@@٢0S�\g�S�#���C<�'S�_��P��~)�ي��Fc&[z����/��hT�:@bѬ`����a���l�A�F�z�G1�׎��l�s���������F�%-X���G�Z�G���!���9�i����=�ي�`�PS|:e���H?����9dt� �fPgԚ���8��;�0d���"@��IW�e��?�L���Zv
�n������}"X�L�d��2�9�<�o��2��D��k�l����uV��Wi2��k1���tKE�	�� �RV���i��|w��.J�C�1A�E	��80Mw-��|8����@0���񛼒k��nP^��x�:F 	�Pf�5������J�A(�g9o��1�_E�&q����v��(i�������i6%/3YB�--$n��n�(3 Q&���"���s 7���A�B10������v~0��. ��n��Mg��gu}�e�\����r�r]���{N�rJ~_K��8�1�s z�g�D�"�/���a���+��;:�&&M����szz��pJ�h_�O���*�i��ʷM-�BL1H�PX��`�g}���̰�֗O-R��`3���*��E!˩����ݻ%[�{��>�P��) ]뢶�[�Y�����J	q�Nơ\�rqn��?�	zC����ŕ$��FW(�܈9�b���* �&E�v� ^u�5[a��&���E^�u��S:��Ȣ8;^���DN�̺%���L&��,�N#�{{[C����Ah����Hxf�S��C�����ϟ[W�ђL�I��I����t⾼���v�\��<����ulـd���)�B�_��^�|���2�{-��#�}gG�Km�_׍�3.�9o���H����u�QVK��m��|泝J�<fX���~�N������C�ѓ�!d��Mm����|��L ��9�f����\��G:�̹�\�&2��b��e)q���N�2�X�!�	�������2G�w�n���u^�L�[J�2�aV��?4i�N�5��?������Wrvv�Ϙ�����k#�Zi��I� 	b6�я������D��z�RV�2�ӟ��s���G*�X>�@~��Gr��}����1���s�M kե�G:����rIt�'A��!X�x���3 �XT�5�O���z}D s�*`�[���M����A�(m-'������w��-8[��T^�|F ���2�X!E��hoG�/�Z�gg�\k�Iz��j7�qf�V�k����}0��G�;�=����X����c  ���^�a~(`���[��j�գ��;$51�D>� P��)eUf��]��`M#�+��1kBK\/"K�H�Z�s��Q�n��4�ɺb=��J��ZӖ�p-�D
z�pߗ;R�G''��Z���) �5�?���#CC�f
��a|���I�K��>z�����t��['aD�[���c�g�|-���o���o�W�T�:����u�����.����Z��O`%Ę{�������ٿ{�����^u��_-4��rp�y�a�}���^b�����< ��'?��:�VD��M ��)��)��. dS6eS6eS��%ˮ3�|g��_��_�;��g 
�W㱼y�B>��o���'� ѕˋ+M�&���A�/���e�;4w�w�=�� �>�������c*��H����Z1ȭ�[Y-
����y���|_��}�ƿo�Ҋ��s�7�}]�ۖ�o��B�Ccm���٪e
�����Ǳ�,D�jw`����t4��կ����/>gVaKu)��q�i��LF�Ax�r�g<��x���eՔ�A���'���3=<�L�<n���B:���.!� �"q&�y{��Sq�0��l�`�'Sd<K��&��Gd�Q"A�[�(��A�_ %(�����ǣ	eR�� �lHdy0�lwM~�*��d,繁0d��5�z}���b&9�K�ȃ�"����oi_�)|���H�?`�tt5bv#|I�ň`��*�U s�2n��5�²,�X�MJod������\��"$p�?� ��XRa$��̘3����ɍ�,[0,ȀA��MV� Z����Σ�j,�����i�V�3g���5H���\�}���2��� BײNN�Uu���~$�dVX��eÚVUb��^�`�FLX�@����x-Sw-�u-5F���}�q?6��!�2j��q<T�K��V�e��������?����r����!gg��6KR}}$[:�r�<������p.��%%D C�tʀD�D�\e�$}ÇkL"KL�>�IaU�_}~x��=,��S�8-��5�iE������Bz���..�}M23�.��z��A�<�r��]����L�9?J��Hd� M8�p6���B��yO��yMT�>/o���Rl/�YY��o�Z��1B����WB@��c0���dSl,����I-u��H}�����d�{������	����X���4��Vr�|�s3��U8���گ�U s��љH �!�����uj�ba^�O����>ׂR=ZGZ������h�c�
��M�24ݖ����D�j��~/�����q�D��clk[D��;�~��w)�Yn�Z��:[���sF��:D��(mW��HE���#��d�2���u�D����#�Z�_I�dIS�%�Xt�������e
������;�ן|"-]�!Q��h#�-�Vl���!�۰� x8�u�R;�k�� #~����g`���q~1[�e0.��������_�5�X_�耎D֦���w�����ޮ|��`C����2�Ls
�T��P�O����[�ϭ�=]�d��=|M�3}9�րvrr�� ����� ��#mˡ� j���,����
L�O������z���ibF��#�յ�a���ӟ����VH�ݔ��faj�����橁��4�D�焁��t�P\ f�rY �&:�'�a�Qh?��  Mɞ�Z��i2��{�w���]NOO��~�o���+9;>�A����Ț���y:�┞7�t�U��v�M���|!��&�L Р~�Ղ�����!���S2���c�����OQ`����X�\-t���^����t�m�\ۦ���{��>;��8hP�?�~,�Bz�,fs�t0g-c:(B��i`�o4# 8�םvS�_�O�l��x��|��?��
n�_:/�޽M�H��Y���8����EǺ�g�8�~$��Y��rv� �h��1�=S��b$W�����S�ï-��g��\��{���� �Bcl�fV�'�Z��j���w>���}�>�t��YZT�7�;\��,��1�����@�Y���Y��~����A9�'���ۅ~�\m�;�MٔMٔM�>� �)��)��)Ѳ��%���7�=>��Cy��>����@3����ӧ��jub�w{dd@.�T8,�zb���n{z��2���J�{��I�^�s^Rj�-�X˟3�7	�ߊ؁ ��G)�	dd�{<L#�	bz��a���w�=x��ň�nhF����gp�_��o���Ȳ�p��qS��T^�:���_˧�~*_|�%�"aڍ�P�` h@ �Ei���{Q�y?P7��)�L�z��ߕv�2:��ӳ �LAd)��Odإ�_HX!�"+@*��U�-ʹAw  d�4,�`6.��2=��p��%e��W�1�`��l5��h2��{6��ڦ�HN_x�V��A�����~@a``�(�3�����ŒmMFNj���R���M�+_�&M2;8�$	<ETDv?�tUa�S0��|�"f&���P:d�,�A�\Fa��BI-��Bp���#���0:�ij鴰!gE��$�Rz�'R�LR+]����>P��������ĩc���T�G_�4U�[�L�:��q�X��3�=Sj	��N�ý��ޑ���]@�f�8Х�?�1��!��X�_g����<���`� �I��9�A	7�3�1�F�g`&z-�hƬ����֏>�+9;=���ceN������_��=�n˭{we�y&�ҧ��$��we��`)�8��6+/p:����y�;��F+��yY���ޞ�X�\\I�W2[d��_�8�ql>��t�sX�`q�ە,�l&�L��'2_��z|M���|����Y���I'n���� ���y��8�c^<%��m�g��ł�Թy���j	�¢�޵L���OO��)1 �na&��������n����E���2U��CL���Q-�vvg;V�]�����=���!���3[������3��&4�F�@��պ��V����nkPW�7|��ޥ����jF����H�/�ub8���ͬÚi�_�o��,I�5J�8���c�s@�>�y�r���}A���I�TV�͠�Lfs��^3[�N�1�����r��=F1w�L�ֈ�d"�^��T�� �D��c��~��X���	�X�ә\�zyv|.����N_�o�Ç��?�۷t�����{\w1~��s9��ӳ�;�H2����½�w�;w��r���X���&��=
��3q�. ���&��ltmă�۲�w��2�E�f��`���������X�˄.�e&K�tc�փ�tm��9�����f�����frԋE��k3H_���-Gȱ��6�0�`=����G � $`���9r_Uzlk��[r��m���%��=�4�^�^/�}�NgHF.KSx֮����m�f&7�`sLf�p"�k.�k7=/Ҝ���;�'��`�>�,\��a�%�A 
��#���%)��4��=�o�`!Ou��5V�Kp�yyD���1`/k����K�qa>fV:YV����L�٤k	��b`�~��r�� ��%%I3H^�14*k�`��f:�ut	�}҇��b��HSy>���u?�N����Ȁ{�1��-� 	�x"��Ϳ����������B殞qO � 9p�*\2�B��7ؿ`.�6��{�}��3h�V�u�ό}'ʺGl�X�Syƨ89F�d�(��/tK��ݒ6�Hw��J6eS6eS6��c��%9�+�k���j_H6��d�4݂ 	����j�<�?<�Z3�q7�;Y$��U��m�gD��{��"�+�52`���G<VU��Ȉo���t� ��/��/��GU�z��!}�z��66zxJ��o��D����	F=r�)In�M� �	E�S���� �lld1�P��ψO��63�K+ �l��J�V��8�u�`2�;v�6�F�̐n�|��R��(�}�N�E�U�������2M��|)��'}"��#����oy��\��h���,j�t�y��	��"�5:b�0�KA�����48::!��j>��|.�5�=m@�Lc@A^���4��|�ճ��6h<P"w�G&9@|
�"<@�������4����f�!׆�յ)ye������C��%M�M§O	�b��׾���H�l�C���"� d&�w��?M]E\f�8��0c4:���H.�������gG��Xl�3��a���t�L; ~!H�z<3�ǚ`%�<����6q��y
� ���1@K��?H�`&q������3(q�E�%3r ~�Y]�Lc0�9���L�*���k�s�F�y}_v�q�hd�x���ɍ�ڙ0�IAQ��(H�����?�����ʳĀʢ1
�,�GI)z����o�i%�������)J�p��g������:�hv5e���},�'�jW�9%A��-; �j$���Eh���!�>Ĥpxߙ��;C�s^�P 
q��*��Z�+	;1�I,�?*%lW2��?9Kot�:,��K_ɶ��n�{��>���z��V�ޙ��������"�V_���&�eimAw� ���I���+x����c�I����g�pY�֎��1T:�`lnL��r.��AJ�?H�6����,b(	<J�#:f;����M2��33`����Bi	�i�Z\���^��w�y�	��T�8OO��>�iC./�����2A�@�Nb���k#��of��B���/Q��@ �si�B�I&��o�_��0����8���ie�SU��(�j�\��M;u�Z� Y$dmC�Ҽ�Zr8��d4q2T>�tr�F��γW�[>�'h��&!�9���j��X�A(����o�S��Ľ�	| ���<p�[:0k�ۦO�IRy|?��-~0�4fг�B}���p�}JY�2������q�Ղ�Aj�.�52�mu���O���t���VW���� ��J��L���@���/��˵���{E���cXG���WH��J�0s���������� �h����5(� ��4���a�$�����L�l@��x�[1�b���0���Ǐ��o���/^0X�����p �h���xt�>��f��z��%�9! �95K��`��Bj�s���%���> �)�a/�`���!�y~όZ�Z K �ZL��^��tq9ӹrI��������8����	�%j0!C�?X�@&�>ܿ�$��]��a�M"�?f�4,V�/d����'H� ���-�Ay/�����'����hGm��� �ج�s�>m�,a��3�~C�k�0�h��x�B>��C�w��o���?�g�=ױ��F�]�de�N��`5�9`��H*�g�{N���W��0y�=��	�����Y:�P<��-}&0'�������@�D������f:}�����O��Kٗ}ٗ}ٗt� ��/��/��/Ƿ������~�Xp |�۰Փ=�"�@�����,��Օ��ϙ�W����Z�$ ��(�p�3���A~�B#HDz<�׼�� ٤%�z��9Z��z��:�lTx2���`L?d�f�'�$�!�;0ߑ��!/�Ci�eD-�6�[��^R&`�g�~.�|��|��;�J!s��� ���(���K�3���"�7�"��84�o	
��� ����K4��y^�� � ђ�D�At�^� �l�8�5������-�䵼��!�\�' cҌ��ȼE��h���Qd#�ߢ�zg�_IgO�͐��f�iL�6��&��Ͳ]����7���%�@'�fk3ǯ��H}��1&y�G�����0�g�0��rn�쩙�w{8ۉ��2o-�^T��%M��WE�d���z��3!w:荿����fw�cQ�7Le�ѰA���T��c5�р)M �}7��g�o�$n(_�2�o(���&��Z��$��-�y>�o�}����M�]]"��dk���_�74�E\��T����!�Sy���9D��1�|�9�r�M<�|6g�}��/�%g����L�.Υ�f2�ڿu����~��H�A�� �<�uczq-��z%T������t��X��'��9{!B[T���U���fa$�����Pdt��ߏ���j��:G�\�S�dP�Whj��� ��y\Tp�j�G!��ck8�4׮h���|��s`X	�6 %<�,#��;ı�$�Pn%���^o0A�u*�uI)���X ���ˋDR}#,>�ӹ�:�@�0��[�(�>��C�0}�7'R2d�ݝNI��;�$���E2�rx<6p��^��@�u3�Vw��j[d�*��L��ϛF@2Bx��H�ჾ^S��(�:�Qܵ�K2>��V˙���<�/d�c��7�h@_�A�w�X?1���/`b1sk ��^E�[��ú�ųq�+|t@$"�L�ߛ��g��R��hz�@.�M  `c�OA���Pn����2Z���u�����,X ��&E0{Hy ��ÚE0G����ڿ���ӯ����RG�j��f�H��3`����D
)1T��$���`.�6�'3�������sy����x�B����X���H�Ӳ��"d�����s`z�{s�Aw�V�&�����`s}�,���vƚ�u<[?�����dK�^`�]�Ll�Z�~��9~�L������D�P���%�՚rR v>��S�T�/9�ȃ�����'4��sBbTh+�d)�R0�j  �U�G&�V�'hHx{�\�����`	ݽ{�@طϞr�.JK����ͻﾫ����o��_џl�H�}4X�1&h��xBM��r��=c�B��VW������Њ^`�<�߯��uF��|�[E1>��P��A�����B�3��Pכj�c���@5�H'�l��^gr`IG`��� �Nl�m	G�.�91�^|:��/_�������?�{���O�r~a}P������ΈL42ö뻍�^�1A��_�o-�{���[���s�h�m��:���
4t�v�o�̬��R^��d?;8:�6$q�C�k(�K�+C6����+{��}ٗ}ٗ�
� ٗ}ٗ}ٗ?hAR�����נ�}t��jF�hfx�b����g2׃\��l0��0�M�#B�Z,Sك�o�4c�{z`�Z���Z��@ �X��n��5����q9�C=������z_f0K�ܟ|��dۂ,�c�7j�#�Cd��TO^��<}�D�?}&_}����:��b&S=tO�=�o%MV��$l2��U��U�#��C���A�
?�t�C>d��q�Y�}�A���C}�aЊ�Q?�%h!�f������m>�i!��_!�rir������]Z�*b�ʧܐ�sZ�n����^�u�n 0�������d��z/����%��w� H��A!�$�l7�)i���ɀ �i��q�ڞ4���ya^��4*��0�H���b椘a�L����c>���m�b0�F�A4`�\j}�\�#pU� ʤ� q�w���efĎ	df��aщ� F��pT��N|(�.�wK��X b����@��%_7%9n�-ͽ�_�*�L#������7�p��p��;���4QU��r�ȧFbrl��������A��]+t,�}��F�Y �."�^2��_6A��6o ��5�ĖL�\�L
L��wSI ��s�W,�O�ś�������62O�5�7��%p�B��^� FAв�A�2�[F�A?���wb�K�7�|<����׶��6vTM��2Cʂ�Rw��}���t��L&�ί�%��$&XJ|?�Ĥ�s���D��y��ҧ���=��ޙk�l!�]&���{'j�$�5��t�"�	�������T��J����A�Q?�M��yp���(��#�^�Q}��l������XBd�}�Urp�&[������K�<x\���e��LS�~�$Ե-��>7+I����ՅdLIsx�@\HW���`up��s��@��D��}�]���#�G����i5������2�H�ܛ�L�%�,@i��r�7-c݌����؀� �K׽���^�.�jcj��g�S.�r,�s9 ��s5}��y�1���(�g@ 6 ��VL�f��x���̿ı	��{��US��(�{=�sR���]=�h�E��ki���l�r=�a���܀�-	�^y��k3]���!׃�b!_}�|��oe9[���k_���Wy�榘lL�� A��6��3c��Z�Z�NA��[�c\�vlK�d"���@d�H6���4OTC*/�wu?$�s�:N�_"c��GY6:�%��,��?���ܾ��kcX'����s����_�  }�����+����t�x(@�X�a���d#Є}�J�ӽ��ê��Uf2���~B_�Go=�}�/>��ϟ��S�l����?x�H޻/��\��o�~7�������}'�C�&���ذ�Z�1�*2�P�����O#�gmx���O��5�r!�/@f�}������k0�������� %�8�:����L'�\Wz�k�$syp����� B�2�֯�c��_g�uO�\��_Q��ӏ?�v�\f�^���K����jl�i�A�@��^�$��	��g ��W��evrr����飇o��w~��l�旀s�z��=���'_Q���wޑv����t^��<$����<U�۬�}ٗ}ٗ}���= �/��/��/��?y(�*L�C�sSw0dp���Oߧ�7���˖\]^HW>�W ; �&�x�p��,S��p�����,ЄdS�x�p8av$��q@1v�0~��G��?����w���.�Q����<���x��{c���Πى�nW��,�����kY�A~8�0�!��"V�g�Y2�W  �� {�<#+��l��;d�ͳ��N�w�&م �鰇���	$Db�&6y�,Qȇ@����3k6�f.P"�8y!�)h<	����6$G��L� Y� p�������~{ȶ�wMoAa��#�D]vxzD����l��$� h�`[\P��ԫ�X��nM����K�9P,�:�G4�ܖf�n��Pcv��Tg9��G�0 �6x?�1�|$ :eE��У�C�?���ڎf��[H�.��9�E����8,I'� y�i�1i��Y�]�܁b�e4S�ñ]��ddp_�dy�3P�"�2"0�u�<��R��L���]a����L	�{¢Ѥ�ٯjf����Nv,xݳ{������e���`�1� D噵�Gy�j�wiM�\� R���Rm洑��:���,]��c�U߃9���>��1��^�Qn��C��E�ku�3ڒ���<�o�P7��`G���k���0����!/ ^�O���*�N2��s�,��22c<�_c-���Jﰯ�����i)��K�Ki��@��9Y)AX�"���7�@���δ|�a�;O�F֪2@c7VŞ�&sDh<I0�ɒ]}H���	2-��ؔ�G� H�#�/
t��k?�~G�XV�l�/��>N�vtN��Ҵc�L��uFc���P����*u��>�����J�G���.�{~\s����63����5�҃V&��.�?$F�3������L�o�=���Ԭm���I�@K&%����L�S���]ϼ�Iǵ���\�jMO K
0����8)b7O4�I�%���f>B2@����&tA�}`�uz]�C���B���@�?����8hwNZ+�y<1������Av֔� hN`Ýls�7$�(�fs��"�����|ޜ˪�I��M����3�kC��Ӿ{L}F��ZG v8���.)��ǎ zm]����\�~���Y������v�y	s=�2Kh��U���7�+��b7�b=2�8�}��]�H#,7�5V%�xdS�&7Df$L�a<���6^C�Reah���F�/t.y��0o�Z&��� S.�r��m��z����}��W\CB�Az���Q�k���8��Ƥ���J�{��H�=��o������?����ɘR��ǀ��"�u���v��;�����X��=~�O�~�:�|h��A�����t��,�Bu�htT���rN�s�&-Ŗ4�R��Ǆ�]^��:Z�����}��l���+|\M��/>��'��O&U��q�;�������N���k�/��g	0|/�Y�w�)�{o��k@������-�JH�o�����W����Y��=������5���N�?���^?z�K9�oȒ=y��ï�^�{�T�{����^��Q�g�u�.�n(lo�:��/��/��.{ d_�e_�e_�(
�'�z���H��I���fhD�p
v����M9��#JD��3"����x �Ʉ��6�W/_�g�}./�{�6�!�vH$��iY��Ϧ����b4�1(;�w~�X���k=4.���AsH\̮(W�>��5���d5h�]p�NMV�P�'��`�|��ad�_0�����r��D^�x��׵�V4�M���`:D<h����v��,�!Sx|p 8��L=��.�mL���A�T�yی��ȶ�w���.x?>�&�@���JE�m�LE��	�CP -\ɷ����8�a��J���z ��5`����<��#���?��4EPϤ�"�5l#�� �j��] �P����Ü&�Q�Y�\_ϵ�yW*A"���u$�-��,S	�HXCz���:�0���� �gm
�ƪ�-�i���@p��uX�. S�-3��:<'�@*g��S:�7`Y���k�pU�pH{!�%[l7���-e`o4�1�@;!U٧� ���r`��6q���?H֒k�>|���,�0��?<��@����G�v���x.�d��0v����NfDv�G�d3�����I���O�귛NA��vl�W;�� ��M�~P#�dl[;sH� �$R�i-5�Z�T�g�������Յ�>�2���g��
�a��#rj)ͨ�:gv@��IR������1��w�:g�`�\�����Q@ Dd-˫\�BY������~�@�s��#-J�蘓�>ۊT  M��!�Kڛ�����7��;?�`Ǆ�����a�c��]2�zu��lQ�W�wؑ�sH!F�=_pL��R�]�u�8��~ ��R$a7���z����B�>ױ;,��[C�^���=�TUK�Й��LZ�Dƅ��������a �����Y!g�]7��։�R�C�:#�W��%(72�y��j�s��X>�ڜ�v�1�]��\g���,�"+��z����d�K���kYK�uRh6"��)���VEe���$�]}�m�RUS������y:q�km����x�[�`.�QN)G?�I�tAb��6�K6n�,v�/R��(�^�K�+%2��A�'v�g���@��an�`�ö�J)���y
Ry�[W��Ɵ��8�yRP ����Jރy���v&<���q�13�}�/bs\�I}��柎�A�N��M�Q�0�*���V7b�ü���$	�ya�O���8V׳���si��k����'����o˲|Bp�XI!� @��D���� o:��X��v����kY�����$�đ��}��A�}�n�&����r�{��rIF��UI`*�<ქ�J��y�0Y�"��xg���>�$�N��D�0���؇��������ΰ� :X����GB������߱e�����9�7J�5�TA�����7�W|�L��^���#����%�b�_�ż��ϩ}�@YtI��>�|��2ݮ���,�������� �h�A��I�y[����\^]r��N��s��{<[������^�^򙐨w$-V�B���
~G���]Mi{	�n�׀����*k�n���`m�rmt��4F�Z����o��֑<|�@nݿ���vc�J.��/��/���/{ d_�e_�e_�(
��n_�z�����b6��p&==���f�{���� �!���˔��#�gd��}���}��������s��k[0��w�P|�5h=�=I�������N7��l"�QO��!
���(�-�"ݡ/�'�|&�����Vʡ���@������͂h�3p6�������|�N$G'����C��>��2����Z�*H:y-����;<��~�9�,�Ɇf�ӫ9�i�I��͋�L�{�c�4LgS}�ɆA �FQ�g(V���@�*4�d�!ػ�- S2���O��.8mZޖM�`Y�����F9&�0S���J0��&��QJ�G@d�Z�f��A�d�� �b���}���B/wA!�]��V"�_U<�ɇ,_��cѾ�\-��0�;�.x0���~��M�D�៍q-�ב��a����@F)_� ���v���`KTۊ�Y�_d��5u�O� ��P	���M1�cd2�l��:�{M������e30��P�I�����/Nۜ���^�DGs���p�sՔ���d��h,���e��18�2C`�=3�- 	�82;��=�\`�٫*"������08.�cCem�#~�����2��\����
��R�b��isq:���5�	َR7�ɪ|�?C毢n��fICGI��%�]�j�?0q�@�vIs���G�.�mII�z����\���d4��k}�`,Ao,Ѧ#�*�vΘ͍y���{7�+�'���A�?�:~c�r�9�] :���EQb����%( =x$��[Yj��m��ޭ6����F��R��ՈJ�6�\B�^x6�y,�ڗ�˵���r��}W���m	  #2�����2�������i��� t��&�^�e�P�&-.e���ֱ�f`ulh�F��!y�h����<<�@�kS�k�M��\��m�u+׏�F�@r��\�#� �'G7Uw�`����S�7}���k��z��'�c}�}K�M�,����+- ��P�"x��A� wDpڣ��v����*L��@bi������A(;/)�wB#9¯���k ���3 oX 7�h����s^1���|R�W�7��p��k�q��y���1�vd�'b�	��t��u��z�J�["�~�-]��W���m��( ���Ib�����hϬ�ai��I%�S*	��l���ؾa�Ԩ#��m�7�n|�*�=�:�ns�WbY.�ryq%˵�����MG���ĸ c������*����9��>� 
�8y/��Qo �������L �:'v�-��Z�k�Xo�G���t��`p#Ձ3���E|���/�6������\��k_?�v'��e�T�/6��F
�f��VT\?�m�NK���_e�X�k��j��ꍺ���װ�E���t�ϹX��hc�B�d���7!X�S�(��{7��s,Y���Zڞ�����Ic&���5I���Z�o�!��:���J"@9]W ���_b����p[~�CM�:��%a}�M���~����G?��[��U��]�kQo�3��=99y-_����Y���τLJ���Tbٗ}ٗ}ٗ�
� ٗ}ٗ}ٗ?h�e���vZ�b����|��g��|>�ΠGl`j����`x�bh���v�7S���L>��'��+���Oe�XH[ߋ����rY���S�?|�C�f3���f�������,U-o��@���{�4� . *8����Ӎ�L�ʴ��9�}$�V$�V��W�X�䛯�I��X%	�I�X���ޖGo?Һx"�g�$��t<(#��7����Q�6$���Cy~E��=}��P�y
�|�,D��R^��S.$+��t���s  O�Y�!�>zX��G�<8��kऴ�Ogx�� ���d�,���T,��]�M"�ٙ��� z�P�h~�Ii�iw[z�k}�܌��0M�d��!�8�#h�~�]��ކZ� (P��������������j���O��7�g.��G����/WK�Q�3 (���"�fw�@�HEU7�X�O)��Q�ۃ$UA�z���8}/�����]4~Y�{O#1���UIx��]I"k�7�0��-��|h��h$��od."S�g�Gȍ8[�hk`Y�����[���+~����q�>��y
Sh^�<6�z\;&c2%��t�σ	��)۹t i�4��?��f����!\Fͧ �N���DŘ+!�Զ^-��[2�|�1*�o��ҁH^R����X
�j;����Z�*5���B%N�6����ܱ)�#c��]��FS0?f����b�(�Nl ��y�����'y�%t��WR����]�������q.��	=V� H��
9X��N+xS|��F}�W�πƀ���˚�hB񜐿!%��� �d+�����_����w$����Zڏ2\�Ԋ�����[�J�:O��u&�gB��@����O�v�<ܗ�׶:��k�u�ѺʥUe���E ?���sv���g��xm�Ϻ�I��R����'rz:�Goݑ���t��Ń1Y�<"��d�Z%�Z�]ڳ�ۀ�`¨�i9g{�(�#ñ�ڐ���o�B���(B@��� ����܂� |�,B{ ��+�m��`�6��gy �.L�sl�x�T��oIo�'�$���נ�q��L�Qﱫ��-S?Y'8~tt<�� �&�R�I8�"|�Y�aE&��9 UWW+ݍ	��w4wx�_nB(ݽ�1����j����-�+ 'Ȳ'���ﾳֱ6�����b����w�ܒ>��������A^0׋��|�B>��S&V��c��ãC��^1���I]���me�/���l�\ ۬d�ҝ@�
w��O�d���+�7� ���JD	�3�6�	�H9@��|����+�7�s���	���S&4ĭ�^!h�T�̓�����Kv'�Z.g�4��vz<�8�t��I �脃u����Q�Y�F�q��� Y3���%��k r2>�1��>{2[�?�\Þ�
����~�	::6C�Gf��lؿ����>&O~'�d��,��?d�+��oG׎v���%y��5�_���e�k{�ka��8`?�[
�� {IY�@�t�9]+]��Ŋ�7X6�3����d�2��@*�C����>�����c�A�b�,S�fJO�F��6F��{����&[���(�����ރG���29:����K�>�ν���|��x��1��/������>_�	(�.a }C�@�e_�e_��_� Ⱦ�˾�˾���R�8@��	�8$/fW����N?:��ËZ3�.��*&/#�����NW,��?�X~��_��|*����ax�13hHy ��Yod����1<F}f���,�u:���fv�'�~[��p���"݈� f��$H�������m=�MCy�⥜]Me:�i$fz[Y�}DO��0��'0����b����79;�3�]�� 6��'�yF�M`��J��.�aV;X�+k2E����>�t�Z̍�[D�2c>���!��x�P�Y�a|O%�.ÏQ@�{�æW2jq�D�w�^Y0*������Zה6��(�Aw���l`[C��C��jd��z(�:cS�����W�9�)�έ ��L�()��@T��9�ĴΙy雇�~'2XS�]� �ݏ���Iϛ�OU9������#K�`=p���=`r�YȪ(� ޤƮ��� �l�(fr�{1p����W������]�~Ā[�C���nnDḭf�%eR,S8pf�%A��x��oq�^��_�!� '���Bm�n0��ز}8}X�������N�ɔ7|�G74�f��o�F���˷Z#xBʭ,;{u�9 +@Zy0� �E�t\�P�r`z�\��W��_�~<&¢1h����0?��6� �z	O�� ���}i�l~�*�>�Ւ�U�b�:j�$h���l��,�
�O\R���ȴ��nt����L�:w�<;�{��8�S��T%2P#}�J�:#C�Au߆:�+�%�������@�|�@�I"g��.%^a��y�6lkJ��,��l���+�g_�}D�?�t�lc�o1�������E��L�_g���uq�j�j���;z\�#mc�iɠ7���9��t�fT�,YLE�.�~���@qxz�K��<(1��Y}(���������с�c�N1��L
�"!)��0�>X#�x	�v c���$�(�qͲ��@�܀c)?��:����Ȩ���a�-N��x�A�P��_�Z�|�D�ܽ/�Q��7��fp��p��� �D�C<�5 s�@�jŹ>�~����B:��Ç����&p��ӯ�^�~oߺ+�����{c�$�uh$�tm��|0����i�S{�x��X�xUY�>��ό���5���x�x�B�����C����� ؀��l�y��Z�n��^��%���p�� ����~6]Ӓk��1M�����L���8id�(Q����ٸ�}ó
�M@����a'BJ��^�@���\YV𾋬tR�-��a)Jum@2��q>]p-� �}X;4 g��[��)��.�`�$*���/uo�q�n�-��|蠑�t����/�ɑ�Id@6���"�t+���`\��G���K��c}֕�f�L?l��e�tþ�Z$��g3�����&t�;h�ʙ5>4��N&nW�K��o��O�EU��[;g����"����M�l��D�G�cҿ���l�H:ꢪ�+ �J�6)3��_1ڏ��R��^��ۣf�!������Z��@����.q�=�a�B�q�^��Ѧ	���oS�oF�T��I�y����|����m�O�_z�ߏ5Ms&����t���{����/��/��,{ d_�e_�e_��
��ρ��3`����B�o�Ј�����p�0��{=]ox�j@����O����Z^�� ���9a��G����P�:�����<����$Y"�4�wni��b��r��7O��n�#�����Me�2�}�Þ��J<�'?��rt0���=�g_��f�ΤIgh�%���4xo3����9�a�!�~�2۰�s澁�Ҙ��p��l\�WZ�1K3�)pA��˹���m�^F�h����u�b�,�S����:}f�!8R����^�+�p���n@Gم"�`QU�A5�ccg�,c�b�m)_Dߔ��l ���Lmٝ8/KxH��Q;b]�����7|.��8W���Ԥ(����m�.�!PP��"�́@"' ��T���VzM�i"��{�zP�,�-3����������]�ֽ�Lwټb�N�Y���7���3�g�A�)�vD	��1L��)0L��A�g�~�|�n��:= :� 4&D$��ѐ#*1i��w�o O#���"���P�r&��������m�n����&��a��Z&s��Yt�Z��m���<��<)��J3c']�!(�@6�e�<ӎ/<��/�w[� �@N�ߟ�	Y ��G4��F����@&�����L6�z+��'3[��� �܆�Q�y�o�jz���x�Ų��v �c �qi����A�<oK��d|r�"�Z����!��n7]��/֕\^��'#z@�V+��ٹ�g"���ܺsO�`��� ��_�SD�;�=����k�_s���y݀�����P F"s��o�}��`���FvJ��9���ח�FǨ��3���|f(WH�Sd�s��U&W��;��Lh..du�Z:���FC�t�i����y8!p�9��'�|�	�e)�V�`t�B��K�����D�_ל�$���`ji��ԡ�o�/�0@��XL0y��D�8Xې"�2Y4XF���L����&�a�|���_�?0���~��l^d�;����թ<��+)���9�c������ݺs±y�u
ߦN�%�'C��Q���� �	0Ї���Z�gW>��Sy��	A�;w�ʝ{�8��˵�#ypߗ;��� �l����j�rp�m��I�Ə*�� <+9�����<��jL�+�'�E��{��l~)/��VV�K�Y�!� ��m-��Zrtt��L�P����q ո^l�{���$!������^ �w�u�g���|P���1pPL��X�`�/��y2\��X��ѵq+&9�=- Y��k��?��"f��AP m�AQư��q�����Y��c�2|ߐ��>�%�X�[3?�<����f7K+ƙ�Y��V��s8Ʃ���T�Uh+�p�%f� ��u�����y��	� h�+�'�W�oz�H/�Љ�իLtY����Gϳ,-��`��;J'{ź�	���J�����Kx �� � �J�#�ވl T����;�1��E#ݦH�m6,:���m�]L(�c�$2
��d��"2���&���4ϳĞ�M���>J�0� ��`�a�ƚ�2�6(�i999�q����O��ҰL,q@X�v�@&G��WZ��F:	���?�=:�$� �۱�����__�4��˾�˾�����}ٗ}ٗ}��* <p��2�l����,�s9>�-�^���!��8��}�E#�#��6a&"FȺ���od�Z�̅o~(>��K�"�� )�F ����p8�Y'� :Zz(̳Z���w.���w2��坷"B�Eeّ"�f��C99>�Go?��[�����޷Y�kC�%��t��3C=��9k�.g�.��x�<�R6B�.��R�Ǡ�т��8�⠸uA]�zZg�fD�
>�7���Ce�Ӝ��MΡ�B�	��m^s�I��i���2�\E�	@~_9YH�!���k0�_m)G�vre�c��N�Y�8/�s�a��&<t�A�٦ ��xVȩ���Q�ݰ�k��;u��p<���!5��Ji��9?;g�#x�4�2k`d�z�M�B��G�:�G����P��ѡG��~�A��{�;LS�]6��3}o�'�7qu���־���`9�D���JJ{��@Q�7C[��07�(��"�p2���@Y���L��KhϊO6Ŏ���(l�����	�3���r�@\[p��"H�8�'$���e��i@� 7��$��/� %��k_j���c~��ߢ_����e����ey���F�[�Yް%C�AJk�̥l�cչɵ���Q�����lҵO_��o��������e`�)�� �6Z�\I����ė���pI������?�`m�d��������]���w0I.��g��ZfK�?:�tub�������m�{p:�$̺/Vr~��j ��G���/9�Nd��������6I$����fzƄ��^c2 p�
w�jƿߣ{��s�V�I�x����4�U�ң�� mȜ�~�:��w_}-W�S}�F?�Z��R@& y��ofz�`(���d���1�nJJ�� �l璯攉���s�b�d�8��a`�(��:S�ɤo��V@�0v�AEK�K	(�jW�չ�c�D��sAV�;��3���
�!o�2@1ꨕ��3�F����6\3Ќ���`�61�еOe�K�w�q�u�lS�&ʐH�� X]l29?���咶�+��9����3��{Xgh��O�n��RO��d��YJs�0j��|Fsj�񅮕�mʠ��gO9/�&����[���c��<֛�}��1y;h3NM�=BMp�s�/��͜�;º�9�<�0��Di:����c��/;d|����o�?�cI)<;�g�D0uu����4K�`��XiX��#��?к��L*��rK�t2��[��Rf����F׀��	r��.A�nӝ_��u�y���$�$B�"2> �B*
�s0�0����`��x�����Q�*j����@�����B"|����5����iŶ�a�=d����>���#�P<�f�5A!_���l)��	>��C��!�	 �΍�w�&�N�����s2�����x)/_~'��'!��;�+�i%�җf~^۾��)��ݴX:/�tm�7;���@���y8眄�lM&�uN3yx�A��69O�����e�&���O�c`��^l����QV-N	:���G�E��b|Ҹj���	�]86�c�h�:�uK>���:�~)?z�]��[��G��uY�!����w�����'x��t�=D���:��\�D m�}ٗ}ٗ}���= �/��/��/t����S� C#�P�����wz|m~5��|*Y��N�E#tj�Wf.�C0�%�s�/�����Ժ�O� �� "px��<�(%�B2��#;�s��g�<{�J�) ����k����
H�0�y� ��Cy��<|t_�f����\N�hg&~��n��ꚮ����9�F��-�D ���2*���|A��L*�����s�r��Fn�>��#�M��.녺�0�D��?���0�@P`8b�<�Y-s�Jg:��<�	N������!�# �n�c!��遴�]���5��&Wۂ����m�,�1�N�M���r X`4,dS#��WHI��<���m���;����G���<2U/..(��v��x�^^�5���Յ���d}�0G,V��Z&?T��Ѓ���3x�kȡ0R@*������l]�F��^�l����U/wR&U� �07S��%e|\D�tͫ��qͬJ YvO�__h]��Q䦁N�zGq+0i^�w!E��kY.�R�2�3���W_�
^`���f`��X�Y��g-�� B0o�] hAߔ�����[�}�@K`�f��/���`t�r'��/�9fKT�I���Եs�.&{U;C[������h��13ߑ]�u�ȡ����T�9f�A��{ ��9)6�te�Ӆ�.r�ח��k�sf��� 6��#��X,\ǀ���A�[@��rT%%Y+D��PV����wd0�Yu�q�n�V�/��f��|SҬrgS��m��x��@ ��N/�"�q���m�ΧZ������o�,2^��	�b��v���hd�<�w�V{@�+�oQ�D�*d���K��(���)NP��B6�R��vK����C��L���VZ�K� !��tn^�d^��B/�m��z	���"�҇ ��M�(�3��n�|r�{�y��_b�<\Z��'�%�V�ery�|,��$�ED���ۀ���Ѡ�#+캯'��ܘ#�����R��*�5�<5`�1�0�y���	\�n�ҹ��V8�d���j[�*ӛ\������km��^��RCAk<#1�F�L�dN囔c�>0���L�*��������rp0���g2�~9�Lt�G~���;�#C]�ȎbHɫ�7IG]Kq�X��+����%յk�d2!e	�q�A@{<9�a�[��sR�܀���k�����HtO��@�✌U�A���۬3ʨ!��L֨�򀁻�ې���r���w����uL߼��d�^q���������j������5�sk���.Ȣ��<1�"��0�;�{����0�G��ܤ�R�.w;}�� �\��^��N���b�XP�f�w�5�y�<���ҙ�ILe��/����d�����"���.|TB�k���mcd`>��|`�#9���U�~"�Ws<D~�D���jI��@}��27/6�#fWWd�xa�lCO�pƄ�f���u(9�g,�y ���������%]�pO02�=�t��k�wb*F���}�Ld&!I�t�sC����)����t�=o�|��[��fb`,IN�1��	������j'��ב8��0��n�.��o��坷ߕ��ŋ��t}���w��3hs_J�$F�$V�̏v��=u�݈nG��:���󮾥��������?���R�e_�e_��[� Ⱦ�˾�˾�Q�����r<m[�1�
����e\�8�ʋ�B<=���2���!���@��4��>�\��Op��0(i��t� �n#0I�K����j%�ř\̻rt<�����ܹs_�}Y/����v�I�K#k�9e�|N�@0"�b����̆C�[��|����s�����z
��8f�(����'[ȏ�@2H-=�e����X#*絬��e=��ԯ-P;�~��C�����g�9��X �Y`2dN ������@��3�j�}]^g�5dN6�53�M饢'��7-pj�Ә6��%J}���i}HГ��;X��ԝ;��wߕ�=�4
�T� =n ��r��Z���o��O?���~KV��t+���q�ȵ�K�Y��Cf4#�e��M������{�,���%dR��Гw�eC&t�e [�fDf)�A֖䋝E�3����f���s�X<a�Ą^�����B��Q����Ec���^���4+T��D0��`��m3��-��f����^em<�7����U������8��^��m�j�!р���zF ��/�!�ڳ�;0�v��e��?Ǒ�3Ф�����ƆB��X�:�r��1�׆4�3X�s7�,����^��R Ƕ��4�j��7��CɌ~zx�&�De���;��A��Dr�j.�� �HA���E�'��J�:'��1�����
t�<�q`��1i)W/����9�{�m�T�Jk|(Q��^���H�.tBL�b�t�#�cz�S�8�,hk3���w2��od�@"��q�@��$�jd���y`3fPn�,��IUY%�qL�L�s���IJ%6�����{F� b�ڽer r|�#���u�k�z��Եe!��X�3��[�|gf>Eq`mW�3r��0���j:��3 <к�FW7퇩�Z�io�k!�ƀ]
-��Y0=l�2�f3 ��b�1�o���ns�,u}�C��u����PB��j�s&�g�|GO��4�|g�i��f�k]LY1J
L�c��ԁ�y�|��iU�>�|�Y�����:w;r��5�5'l��+`�F���?{_��_����ޏ	�c�>��ފ��o�%�|���x�\ǣIh��9}Ƶ `í�'2����\^_\r{��!��T��_z��mJvb��w�AtN\�w��z��@
0�P�mh���t�3C�Cw�d�}p��-���<|�H���w�6װ��K�I����a���˯e6��O��:_�`%:�ⴎ�>Y�������u�=h��1}��o�?�NRS����]s=��z��׎�U�	���� �6�6�$�,n�s����Y�� ܎�\B� @�ܣ�W"��z��1�fHǝ�I3@���Ƴy�6sϭ�q�^�:��t���gEȂE_=����eV�%A5�E~ʮ�C�2p��PX��;V�?��>S��o�5+�|�g�{ڥ����n��v�"F�t��"�J'�ş��P`=E
�T%�{�;f�/H�	Ț1veaTV���֟����#&M�?�x�\���~w�=�ݻw�v�lΣ^�] �"ƠO�z��<e���i���FgOo��gP�eK�e_�e_��]� Ⱦ�˾�˾�Q���k�t�p�Aٓ8̤����̦�r;pA>��dE�l  <�%[�
J �4bd2}E�jfh"��&�rXYjq�:��Q�L����lUH��Hԍ���O~�'z �H��u���wF	 ��z�����R�;<�eYEc�WS'9-%�鵺�B!pل~��?��9��N��
�o�<1��݊�p���+��l�d(l�R=0��E^�!ץY�@�̼�G�*d�g��H�Q��j�����5�����^�c� ��L}��·��-���c��{���f2^��5>Ɣ�����q����<z��<xp_nߺ'��Cyp�"hg�'�~��3ф�e���������`'� p �޽{2>:�G�Q�d�M��B��)* �"���̾���(հy`�9�� ƴup�{ �A��ə9��F��4L���H�B۵}�����ȝlGT�M��I� X!�$4VT��9�_!u ra ? �QT�a�>��hkǝ�A��,]2�D�`��P� h Ћ �M���5�� b̗> Zϣ~_z��eh��4�n�B� -�f�54�!�����]0��kr�	L�)=u+�	u�{�R2m�L2�5��t;��|���q�� J�Y�4�}�������o���O�3�!e���q�O�GZm���,����7uU2�U2��Sy-pL�q-�#��Z7��}�s� ��>�K�G�M�%�%r�e�]�~g@9%�_�s�c�% ����wE&�����F �Z�v�J��+�x�FZ�!�nn|A*7F��-��P#��?N��p"�3B�LI�$-C>(�����k��E���11%�О�ו�=�kB�mK��v�r>z?0y��	���E����ȝ��2��2S��JR�]ZC���'�r.kYHOo~4B(�L�����1?i� =&G�g�@��E��B�Lt"��:�w��mS��� K���s�3�r2Y0�6� V��5�]S|7\��GC4�G�$�j��~-~ˍ-�K�\�*ʮ�Rҫ��N�0a4�g������1e��R⿃�`��ȥlҀ�Pf�l�B*�$������$$C�3XO<|(���o��+?��� C�������9﯇9J��|>��b./_���?�P�|�%?�� OR9h�>��~WVە\^]�.������C���c�/���w���x<"�������w���~�\�_H��mӍ�8�����m�|�9�����rt|"���/�g?�͟o߽C9��y9`��`� ����+?z�9��	�9;}%Ͼ��Ң�˩�r�@�ў�>�Hw��ҼxM���+�]�c2R*��jI�5�d��-����V F]����&K�n�6�`@��Mה���Vޖ�a3Ѯ"'ل��߀��u$�C��ܙ!�2Hd��lt���z�wvt_����]��,��w``��_���]B�1_�:U��[W�s���g(���%��5Y��~yݶ�'�y�����C���&��u���\����ef�\ ­��|m T��e%][ն'�ɼY��MJ 	��իW�������g�w�����ʰוh4�Z�տCz}j�{5c� d쑥�������!]ؠ��v�,��`�˾�˾��� ٗ}ٗ}ٗ?h��&���+����c$Ԕ ��7R"=h-��2b�лF6���q��g)hPP[Uߟf���>�Cj�B�^���5�4X�rL��
��aG֛5�Y����A~8؃����l�z��j�]-��r.�J�k�H�9yf=|���s�7�|-���Ƀ�������\���}�b�3�Ok�+. �<eiF^lKI���NY-W��� ���)q��S2"��-CȂm��9�e���-��N!�3��1�pr@0	A��fc��G�l�mb�W�FJ�!�����h-����ϨM�4s� ˖���^G�^0;`TZ�����D?����+���/��ޓ[��P�
A ;#`�W���j18���t�y�42I�%`� �r��`$�c}��H��}J� x��������'rqye}ً�w'	���pM�v^$d89"0t(�R�V�X3�$�Bg
{���`��
�c@J@5�Kq�pHFZ5���@O���GE�+�
 QJ��m��]bF�1�uq>��j���(��r�d��=`Xp,���mײ�2��"L �L�S��]�<�h�� %F���-kS�k�$��e�S3zP��G`��xnf$��!�V��F��Ȳta�� |Q��Bf�f�����3�S��~Cz�3�����u28���Hn��`8���uK���Z�)pX4mh���_�@ @DS��P�� z�OB?s8�:҆!=��s�YǮ�%����@�I�|.Ip!A���	�<�9/�� �����0�㓞�&�:�P�&��?� ������7%�Ĥ�j�:�c��,�N�	π@�M�W5�<�xJ�Ѓ$"0F���7�j�XI�Rd���pM̝c83K �|E��өt������ 8�P���P�谣�P�Yҫ4�$�m
��{zMo|�}�+)�ڮm�|�Ur��,�P�T y��1��@Zn<$���������[Z��DE�}*ӵ��qG�J ��>��aE`�Ӌ��>X|����N;�$�� q�+� �-X����h��&:������.�_L*�+�^�pg���' �WA��;�y;�=2���Њ}3���6��J�e� t��y�E6'��!�V9;?�M���ѭC��?���˿��"0?�����Ou�~.���Ċ���Ϟ=%�b�����B��S٦k��"�|��:)2[o��3���n�u*/�/��?d���_Ur���3�k��_%_�>���o��Cf�΍>�RRi� A��R�}�@��HB@��/���	��Z�v��L�j7?�_����s?��::��{���A	�ǋק�����~"��9e�hP�sT�6/��]6�o(!N�f���v�$ ��[2��1w��b����ѹ��@{-�|pO�2�4�M��t]��f�N`�7V&���I)�����6�vIu��2��h{���f�$���N��s^o�!���`�Bj�+�����m��C�ӗ��O��h2�u8��'"����o�����"����5�'i���	�ׂd�ۺyM��e����.��i^�`��M�ύ���gɜ(zY^KZ�7�����&��/!��{a�9$t���I�:�x�V��kt��Y�5��7`3M��/��/�|A��>��W#��o�q� ��LX���\M�:�zdQE��4����o����]�����Z�'� ��q�}ٗ}ٗx�O���/��/��/==Tn�3IJH-)3׃�����ɽJ���qʄ��022�����{��N�P"dB�H����g2������KI���yL9I}�����M�l�$?,�]1ӑI���z������$��Жu�2��v/6٪N ��>O,�N����3=�%����*,����rtrK�-���sY/7r�ͥ��mQ�%�д�&09�����<d���I;�56���zN�k艛~v�̒�^C��e9� `
�3�4���j��IH�y����c009(>�S���j=��&O�A �%fƉ�1�ӳ2��u�m�`3�x��%2�g�;��������c���K������}ׄ�J�5�-�%��9�B $�z�{ �T���2A'�78��^�~P�Eᛱ����ё����_����W���s��%=f���� �� �� 4��<�P��)e���-+4���ee�A&#�[&QC��@'wp_���'
��V)��͓�V`!x���#����[�Mmzh�[�p-�Ŕ�����΢���i{�`���WA�=�A��Z� w��9���(o�z����*��<0�K+lSW�����z �i���k��?e�{��u�X�l��&��$і�����<hK	�=�"pL���r�����%�c�:.  .]D���l��II`� GZ���l�0��:�7r9[�4Z�C�"�:���I�պ��<zK����R�%}�o��@?x&d����@�� �3Yr~�{bii�~B�'��ҰW�K�n<�J�S��}y#r0�όc��5L��} �F! � i��gr���;3�+�.�it��h�]��09����	�lB �C�P�h�ֺs�`��P�M�$ U���%H>��o��Tv�A��MB)7f:����Hv��D��a n2^�N!�㖶E����b�sm G:���C{�h��o�>���rrO/N��K��;P��:���#� ���<��Y)w�r<y$Ug�u�'R��[��^�\~�sl$��ʴ���W	ׯ� ���$���g��6$��T�7� ۥwv�k��sB�� ��k����@?l��v;��xZ����()�F	cYi�`��Ja]k'�y�4��C�#X��������͒e�uؾ6�{�������� H~PP�_�5�TH!� aƴ类.��K��^k����1��3��ӑ]U�e޼����^kQ:N_��#��-�6̝k9]��`��؋�#1��Ln�#� ],S;�P����a��#��|���I؍�^�g �������RF��;'#d��uy���ɿ����ܹ�`%���3��g���~�K���~�3��r�H  ��IDAT�p�(%XQ���e�	q�e�jE��y u�AX"5�^�B�|4�v}N� f�U��O������ޒ���P�5'��l��� �\�vC���{d���ۑ�^�$.���Y�D�u����yQ���1�������IJ��{pE��˃wߒ���Hog[�=}LO��bBIQ�?�����L�)d;�z9�-#��4jNڬc�(�����2��o���j>�m����΍=�/�K�ݡ��x�I?�j��2��V�տ�>9O�ї���|�ݳ�M�i>'���϶u�t D�<?����Wk֤HCJ��tM�օ�u>�K���.�^�<�W�'2�}M�7�=@�{�4�"��$H 9�8�:ֽ<T��Ś�5V���� T���Qu���l�uЇ�/ȱPK3B'��ʯ����J���������x���0_�,{�g�s���1!Ԝ,�H ���>��B��?�^"y���3���?!舽���1���s�����ov��d:���:=9��������ǿ��wzr����b;�z ��K��lʦlʦ|C� ٔMٔMٔ߉R��G�3�'�V[�W����6M�_�23kI��.Q#ܯ;�H����IXo� {[�o=���?~,����r�ꘁCH�̃� I�l����@��Yy��e"��}Q�8|&����QzH��>1�}����=09x��e�����,�k=��Ȁ�u!wuq)5@-�$��b�����nG�w��XΗ�hB��n�� ��|&�<x��o�}:�zY-fB��2Pf`G� <p@�O��!�N��٠�g�Ӑ��04e0(/i�Yx�M��2� IA9-�ڹ�ff�3�ޓ%�Wf="{�5pF� �� ��;\-�g��ڔ���d} +��w�f�lԨQ�Y�����Q?��;zu��J������Jd6]��k����;���
$�ڭ��>���P��N��?�Ih�<I �!��X��I>}',�>Y�$�M��ѿ|�(!��>#���΁��`���##9eV����#�K�v��LǄ�����"}�wn��C�[n\�.O�>��ϟ��qD}�C����S���@�#�����l�T�B#ؼ, 8؄�d?# ���� ��o֛�P�������' mY����$.RJ��Z��O���I��m.�!{���
c���3��'r.��z�Qx	8U��/~d�$��g�F�󂥎��}�M� 	5�J�K?d��{�#����w�����rr�չ�dUB�|E�7����9�1�#_���h��_8O��t�{�I!��c����t/R�-Z�U�u^Ѻ�>!���wt�����ޞШ׫7s7��������b��h�t��ֺ�r�C�������`,e&y��S��}���{-�Vy��,�I}�y���$�ں��\�gl���{����0��R��|.�^�|�`�d-G���_?����t��~��� f��Q���`H�#�+���"@�<�u���k7��;�nT�z����R�&�y<���$A̽�k�5��t�k��LN��k��õ�����֥9Лi�U��0YI��ֈ�_%�P�`@b*����4��"��/���A샨{���o0*�����O�j����?�Z��qA�"�4(�V�Gg�Y��iY1�J�gc��6>KY�F����@JyEl�ޠ��(V��]�zrzr*���A�#w����lS�2]��:����<}��|��C��:����~C9%�Lbi�sZ�&�f0�ߏ�}��'1���"cI�Y��Y&�J.�N	$�L[&���<����]o<�>5�U�2���C����G4l����B��\���1(l}Z���lC{i]�Zm��S��`-F���jR�r������<y��<~�P}�P��	�FI�\�y��I%�����V1�Hr�G���"�
�:Xz��H��&��������r9��},gǇ����u�`�
�b p�@��沽�M�a�X�+��f����t�5�۳�\}�Q�iե[kr^_L��ú������/�O���Ԩ�dV�vp�=ڽ���.�W�I�.�S<s���\�5H ���ϔ�)�P�X����G+� 3�����o?*I��������+��N������}
�9�:(s���O�������c��-9Z�*X����v�`��lpzz�6���ϿнّΟ��L ���
�n:�'����]�?��������z�_n �MٔMٔox�  ��)��)��;Wpx�y붼��;�w����S=cz��(�'���F_���2�=;h�qlF��9e�b=�޽�@~�ӟP�b��m9>;���c�S ��KP�`@�L��L��d=|JA ��픲3��AŮ��awux,�AVK@�|� �d�H���{��`�<�=����00N�G���-�~*Gz���gZ���.�!Cm 5�$̦��r�FгVc 4-���N����p�o0P�Ϙ�F����3<�yF��<��ӔY�`M��!&K "�%H��a���R+$wA��������M�?��e&����ny�# �Z�R#C�����+��{?��9 �0��tI�,Z���j-G/_ɣ/ʳ�O��&��_�c��1��.v���9�:��ߗ�k�{�� ����f�^�q�"��|,|ks���I;� |���[ìb %�V���`��{�Ze9eT*����ؖ�_����d� ��S8�A�� 	cޜ�E����nKw0�q�'�~�=���ȃ��hV���W|=y�DF�e��� H� �Afl�4/
�,��'��ez4��������K�Ч`t?�N	P��P�J��ϖز��3�M.���8���b���0��	+����fގ�7�D*ߑ�y��D�`p��1����}�0�W�&T`#�n]��5�< sFP��b'��,w����v�8ju�r��M�я~�����m��^ 6����kU�2�޽��e=׼�c?�}fL1	)��LKNY%�je��2/���D:�i��G��@�`?��-���R����{],�)��m�@j���#��+����t�����fC�rc���ʿ4>�����Ƃ2�.�3�� ��C-p�3��4���uKg`��ri�S��֋D��@�ѥ����x!��3�=�1�ah���5G�D��?h�s��D-H�9����Orr���Ș:�s�'�HsԔ�eOZ ���y�:�/rN���"[nC�j_D���d��m)G�z���S&C��W/��tN�K��}��;����G+ ;d����^��mT� �K��ޔM{Sv��+/�U4� .查� L�N��Y�!JH��r]fj��im��%��K~Σ\A�؁��A���H	����阁w���ù��Ϥ�����tt�������_������Y��s�s/��^�|)��������Ϥ �XI����O��h�9?qgHr0��j��t'%\c  
Xy FJ���_�#����j��d{'�ugNٹv�/W�� +�ƍ[�����))%��ܗ2[~P����2	'�s���:�+�w�^��3�Iyz�D�:��=��ζܹuMn߼!;;;�
�<{(�d�d	��&WhR�y>��nL�w��M��T�S ܂$
 ~�Ѽ�� $9*����k������%@��~����g��$�a<�� 5Hjr��ra]���f�S�:suL�A���+Nu�ϖS�[;��>G�'@��5�2�/��de}kυ�C�ز`��:�/Y��d���7;�DH�A���̺������_���WR��o]*i¥3I �뚌��/���f�p�p"`�΄5&+�� 9{#�ݡ�p�[!eh��@���PZ_5d4��?�?�C]O��V-2��J��S����dS6eS6eS�Qe�lʦlʦl��TA(������ߕ�o=`���O`ڋ�=t�hH	S�n�+�VS�h68^���	���~K��{��6��N��x�hփ��CWA�"�]K3�\,������^��H��tӫ)�7\�(��{ z��h�4�\�)?�����;̮}���$���]��|6�.�O�,I0S��oD�Sd�'<`�Έ�$+JsP��>d+��t{� hQ�y�%�R��Ӄ�zIF	J�U��J�f6b��� C��cf3��ٚ�Tfͺ�����LJPn��k�5���\Qv�
�X3f�B�e[vww���j�]��6���%�DP} (���8<d��xx.���?��5]��.�G�c�nݹMi-H!`	*��P��Ne83c��������z��e )���x�a�>��9�fb3A��X�{�<* 2��9��܂O�9��L;ԢX�_e�� @a�ɕ���� ����|��?����w�m��W_�����_�B�=�uc>�g�%A�JR��c矂la�,^Zp\\��b&�Ef|0���A���|�3X�l�,;[?S�꒹���/칲���t���98�}�.��ߙ+�bA]�~#�d�������2��ߏ�}�`o���"���η��IŌ^1\�|�5zP��2G ��O�ݗ��yG���~ ��%U�NOezji��Kha������Tf��e¼�f.]�6���|���Bq-h�He��8Kd4�G:�L�iJp���,�4��4�:_�mJBy��[�؅�RN��r��
,��~ �ޭ&�<}&�t,�V�U6g�0vL��S�q��� �Q� �39�<3'�D��(fߣ�t� �m�hL�6)�P�>�y���.`8��t��-�"�T�V����)�S�0^��y�D��@�:�x�mBe!y8.�;�_����ܸw]�nlSJ��lRF��/s����R��_&��b�_� 7�@���1=�:�A�̊(j��;�u[5��I�`Y�����X��=�#��G� �:]IT���xC�?I��9.I��J�z��Fn��K8��,�����Yx�n�ü:ɩ�I���IK�e�ucXA�)Ie�_Hڊd{[v�tM����M�K�kd����+/�����|���rz|B��d�)�sA�]���qh ����V:e}�(�S�]�y�LHQ9|�@J^���H[zn.����sr~*��>A�v�E��������KK��j^�}�9����D/��s̿��C�w��=�����@����;�{:�gȘ�aX:ͺz}}��02Rm�W�0#2(QXg؟,s燝��W��)�Y&�0�bn�o	$��ߖ�\�O��;[ܷ� �������+�/_��䣏>bP��}��9ء�W�W��#ѵ>b9�[5���c_���p4� "�	ώ�Wֺ�Ou@]\���i��1���l�-}�f��ӫ���ra>+ģ\hA�����o�f��a�N���&�<w{F}H1b�� H�N�(ʯIF����_���˯����?{�L$�����Ty	Σ,��@�5�lO�D�dD���=�2L≮�{☉H�@]{�g�G �ct$����0&�,�9�2��}뛺�]�����ѧ�����7&Amʦlʦl�7�l �MٔMٔM����=������V�q�\�~�2k�����m`�+�~����`-�8G��,v  ��mfD�0�?{����v@&?�b��0��-����v�����P��o'���)�f���de���/9$� �Ĳ�ߑ~{̸<88��wn��ޞ/&�2XU9:<c�.t+6�S8O#w@D	��(��L�,�� QS��ڒgk�)9�u�x>�C.��3T �)�Tc�*u�TZS|�Z'AYƞ�k����PW�|���<�h&LߏlM�@�]g{@!u�8���=Sx����� ݼy��vzr&9�+�!m�@����2Ȕ�����C�z�*Z_}���+��܅ˀ+� D����={F���;w����'�L�ZK^�x&�~��<y����u¾��)��uF�&�_`J�����NSg�*�D�٥���e��ja��Ҕ4��?�y�\$hPo��c>����}�[�j7����_�_|.�٘��YD%����Pe\^%��O߽0$��21v�~�K���,��Jp�b'�]�/�^G��h��V�'���Y��������x�������yh��p���<Xiᚎ���� �l�d�Կc.I\ ��[������9�u�'�)�+(=�	�S����
�� .�>nܺ%��-y�������~�399�RZ�B����(�?ʛ�e����d�.e�.�Q ,���%�L/r�8�{!����t2$��{�����ť��	!�K�Q�E"���,��\���n��[��J:z��7�>�mSύ��:OQ��U���A0������>�ÔF( �:���,G���P �$y��Gd����W��k�|�5d9Z��jH��f�'���x����+� �tʊ�@o�':O?9�iuuӹ�L�29պ͎�;�.O��o�Z��bz!mF�w�:����c�X�:rz�|����g�gVS!8�^=��������� �D��l҇�/1be�(OD?���~ͺ��z��9��Fa����L��<e�d���~hoȸ�fZ��I��}"G6�3>'C	�A�p�5� ����=�}K7 1�J����8���]� #��@5����4 �T�3��(� �?�mx��8`��%�>5�($��t�r�>��SM�P i��'����f�N��! g&ޜ����5A^�0|���	:�d`��y�;~ �-��c�&�n�D�K]w�<~$_}�%׺��OF����,��	d��͋X��^�J#x��[�i�bJJ�αfzڠ-���޺+���|�����g����.��ڡ�s�lS���7��� ��u�@��w�cru�@�g��os�g�P�[�0b�ׇ���tb�#�o����#y�<!���o�u����,R����L>���<�oB����d�����c}�{&�H�+0d ���|	���c�>��u?g�v��=����9�D[ͺ��:�՞^k��}�v횱������;$�0F���RWL<���k�I�N�,^�����߲��$����~���;��������Wا�3�s�#�27 �>�pH��0��'K��x��i
�8��,����F�W��==��XW�'K@�2�᳨k .`ݸz]6eS6eS6�]6 Ȧlʦlʦ��K���C��Ǥk�nI�;��EY�S����	��3ȴC0�� 8���z��K���5��,��˘.sA�`��\�f��3�\�L�K3���z�)"�|�e��=�5�U��{�Y�Hh��;� �����s����ag��,�������`��ȡe�k�A���:���w�X$R�#�Sg�^(� `��`/R0���4�'^8�F1��`ɚ�%Lp0��6� ��S�*4�ܙtgf����e{3����1�@�m��F��dO" ����{_�Ϳ�7r��5JZ�_����/~�3f�6��p-�!�� | ��f���V#�i?
$b_	������28{C.���a@���8�����<~�X����Y���@����\���p8���(�#HF?H.`�U��#�$��b�qh���e�1ώ*�]�m�!`�3Fp��9����1j�����e��y�dɠ�?��ah���399}E����g��kq�`f�7�b'A�/�Q�oNPǘ:���	:�l�� �� �g�&uJ�P�&���~.������{8�F��5�s���U0�E���(��
*�憈I�-�B�Q�2�S�~PE*���67��� ��PJ1��y���1�B˝NBc�������l:��R>�@�\�"?������G������=�����s9>���e�����׶`O�wQ��ݯt�ykA�&t	�x��������Td|:��C�G��ͯ������\�殴l��z���d����D�܌,'ȓ�е�~3y�8���փK`�:����RL��	��
̩���Ac�+�J�*���[8�@��/����*ܳ��$$ڳ+�s�a0M4+�~��)� w#4O�-H���1�����+�3��ob�b�)�0H	Ϗ�4�1����(�z���?��9�vWGU��N#�:�{���*��=+���`��q����wF���8Ѷ�Ou�����ϥ�7(�AN�NY_f�[��-����'�?�k�8c���y�[+���'>����ђ�{�H3����Uc2e�t�vt�o�:�s�ڝљ�ۅ�.������o����9����D��1�NNNd<��\}A�z���V��`K��C�_��fM �����P
mc���Em`�^�e����@*���7�+3F�^k�Y��k���`����� �`u�ҵ��;�����|�/�U�+5c��O�\�M����S��їr��	�\�#`kb�#�OQ�g�ߑ�}ӗ?���~���W�ݠ���&��`L�u�����j���H��xiI��0I��akְV�5 �d<���S�}����\:�ç���'r~r&�Ǭ�g�vq�2� �@�,X�PoX?
ǂ��zo�% qH�z���^	P
{�����o����y��Z׋���\�����&���Q�6h�]��1K2z�-fs9>=��_�M\rm	��{�ޒ���ɝ����H[����pX˦��e����*֜��<�*���<� �=�������L�.G�@^@��z/H��4e2B&&oe� c��wX����^��u �Af�2�H`�X�	m<Ӷǵ�QVPV�`"�:/���z��J6eS6eS6�_6 Ȧlʦlʦ�Δv�C���]m��P�аgN����|a�G�N��x\�K3������C�K=@/�3ɐ����:��@���� ��I��<I �� �,oH[%��a�3�t�7���挫��j�O�i�@���2[..%;������:$'V��^
�~� 2ܐ��{B+ �Ug!5�q�o�jq��'��^/�Tu�}3w%>��$�銺@�"|2��/	��F�k:�n#���w�>�����x���j�h4&�s��̤�ؔ��p�%������?�}y���0��ۃ��Gr~6�F˘9����%5�RD��2���@F�~G-�9O���(�� x���U�j5ӟ/%�V4х�8�,`E1���O����s 紿�]�s�kf�" E0�yCx53[�9rd�?y�f� x������br�f���ӫ������@�'!Y5�fi4j�+�!`9y�s!����5&E���,%��;n�jߨ9 �XCkg|�IY��sBBj��Sd��`�uĬh�?ߘ�^O����@_D��rNPRoZv;��9Fc���)���g��`��(���s���ƧG�Rj�m�߯�7�$1�J2���P#��e3d6�*�c>A���X�����lf�����W���}O~�?�������O>#���Ç2�����-��҈�����e�[�38[�\U�;	�7:FQ��\z2Pz����k��j�]�2� ��`��n���y�>��LG�5�G2Y>�����:ϢuL�������e;�@.�G��K�<�w��Z���o�����| TT O�dr��(�����>30���6���� @�G��e�We�0�U�:��R��N�'2��o��w��c.����!�+:���Y3V�ؼ�e`8�5����D�.�܎��K�=�^�sI�~t
��5�$8_ק�b�/�P7?2l���NK��arY���\@��z�i�� C26��l&+d��Ml��A����%���E)�l�@\A�� �S�_0��E�]�zK*�_#�%0��x / H�E���ͧ�XW����z�5���TM��'#ML�.���6���Hk#7�{}�e2��U7i�6��`E_L�����>��?�s��<��_����s  >�A瑩3g_�ma�<��P@\���Q �P�ߖ���1-�O�t|�7F�{���al��D[�����D>����������g��v�E�w��b���)��[�.��ج:oOt�q��<��+�r��{�]��ߗ��}�J@��@��-l��־/��z"��T�_�j:�ܗ @���q�E��vd E`�`��,^  �/��㇏d:��\?�. $�خ�F@������t�����i� >Ӻ�����L��뚭?�����̋��#�۬���׵�d�%?��6��Z�L�@�@<A� v- 7 F�}����o��d�޿_��^���g�`��J�!��T���@72S�(����09��W�y~g
�SE���?�}��	��Q�5�>:f��1ϰ��8à)3K�(�ˣ��aƄ�3�IHj�c��8�������zm��&����?�Oľ?���r����R�bz�4���뭞��c}o!�.��)��)���. dS6eS6eS~'
\zz��xu(W��ԳY��d2���+j-�ef�8�����`�ի#=�?������ݪ끬E=���3V`�X���������L��$-��8��2����$,gv@o9)��2��HPz8{%v>������P��dp~{�/�����d(�Ŕ&���2��&�u1�Q^��.Fr���h8dF 0/�����H	���`�@�ZT�dI�$HW!�S,e&h�m��*�դ�L*���4�a6�$����YÔ���pM����Y��<*��JDg�C�+�n��B���fE�ޏ,|���W����8A�~<��r� 
��qP�DM^X  ��
�����Ч<J�Z�sN�l�@Vo���^����i�#c4�[�-e�
˼0�Yŝ^�,d����;�20u|t"�})��ʌ8#��. �D��Ud �a�>�C{�2B/M�!qS2����;1�3 ]����6���K��4c��|nP���$$��!ea��	�%`�݈��eVlS��"��m�X�7��1h�ZX@u�lO���3P�"B`1�D�I���*B��5�ӑ�����l���g�c��ἁ�6����ֲ��2{��Y��I��#}��~������_V4E�3�%Kə�bܒq��><>����MPC)ޔ-���Ctw����}G�>��Lc�0f>>>������:7���Z�J�G`~A��L�H?�
��W�T�93�� H^!���"s@�yd��2-S^�FA����5�깔�LZ�@v����H���9v"C�;�E���`{H�B�r��«C�+��#��,`i1�߷H1@}3Rf{�H��/}V<�� J|� �o2���}�t��+L�h�(p �U �N)���:<�[G(�E�Pz]}o���c�[��Qj��Z��Fe"�^.�W2kԃ�O��`$��v�"�f�soB��R[�ۘ�9� �K蚗-������R�~�vƔ��z���t��d�2��Q��b^���`���w^ ����g��vx�Q��\��\6��/d�����1YHk����K�3�!�Y���	7�f�ܞv� 69: ��4� e�����n����w)��y����:�\���ø�TQ�����Z�6�7��<?XzXg0�! �>�������ԝn�l�v~�2��	�p��|��	y�f�KO��R��
!	 ,$ �A���7���|[�z��/��/����OlnX�d[�u�|���ժ��U�哏?���˿��~�s�ۥ\�rM�t��n5Lc�\�R����'Y��n��@�J�+1�CNp>��؏_<�R�ݼ%<��o�5�l����W�^�?�������g&?����D�7q��&;�U�<�]�<���u���D�}����ń��ؗ����*1G\Ҧ`���!Y�|���	��@�W~c���cmoo�; ?��j�����d����u&b ) w$?�����26��Ru�mɰ�)�/��osm�F�~E��;��ѽ�Y\Ol{�Ct�K��s�1"��?"(X���Ϋ�V�<�pR� �r�s���~�|a�{]�<����ʴ��d^S�43�P)�z�fL@A2��w�oM�R�5��#�>�NA2����>�߰=��4��"�6�^"tl@ 452��ä3�_k�h�U��)��)��)��@6eS6eS6�ZZ����I沚N���!��w���ެ1�z	��$�P�8���:)�ϰ��À⧟|./_����ܺ)����딜������+f�O�nvx-h����`<��z�F�/�1[�l��I�Ֆ��_���)�+��gO_0.q�T!k�����_����Tv��h�}p���ϟ?��>c\(y8� h8V�i���gQR��lE0t�����[-)uf�ès�\3�N�k�2���V�̓��}�J�P����Z�w�O@�;1}u�
Z�����#P5�Ϙ	IɈ� �	Z8�6���fsY/Wj ��'�#�8@�(�;�4���~���PJ#��h
?׶AT����)��荢޾�;�1��9�&�Ǳy�t���\������,�}�=ڐ^��}�+_=�J^�xjZ�q�$C �wC7 ��a�]o�24���X=8ؓ���r��[��'��b��ˣ�?�g�>O�1#��Y�qh�EB�Nb�$r���g�2�h(��E p�/a�n=A&ḣ�8���o�Z��X8O�o�P�����B�W���6�{n�:�f�� Bll`������4x��l����I�	{f*L������L�FD�;G�6߅�Z� C��^������|����81zJ��3Y��h�P;���;u� G���#:����Q'�&}�
f��R��Up��{�������)��)ϡ�A���w~&����P{��徾м_.�?�O黂@�Y��KH6N�D�	�U�����\f��}x�Lb�ҫBҡ0�����7�q7X��A�+��g�C�`u���iH\��]ӛHM��~W�Ʌ,�C��A�0��qN��[�K��1{�K
 "�_ &��@�7��I���i�-��Zs��	�52bJ>�����@mG�R�=���g1��"�����ɗvVӜOrp0_Fi��=}��ݘ�O�]'o���%e�/A�'��D�:��זl
<7$��@�S�)z�����S�[�� y9'��ֺl�y��W�4�L��X���!�1Jf��wZdU,���I�\m�u�9�n�ZY�c��_����d����u�w��3���&�Ť���}���,�҅E< ��N�gft������J:_�e�Ĩ`���9D��=H����� 1_��b�e�Y��������k__���g�w����'@��W�H�b�m���5�9�'�k%�������4�\��xz��]�w�����ӣ�k�r5�b4R�,O^W+��)g�����Yh��>c<��盲��-���������4YL�����S9y�I h��?�X׷}��� ����C�<�=�#���e|~F���	%��-]�v9�!{�78~Vd�e��!�q����`�j�{��G�<}�D>��#��{�����d�#��2]������kD(NO^�K}?�8�	Sl�����j��u֫�?�,6�ǹ>7��ںº�n ѠN��wj��$���Us*���&�Üry�% 7a\A)��B��B�{�ȯȌa�
�u 	}�� rg�7��,����N������؛0�F�x��x4�/��R�ھ���{��5��ׄJ��/��E��3u�y�1!!sr��T;��~�z����zK�z����y��],��cx@C�u�u #�Aͱ1��X���xR1����l p
8�������,y#g[�:ϘlU̏�)���׶�tL�NB�\��! ���1�unh�dS6eS6eS��e�lʦlʦl�o� @k��|O��rv�z�'G���B�&���zɃ�s�3)}��I��a�&2����j�%]�%Y��a��/�x(c������+�N������ ���D��<��N�	̏8x�����]&#���0�3b{п�F#9.��湁��׊�.K`����CI��tjm4����S�1�!��l�z��a�Q_�A��s���%+A  �E�b@��:<�V�� <��.�3`� ��� V
��$��^H��L�<!rAX�In�@k>!��·KH H�����b3��hw�۱���|�k�"��
��1��#���5�]�r�/W��2���m��t�r��]�j!��?��� ��������0xLa�9Ե�4̯�]�/��tLB&���Ȯt���V�&_}��I(.a�2��L���@�i;���U��ƿv���``������kȺG;�=4֋�e�6e�9��4d|�S��<���J ��YQ���O�,)���{�M ǽ�/�I���� Ѻ���	@�t�k��'�����>@�^[]'��S������F?�	pA�7n��۷	z�}�8���e��\~��f���ѿ�?�1|~~ʀ�����A7`Qz?����i	C =F�g:����a� 3�Da�^.���Q��`��y�J�(�V`Y�h��e��{�djde"��Ȋ�3$���Ե޺�{�g7ֱ����x]൤�Fpp E�O��rx��)e��CdQ;6�� �����Uc����Q=ge�?3Zwu�/��g�M�&���k�DJ���Mm��64�$,'�����Xǫε�%����}^Z�m��� ��5�S�LV�e;w�o ���I}��q&�r(�ܼ J�s|,c
s�H��N������:�ևhCn� �f��r&�ٚ��q�!;��ˈu:4`N��۶v��jK������#]�<}�Ɩ� @����]IW3Y�Nl.p�Uк�a)́��b�~�?)[��Q�0c ���}zpy~_z[;z?}�δ����m�N^k <�bUm����˻;[�l]�"�_r~v�~S]���_��Ayf��SYR�+p<�z�g�����`�G�	vR�;<�޸��%&�c�B�߉�,�P$`6`��u��
g�}ok���^�G�ý��������<��o�#�y�}���R�:C�� ��/?�=CZo�k6�Ώ���@�&�O�yNV:�-���$0~�(�9`����@4�0JTzU]�d����J(������<����+&�XewGn޹-7�_�1}.%=��"S�4��3��9�i�����������k�@���3b����H�m퀐�Ě�l��L�쓘�D~�{����lJ�ixr=z�Hvt.�7̓'O�'���fX��X̗L�;m��1XF��R׻,-	l������Ҕ��f��<0f�?`��.a��dW���x���A�� ��ٚl%2��Vq��}g�d����MN���_@��ϙ������@�\.�w �I؞���߭�!�:Ƈ��=: �5�
�Vb��O0�d�A�s�l^*9/E�c��q��*���G���>��%�V#y r�&U0�H�ʣ�}�KڔMٔMٔov�  ��)��)��;U���,'y6�H��a��Y����4�ӡ���|�����A����2[�E����\>����8�1L�q#��'�?
hv9.&�Ǒ��P�MF��y!�ј@JT c���R�f>���0X3Ӹ�ky�YL�$C񞯞>��>�H�Ǽ>z�V2�/��Q,��'X�ǫ���?N0 ���G�����48,֣���ly%YT��5��Y��CC �\�}Lfӱ.Jʂ�@� v�چtjƬ���l>%ɢz�yu�!�����52*�!���4��B ďBf�3��W_})'G��}�j5�'A+��4W�f���9�i���l�ʝ;������K~��}����5 0r��ԑQ��g_P�"]�L�� lB/�0y0ov[��Ff�`�,#��!�d���l3���S���Oą��7tb�a�
�h���{��X�b+��A���ԅ��d�/%���<
� p�[��Re�� �\2���6����踒.�Mk%�$�.��GQcəˢ0�ٟb��`� ���rhQ���@��� ����׺D �@��:���LF�����ˈ��AP�����`$ �W�����S��s��\�f~# ��>�y��rm�Nf�J��w|d��3�O�~n�{(9#.�� �ɺ�a5nb2@0�+y/<���B�:�����xm+ehL�¢���}��^����zS0��c��e���D�q)�#d�������#�X�FB?d�"�\6�c��>X:�w�4k:�̥<?�TS�����}�%m�+�'˅t�bh6MT�.��)ޛOE^uT�w��Z����P�"��2v��� ����̜�b���h3(�D�;R`˪y���SY�Oe[%3eC2	�:}�D�vb}<��[�39=K��:����]�
�1����eU�t�dZ�z�d���|D�\�-m� �u��=�j�KS�ۑ�u�l�@���dI�.�~Bs���`�]��c�_\7h��t:Y��>��R����`��O�=�\�=��2_2��*+����lB���;�4�c#	'�o�y�����ȍm	;���o똻b�q]�2�u_���S�Ȃ�A�q���s���v��4"�ϡ2��V��\�Sޫ)�.��Ȧ����?�y��������V'��1c�=FV�g�b��QQ�J�Rf`E���1xi$ ��A�픠S�`N`��3��O�.���Y��&�G�� ��}.g#&U i��g�s��u�0�8�����V�{�����Y�.u��Ԧ_P��$Ȃ������LOd��Us��zO	<t��<��{)�ut�h���L�ז�����ӛ^Ѹ��mN2�Y��a	��w`����_���_j{�έ?� @. zJ�&����K��Da�LlNm-�B9�x�!||�����S�EbZ ��g����	B ��N�}	 �ʲn�x�M�O:�'R�X��W���)�D�HH��Q�[]&�Z�:'ʧr��M���;�6�K {ν9����8INDb���8~�� y�H���M���ި����U�`��ܙ���{��s���w�ޓ��ۜLF���0KL^�����!Vu2i��DzgN�;<�O�/���(���W�76�cw��.+�T�paF>��E�o=�5GP]22�@C��b��N~_���]go".�aS6eS6eS��e�lʦlʦl��D�㬞iS񐹾^�B_Ñ��s�w��$@��E��,d��2�>/��ή�o���A���;����Y�^hy􇘭tff(��A�$60�ft�9�d
�(�4�Y� �s���wdoO���L5��-prr��yA/;�Bc���R��������KOF��	�X֝T���D-�i��j�ݻ7et>���A�%3Sgd{D��h�����Q�W�^�P�Y�N���9�.���̓�f���@0��5ͮK3-�1�oL �Q�;����^��=2$h^�M��0i�/ ˴Z�j�5k�?HZ��w��G.���*�_���</){�:@����� �]MZ���l�8��o��Jw�P����[r��]�O�s�<_��²=���'^�P��?Y�8�SW�	&��`Knݾ)��@N�_�tz�}O�ݟ�lw�� ���a�~�`]��"33�܂�Ve0���f�Y�!��*�̀>7Af�:q�@��5fW�t�#!��%�v�x�I����-Lrؘxp�^�ʄ�fƥ�q`���$Y���M���4��g*�ŀ3S��;����@�}�]z栠�`�{vqJhgoWz��15`"��X;����Vh�U���`�����Ǭ�����@�m2��<i�z��4eY��ڝ� e��t��y�{f���@��򔴪�'��@�y%��Λ>��G�?�X,���k?c��ȫ*�4}4���̤�l�x p,4�EBz	�|�f  lQ"�X�Li�70y)����:����h*��W��ݓk7t��� ڄ�-~m$am.�Z"�&�̴�.=�⠌�ڌ�b��K_���C,@����$�,$�a��=3�IeA|N��"�H�_Ȯ~�d��+a9����YzJ����v`u����#�:v�٪�󳱜A�Jבzf��{ ('����Sm�����# f `h��:0?7_�"�e6.�.s ��\vW��4"�$Ժ�"���N^��S���{%��,a���P��Ი.e<�p][.��:��~"�/�dG���J���t�������-߰�Ʊ��k��W�� h*^�8���m\�@��ߖvs��u�*9/yi�`y�������� l���#X]�s4�)h�]���O��_I��:i~������!�zKB]}�9΀��2?����c B&	k�*�>��������$�p��m:[����`�u�k��t�Ĝ�u�b���_��%�R� HS&�՛��?��O��ի�����������G�\��&e`��v�Ƙ B�-_V��{��Dr]G���.�ϣ�
Du�X�Ebk���$M�a|��u�c�<;9Ѿ9��ƞ�Tf2f5�7�$i':����X�|ǾÚ
@����<|��<}�D|���"�`Јd��_z_`m�\n�B��;u"����o;�E�WfNzS�m�s0<B�a"���� `쀩�u2vσa����Y`���=#q$I'd�ֵ?��c�����2��l��$�}���lxsqv����4M_�W���u,{�+���9f���y�uPTs�`�?RbJy�*�Q���ϱρ|��ױC�7�� ��-~d̮�IQ�W\���.��I�'1���@4�h �F�5P�ҁ%����{�ı��~0��q[�� h�/�po��ד��y�Y�	�Z����ƾ#M�Br�?�3��:��\���a%��)��)���. dS6eS6eS~gJ�ѓ�l�_4�#������G�ZԠ� ��x�L����
=��!���/(��m@��{۲���~��P�&�y E��p�*�K�8�)ݭ5��k7���{w��z｝�ܺy�p�g���'�Z�����L_g؞°Y�2y��[� y��@���^��J��<��S99�s���h��~��C���3᱁�;�ce2a�-��V�IP�y��g!�Y��O�8�2;3I���i�@"2�RT��wf�tz�s � ���5� �x��䏌����08��q� Y�crɃ-�o��e�疭�lD�J�蝦l�wxp�G2�Le�vM��7Z�C¡�SZ�Ȇ�L���ݻr1R*��L��J�[$��<~����v[ۙ�)�r��Zӹ���V\�z ����|&gg��"Y.V샸��w~��e��H��uV�q���cϟ0�6s����������z.UB��=�5��ÂT�**�����-�PE��Kp�� �����\��~��C�	���曌�zM`��4��/��~��>7oߑ��yG��ַ(cٖ�r�`X����=��ƪ���}�KA�� �M�w{�|�F�/'�lFƬn�B�'d�DN�#�*�)2m�$Y�9��cd<[�7�=V`�����1�K3P�L���65G���C`h߂��IV��}���������a��y#hMy���y�}+�q-�� jb��B��z��e3!���M�+���*��j)���?��*K�����r�9�P�d,-o�@u^:X���)	�$��g�� ��Lӫ�`��R�r�Y*�>��B3�Ɯ?����5Kf2�����~ٕh�f�\�A�%ER�1H���c�x¾ ���N����l�������4�k�D�/����ރc�4�;R/t��9.K�$�qc��f-�6 d�G�4��8��9שD����ѹd�3\�p�Ciz�.ϴ�ϵ��:&���c�EեK����X�5���D��_���vW�m��_K�+-P��&cTk��}*4 �x݇�&�){�����@��ηޗ�[ߓ�����i�6J�n٢ ;/)R%��6����̑^:_#J�A�������}M����W:������g6�	`����˂�{X��֮�-���F9�  �~n:�Y�+ lLV���ZRb�1�`�������ϗ��`�����
̽��=�T���5!��չ����ڵk����s�;�%[����<����$dZli_�_?��~|v"��k �#�O���jp�Ӏ�E��z��0[�NJL�P��e��-��ޑ��@��Dפ���1�0m�&�GƐ�X�X?q�Q&��5�b?��?� z�l-�:��~�r�h_l�Ejo��=��d&`�r�@���;r��m����h��h�c|ʾ�Z%2M���L�<}&�ǧ��Ϟ�5�LFu�\N)��pRX � nab��̵�[Mm���'`=��/��^���+�uG�C��t+ /ȵ�uca�ǟ�G�S�u�O�7���{� �{?(�����q�Z�=�C�!��ׁ&i�g_��D�y�CojlRZ�� ��	0#�������̒`�g.�\�(9E��^��3?`�����%U�R�u1�w)��{Ĉ��a���:�Qx�q�0Nlp����T�օ�cRc_oȺa�oĕV�I�����V���_dS6eS6eS��e�lʦlʦl�o� M0���r�р�tHF �)���K2��e�B�Y�4`������ z��|s���� ��Va,�A��7D�u�@F�2�`���P�`���� �rJ�lmm������P~A�#ó��n�8#�d�df'����y@B�)2X�ͺlo��p��w�Pi��d!/^�t����,�Z�E���K"@@	Y�[��~O[N���m #P��s9���^�M҈� �"vqOtx�L�g���2�Ъ�u�PF��WI������^si� �O��@vK� I�_��"����C�ΚG0��������<�s�P0���f�%W�\�{�:<<�c�Y� �Wqq����A�?2B��]���������`�fk��R�z�~������?����9�FK|��hc�IւW��뭆���u�����L�{���j!��1>
E^豽��34[5W裨GH��������c|?�;dCV,�T���z�jE�Lȟ�W9eID��֖I?��A��^��w�9��҂l#�* pQ�����D�g��lK�dtҷ�`�ߋ�\���H��c� <�D�e�a�ϑX� �hͬ@�	���]��4���Y��\D�����HZP
��������o���p���@&k��È�s��2��fx��b V��U�U=�4����
��S��c5�=[`@�S��y��"��p��_{�����uF�|�+c�u �����"D�Ć_��ج�Y�1�,���Z�,;Q��Z���!�4�Hs��V��yl<��K+0��ad�!tAt�3�S��z�+���$w,Q�6xŔ��+���2�X��&"g���}�&�:���}	�l��%�ەfq��;�T��W�P�h�ɀ�d��D#�O�����d,�>�X�U&;�2!�����lH-�>cwH�	��0J��<��.����z�նԟ=�>�'�O�ƽ�<��	�ɷu���t~;��t�`^�2�E��^�Y,񧵳_�d�L�0�q����ʄ�&;�m�g�WL�Vu��I?�����{��QV$�������߅9|G�U��$PdqGdDiҺf�6�#���� ��ܕ���et�e%�;I!����40'n��DC�D3���F0z���i��8�1���tG��2�ɒ���I�W�b2Q(��<}/�At�)0��k೫Õy9�_�Ե�{����c󵎥��sW��Yg���t��[o�w�W�u-�|��|���rvz�펾� �'�<��Lܸ�>���C�30�{�����P�o�ݑV�iI���W �"�{�z-�W���GrH����ز������wt�(��i<�S�k�90�z�e��	^/7oܖ���5��Z-���}����'?������9�`�j�d��Nf�߸�'�g���6�.~`�G2 �5��tΊ$	�e{kG�:f��^�08Z�\�~C���{s�7�o����_�Ge&����T�eF�`Mf���Z:��8��S0_#s%�R��lHy����(NU��*G=U����_/d)��R��$4��~���A�{F�����r6�paI!�GV1&�U���}F����c� $�����HF1����1�� �u�~Ϥ������O�$J�Y"���'����z�a�G�$:�~ש��KF�)�ǸZdRY��,�~�~Y���MٔMٔM��l �MٔMٔM�(����ٓ�eD$�G̬��K��L���� �b2��vI�S��y��#�fq�.x/��0�F@�g�wƌ3� �v	�_�i"��e��lE D�܁̖�C=�����x�����
�"�J�z�?�8u�KgԶ�7��=9:fF!8YB�ׅ4V�Pf���c9:>���s�/2����'rz�J�z�O�\VuX��SO�^��D��T�a ���SZC�}�tA���a��`4�q`��.HV0�8!�A�v�C�+�χ�:#���F�;H2�\s&��w�[a�>U���o�S�5�&o4�fЈ��0�z���{re�@����^"M�	��i���LF%A�41���� P 3�N��@����]�%�xO��*Ͼz(_|����f�G6��� T@`���E�^%��Nw��F3���	'�g��B��l�4q#�9���ܴ�Ų�+�<��d�⠏`> ��95��o=�=�^�'�GNٽZ��؛"`�@��x�����*]�)��d"�I?ч"��a�~->eT(͂ E��ϾlZ�~��TNp$dڠ��Q�3�aT���cD+��`~��Q�ٵm���`�a�3mX�"p��SkԨ��&������h4�t���y)�#vG��'ǐ	����E�ݐ�������� ���Ȏ���L`*�e�`k�(~d�/��rrE���9Z2���~��>�}�&�PV�Y�م`�[���5M&��hIRΉ��L��"�9zB��d�F �E@���d:�X�Wǲ}�t{����%eP�Uisq~x.Оf4����B/�����9���Ș����7�q�:�������3Y�4\�5]<�l��k�r=��v>wR&�s�xy&����z����E":�j� P�d7�j:_��r�m5Mezv*����}�Ʌ~׈� �#�G�d�p��%X$����� ����`��|��=O���/��*}@�X1sه�cR�uW�g Ҝ����0���b�_�ڦڮ��Q����ʎyA���ɩ	3Ա�UsAEtBecI�}�.�����l�2X��o^�1I[lR
��>�o#�f�*�j�/zo���!���b��GV���	�����7�$��Ğ/�{D�������pHj��:���F�f(iF���&@�$�������c��E��g��@����ITgfd����3�{߻�ՄXo}]��ŷ���`MB���!֎f��1�&���M�\]]1����|�}@�q\O�d��xo�W��v�1�/d�V�R&S�`?*L�e�#���~�+�l��B���bma��M�Tf4b����������|������䧟}�c錒��N�����@�S°f�3�M��zj�I��>_�i��g��8	w�L4YCJ�$s�u�$`�*F�,@Lo蚻/<`x.��Y�D!q��!�'1��NO���ɩ�݈k
�ޛ�Uf����M�לի�r��y}}-�0���>��-���d-b��bV�y?ijRH�d�H�ृ����2jx�]�f��zN3v}�wNO�~sy��\������~�h<�t�о�9�7	5x�vwu�/4��?&7O
3��~�_E�� |�ba�+�F�
����H�a�$�I$ �p}�ߪ{���n��9� GZ����X;6[��ǽ�	X���O
��XwlͲu	9u�w8�1�F���Fh������Q��}�6��t2�Ŧ�D̯�Q������&�p?�΢D�G��P%�1���	o�{������r!۶m۶m�mK�l۶m۶mۯ�A�ɞ�
��
�2�MiB 6�Y�^R�	Y���_<`6�1_CJ �,�׃T���Q��6Y�?;�1{82�ϗ�v����AHHB��T+6�o1Cj�'�y�fDYxH�^��8C�z��s�C�0xyy�u�!q�a��k�_ �􃠃�,p��4Kn7Y� ���Ꮌ|u._�L=y"W���\���0�A��H�h�ì?=Nf��Ŝ�چ�ϯL� ���PNs��K�7��  � i@ �� #���5� H�A�	`d+�NW�z���F ���:�Y���!��(Y�Ѽ�w5x�q���}f"k@��gu��}~`��KP<]�v
�5�l[�9 6��8i�0��7���>3� ]\\�x:a_�A�uҠ�3d�|ٻs,o��6M�/G����3������ّM�iS﹍M���^��G�*�()囶�'�Z3��}H�4J�.��� @	 ��:Q���������X����oNi'��+ �#W��꾍_��C*�8�����8y2G�TfP��x����pG���X鱺�:H:��*�r�Q�x�2" �P�QC�pƲ+LS��p�øo#�tlC�=��W���\�πd�r����i��cf~�A d���o�.)����6֡�r���W�S3�� A5��xxS��b��@ۑc��Uk�.����`��&�s�����'hF�0<�)�������,���R�;�ߍ� 8t�I>4t|��#�URPfO�X?6��,��LF���_��bɹ
�(����	*�6�F�Uf��<'qTf�89&W-�X�;��e �����g��Z;�1�2!�]�U�Y�D����[�i��g��L�O%[���;:�5��b|L��6?�
�[���2I�D��2�غ�F&��u�;h赌��o��h�cČ�s�H/��/"�S�1�0�fPмyr6��h��y!�^I��<�H����
4��d��H�@��[%�bb�\��0�+�A7�qm�y~s���-�s,UfJ���~�j�W�׸*#�D2V�e]�����Q˳uq�4Ұd� d*�e� ���ǊH&P��üD��Vs�T����)*�Vk���:��4:�bF�4M.+�Xd�W�Y긮�5�1 ֹ��uq l�[e��鄼�M�].f$H�h��}ҡ�i1f�FW�EU2��Z�����,x��1%�`T��4Խ���I�
H|�PYq��1����u�q%7�7Fv����V��^��s�ϸ�
Vxn���9�չ_�:zs=�/�Ɏ��Q2P+#�DnЇXP��&UAF��^�=d�h����%2�VW:f��(Ը�9��5�ïm0�o�X��/2\�lI��`�s�'�SH����Z����x6��dƘ����&J����V�ch�����s�Q ���ѱ�}p_��C��#S�T�6<c��}�=��3�e,3��%�0Q���*lM��� ��\����ˣ�H�M��c�4��H��*g��#�ׯ��/7���燽W@��!�X��:�*�9*��s��=�c%�S��F核�0� ��ê3a��^��5���<�Á4u���&�-H`�½%���NN��۾��8�=\��-׺ҼX
��~n��-�o%/m��X=[;�Ԝ�"����Zk�W�_�"W�Z�/{�l۶m۶m�oF� ۶m۶m��Ϫ�`1M�N�8�n8@��P��dP2=�MM*�eX��z��q��c�����<�_^��\}��YZ<Ɓ`P�f�$ ��{迯��z��Z��#Qpy}AY%�C�B��Jb����L�v�+f0���=�Cn��� �2�Ι�7j<�Χ3f}R����K�Y���<���t �<����H߯�iQ.��f,�H�z�^�V���LsQxdHL����RL�>!�'}_���LU'+V���FCn+�� ���Tq��B�L�;R뾬�K �á�GC�i-7�9�;{�A�����6�2���hB(�X�Ԭ��:�a>�����s�	�ތ�e8�1q>s`��!�T��6�ƫ$7���2������O�ra�┚�a��c` GG;No>���Sy����Ƹ�0˖`�����|�^ʰ����]�Ϯ��y���d�����}��9��2�N�e�?�&(3���i���"�~AeS�̯7�� ���L�!d�AV���( �	�Tk��#6Y� ��� �`��J�e[���K������ 7M��b�(ޤ�(PQ����H�z�C�J��5�a`�[���{��@{?͘�Oi�"#��Z���b�lUf�0��.g����ј  ��OEɬ��άa�����b�o�#�Ɍ�%�8�=nkl�{P�B~9 �q��*���4��b��s�й���P�v��8nAέ�
�Џ$M4�1l�8�:X�a�=�@���k� ��i��V�ՌL  ެ�*Ec�r�o�[5V����c�J���-d�� ��Y�e�V�����B�L�����+�_S��	��b"��J��vu-���e5����qT����!��A�i����
8P!Ar ���d���)�,�0�[�I8,oM���jZ$ Go�E��\?}"�b&W�R�rĪ����@�߅#�)U�1��T�G�4���s�+���L=<�z�ȥ>��g:��0P���揀�l���<>0D��1 �V��Uh$�ٳ�2n�c] �_oG��k/���<��lImLD�De����kܪ.�'z��F6�"a����CH����L�2#IP�Xq��W+$�=�x���1�'$OH���C�s��Ig�F��8r.s>	!�,����T��'mX3� T�5�����0���r�@�:	���%3�a5%$� �6�x���[�^W"]]CV�T��
"���,���2�t��X+//.d�k�����m��S��:�v>���'7�Y���K�����<�C>.��|��ƚ錜g��j�|#2_wI�<y�X�.^�t����zԉ$�V\�6�2Q]��M�/Ϯtܷ����
����"k3�Ji��TD�ܠ�#�{�eB�
����o�t}qMp������٩�4��$����0��O�3�=�R7��$-wv�)+��v9�4ѹ6P�+�W���x1�����S���Nt�0�>4@�o��h"x���'���c��k��UԨ�:�W�sC�� �Ȝ�c�6Z����)���������+���rx|L��/�������%����5�r��H��%_?�J~�ÿ��j��!�-e��J����@5T�rz�f�UNa޷�@�AB�V>�L�Q��*� �c\E:ϳ"�O86V�l��_&H���㪆Շ�2����r=�t��!� ���lr��,^AK�+*A��9�6����g2�-�G�fU��U'�H�\[��j`}^���@vz���HV�r��0�ɵ�(�����B(�����~|˰g����C{� *�X��օ%8`9Y-T�U�I�Mt}�A~�ޑ�������ɶm۶m۶�f�-�m۶m۶m�ֶ�俞��Nٓ0	Ye���0��C˚DU��2�Kzj���`+qO��6f�q�,�����<���擐h���o���6��T������M	�x���m�R�����a7_W̞k5[ԇƵA����>s2�{�9�������%�p���~_z�~p�T�����J.��(� �P�H��,�9w����L&cfu�a���� �����HउLW���E"3$m�1	f��HH��`�^��rX�~=�����[rpp(����	�2��)O3{ϙdC�Dqp��4��t�=�$��H?g�Ye�V��1A�ʥ%�f�l � <�� ��W$%�%���4�} s@��R�A�yrT������q:>�@��H���|G�GW2�����WW����w����;2�'`�@�f��Vv
����|��)~��V�)�H
���~R�`!��*��gn2KV� _�� �8�^#W�<�:��( ��L�A^����?����MF�c�*\:��xV��0mh����\ݑ,�� F�� �" A�Z�DR��5$e�' j��#�yC�P�mMP&��@(��a�����=�|Vo�}y��4߁�q<�K0�h�RZl	=G����������Lք빛�3�Ie���"ܱ�<hf	��h*�/�E�	L_���3�o孬�!�'�I\��$���=V��T
��L@_���5H���=����ֆ�� �&x��F�J��[VT̬��L���eN�/��\���ɭA�*3�3�dH�m�|,V�̬���*H�Ӝ�L�̫�_4�vmSi�8-�P��e�QMVX�5לN=�7�$C��/�4Nx�Y�;��vg���q��#���;)Ȋ�}A� �l��W]�r����
)�����I(|���84.��2.,�ɍxh7P)gϜ>9�H�U�t��Q�*����[�4�Q'aFߦ�$�(�Db&�
�3FJ�"���J9/-N݀q�Ro�y��������:��'H5FK��S}mΉ�uzo�f#f��+�%m\�ꑘ��u�Z��AvO)e�:$���R�=5nM�S�e̹�)��:�u`=�l�C1�P��
"VT�/d�r�)Ԡ���^��1�7�	�IXS�3��U����}�b�Y͌�ݺ��Z�L�s�G�	)Nze%Sk�^Tę����yV9
��ų��s`��Rb8أ�%~b��,Y��`���w��A�䛯�����㯿v�p�ׂLB����#/���;G173V�h�Ɯ���LZŽ���`��=Y�1�؇��7�{�3�� �$ye�;��X�ON�d��d��sxڡ�,���?��V��O��� ����ﰶG��,3艂J%�������孷ޒz����60��w�m�:�w%�΍��d|#�''r��5��:라*}_��� �2
���| �U����Mm��<Η�$xۊ���O�d���Cŏ{OT`� �P��Վ\��}9�\bE�(�]�Yͦ�Us��x��3 �0�0��nC��Xl�|-*�Z����c
����^�xb͞Ũ��v�o�}BER�w6��s�i�e��n�&�q�ss�q{��C�E�&eÐ^7���|�6۶m۶m���׶ȶm۶m۶��h���d܌)���2B/|��Ȍ�$���� E��5ό-��\���enw��.�� ���J&5�� �5%q �3�.����F�#y� !,d�w]�8(��= 80���0�u�k��4��\���B���2��e�̙!��\_�$nu����ߑ�;��/���?���md�EF�@����Z���h8l�k�rt|$��>'!�c��i�u%p(I��`��:�_��_� �� 	�\�IM!����ߓ��=����t𻨶�J1�' Y��IL���D�,�d����y4�M����L��Qȿi��L�͈� a\�D�}2����f�d� _���������"3�I����W�@E �c�s�|���r��Bί����BV�y��y���ސd��o���F�I����u���,H�g���'N�~ �~'�ja6��҂�ص��h�F4�wD
�{!OR�FlQ��k�}�6��"�s��0�2R�ɥh��꿳�5�ِ#�^UR <k{�q�����d�/���ܑ`	B+�4]�ϕ�-�� �QT�k@iMƇL }B�$��� ��AP`�"-70S����2d ��!�1c�������y�����?#xZ:-!�^���N7FĔ0L��Cnn�1,l�$4Ι���餆6��"���+˒�q������Han�נ�Ç�{�1�����3�+�W��׊h�� jٸ�G��U Vh���I�2_�:;=��.���$��S�X|�$��c��
q����C'��������H_� ��Z\7(0F/�e��$��la@^m�F�z��� ,I�(����䠯1}_��J��Ȫx$H�1�N,��@[o�'�b_�������~[ZM��>d`��+[��hUFt�k�!�E��i�
 �!,Zt��`��Y ?��:�\�|&�N.H	"�;�U&�Б4���/�Wpa��^;�EnDH��/�	�J뮸��/zf��%`tpLa�u��j���|"i0�u�+��`LgzM��GH2�L��|��X1Z��������V���k@.�3G��5��(���*5V6���
�ݍ����`T����˅\UC�w�ٹ��U�5�g� ��~O׃:�'�r޺�n|�ڭ��1���V�>^�|��,~jG�Sz�,�5[���	�k�{ �.T����%)�C�z	��%ڳ�R�>{.�v����������M�[��VV���ق��������9�'o��.�f�8b�d:��Ս��-� �3�$_;�&���=���cRfqq=p�Ӧ�r��p����-����i�@L��7����4Y��S���m�~�@���Ր��E2���>������HW��+^��V��7H2��5��z"�a��$"��s�������F6*��o��A܀LB������W4]�ߚtZE�6$c��$����_
�q�m�$�%7^�10��9B�W�_��C*5�l�P��e���w�W��a���7�����U$5�t}�(M�q�����{Y.SV�;R���%`a�u-����jW������b=,�W]R�qqI+��ؿs���-�lS���:�Ã}����*���׍��dr�c6�������.�'��'������B����l۶m۶m�ov� ۶m۶m��koYa�:Sht���^#��. i �8`#���1$���6��g%Bᣀ$C�j�-+��+#>�5�3�z���8�^?��p����P���5�	����Z�'����_\'� ������q퐢x��ү��3��������g2�L��ꆤF�ե��?��&��E���'' �������J��ٕw�ޑ{��2��ŋ��㧼�uf�Ʀ�?Y9Ҳ�E6(���3����A�Y� � 8���S~@� ) -��y��8��YTv��׻�2� �B�ڀ-� Ԧ�^�gm���Hb1͖Us8�f�j?O�cf�Xuۼ>�8z�����ې!�L�̞ib�*U���y2y,ϟ?�x<=9��ܕ���˳�ޑ�d��lJ#N����]�B	xX�{]��,3y���0�#G�QVK%Z����Y	4�Z�*c
��0p�]�Y�3�T,��6_�C��D֞�_Q��#�7��x�4.wrRU������b�����$7 �T��(8�\�?,C����z��P�o�����0³���C�Ԟ!�S�ތ "P9��KI���7	~��%%�{�{��D��.�T�0�Կcxm�H�����*��Yy�IK�����Ћ`������X���rI>h]����ӆ����}��?���U����]��RUF:�0�$��k�"]yT��j�V,A縡�x�*Nj�2��AӨՒz y0��y"�ťTA"��0�g�L�4 P �&5��,$p;���?�iGB�ϡ'u�הZ�&IU��0�p}\�z*�o�c<�'�C�*%�6� y����FE�o�6�� �<���gt;�@����	X%!�9j�Im�@_ܓ�!�ɥ��P��L�I�k�e��(���I6���rt0�t�X�]��m�=���YB9��ZI-�Jw "%�%@���3�լr��X�{?�oGH�w��	B�AsG�:' ��X�$hFK!�P���*�x]+� 2���'���H�
/#|WE���j�� �m<h|V �[D�c�auK<�6�U�џ�B�UTT$I���k E	^%�bJ�8���x�e���zŹT�V��ױ
�p�8XG8�gc���H^-9�{WZ�)���Hl�R��j9]�Z������ �)��U+��u=d�]j�[zV%��A���ށ΋�kՋ�O���'���cf����ڨ2����oai����-�<�*���y�/.�s�a���	��t�;<d�ֹ�^{G��D53��� KUA�Ľ>�K]� ��� sp{�NW:���z\�:J$:���	�*V�B·!�۸�9)�
kOXs�e�PA5j�W��3���h_�x���{%�e �w:M�5�����~���H><����fB"��6^֕U�����`���2�0HJ�Lc]��2����U�xf���Oo���+Pu?�W�^��+����|��B� TaVF�.�3ʐa��m�{��d,q�-#�>�n���׸[o,��RS���ۣ�؁�/�q���H�d���Hl�E@� ����;j�����z��~��\�A���0����������眳Te�C�5-pg�ѵLg��r��T�~�+��2��O��jx�h|C��:߬}%�OvC���o�'��:ޖ��}�����?����=4��Y�
XT'��ߐҩ������?��������m۶m�oO� ۶m۶m���oef��z���!Ȯ��?L�E���bE]=�9����g:� a����0�!UB�8d���A&\-69�O�Nz"�A��ij�Z��Aq�����U�C�:z@�u{�L�srW�����`י~y�B�(I��F�uh����;�&���6���L�=},O�>�O?�T^�x)�^��1�O����5�~_�n[v���������^�Yv��ϐ4�x  ���zܠ��\���#�M�N$ '���9T�̠�d�Ӵ[�2`5jJF�UJO���4�)+$ӱ�=/�9���I6�r3LK�ʒ��:��P�G�g�����~u��lI�d�
$�pu)2
!���zD.�nXq�嬼i�$�Q+UkJi�6ʰ��3�1	P2lo�^�ꫯ�����?�#o��|��3��Ϥ��<��+�(����m�@��eww�Li���-pM�Q�
�.#�"��	�V�F  ����9�> pA�a]��!0����_ȝ�T?3��]��3��[�%#�DB�4C�M32�#0S}�ِ4 =fb����(���̴T�c �:5)��:��r&��ز��3 S_d�f�-��
��_q�Ep�;�[�����o�3�UN�
���x$�����&�uT�q]%�[8��88=�?��?���K���Ϟ��SQcK��
t�����ތ�A�xK;��&��9DĪo0�O�Ջ5�=���5����J��Ƌݤ��E��P�cO��݁,Z����j��կ���T�ЌʫI��.2��˙� �p�H�H���蕵�Q75>z;'FЍjru�����e9W�3�6�X�x"F�Aҫ��)��~ict��
A��Alg�x��W�s�[]�����A?��ҪX�l��AeƎ'�����A�xxO�����Hk�}]jK�+A���; �"G�����\��I�X�⦴�HP|9�Tc�ry%Eh�r-+0��:�I���m����t�Sa�Y�'�.
x�Kgؒ����{,uz�ƿW�aVoE��g��=�JY,��^ �.d����H���(=VVIo3��#�\�{.|AX�F�	��W����!�V!������U�b��ɵd�ѿ�t/XQYQ��O�0�q�Ճ%o ��D��t$�V$+�uP�����U��S�6_�op�	'�Bx+5���@:�LS8��5I�N��qy �w��d �B ��YG�%�H\�FV	�A桵bv<@�v�#���/|mj,�<�k�S�O'/^���r�k
�z��Xw!u�km�3G�e�;��vy�0���ȼ�P�jv�� �CX�f��{L�sy}v���\��������ms�5B�����j�����Ř�Q��|;d> ]Wd����#�|�s����!W���P�3+�oQ��׉J���7ٟ�}0�#Q���GR�@ๆ�~�C^L�2X��X�����X�An��]��&��4�`��\6Y���,������/x��k<s��~���ߧ��Ç�t�Z2���7���oT�h�yՠ�V�"�_T�I�`�Gi^D��L��6�YD|0GX�d$�X��0�k�l������(w�Jo0`e���g1A��X����g����ח7�?� �����R����F2�%:�F$� Iy}qN�G<�;w��;���y��Z��+]?1��uH���*�1��B����*�>��c9��@����e���F��$T���7j��8�����vk����Qx�����(�o�������m�öm۶m۶��-�m۶m۶m�֖esy~~y�=$*V��t��*�l����:#`	y��e�C�wه @`�lR�e��e��̅+H�D�,˕,晓UNL���eLX�g��lDx^v�rr�U��G� �n�2#��	��]3����մ?=��PYi�����=����T�{�C��O~"��/��|��O�铧2��$����{;<������!�V[Ȟ�:�6�3h������D.//��hZ�Ȧ�	;<H��@q	�F�������Nd$AI�� &�Ip ��'��ʖf\�!  �
�[%K�U͗s�hx��C*��0�~��|�,���|O�=J5�2�]V��nHP
�	*L�o�����B�H�1��J��� ��"�g�:�V�����(Ä�H�볟��XM���i��R}y�Z>��s���;�'Ϟ=���� LB�#{�����Z�����Pvzz��#�H�����̓ax\P~�@#�`���J�g��$	|H�|C�'�p��E��
Y4�����V���Ƞ�F�$��P�rv��*�7~�����)��FN�r{�u���#g��9�v4<�LO�<��u򾽘��|�O�r}u)g��e1�&ŹV�|V�x�F��P�J��4rM��΃�M�`�HJ��<#m�q+�e�S���}���ʟ�ɟȋgO4�Lt��(=��G��oٰ^yKmdb<���,yA�9ϝ�S���0b��h�f�Uo�V}׵���jC�t�e��c�T|�a��X��&	��B?3Mt��g5Q�ѕ�a_�˞L��hl�����D>|�FRN�b���`�H=�m�L��������*|fu]��@�M�I)aB�}֩���	��X�ܽ8�~�@�(�7�=��"Әm�I܉����y��j̄�T7�N[c�ۮW:�D��;^&�C!���`)�\&�H�G&�f$;й�'�?}�����J�>�6�!�Xd�'Rkg��ӟ�wi�$X�r�:��Wc�����|����k�Ɣ���H�/��B��*d�}tx7�F'�V_/�ٓ�v�J�׉��Xб6\e41�5����毂�Y�MeD�\M��/Ȓ����g����H1>�|���R��+(��Z��X��z6 ߹�)&�1V��z��	+ �x�����gK����j�4M�� �V�����f#�b-cכ:c/����?"��9�nG�q����`���X� ��UF ����j�1�aU��CJh��R������ή^sG^�|�jO\��)��,�rC�&�Z�+T�s��b���Ƽ �?4�s���A�����n��Ջ?��u�q{���z��G�%~e�d~b��N�ʬ�|�W�Ƽ��k���Wͪ=<��Q�$~K�k�~
s�3��h9	$�D�������B�D���-)�8����[Wt�l�
;�Ǭ��D��<hQ�ҬQCI+�����GVy&[�ʏ�W����!��7���|�;|.H��|���S�9�)0�(W�
"��6>+K�A�G�+�
���1�y6>�M��?Ѭ��|�P�p����55^2�Nn_�߷[1��;�#}��ܽ{W�����>s2�6��:���G2 ��wv!7���֓�S�e�����K��<�/?�G)_h�Խ��\��|���%!h{��w��ӱ9f�^,RE�=�J;�	C6�|����?�}����C�?���L�<�|!�Uf��Ƶ&�(�n4>�m�D��&�%;�m۶m�~ۖ ٶm۶m۶_s[�� �tʃ
$��^�,�#��"�0�a>�<fKӷ��yc�%��B6ff`��6r@�!k���I��Ad$3Hfn�Cdwp�şU��Ä}w�#�����7�+H=!�@)���x��G
��пi�-=���=fͮRO�lc���W�� sxrG�N,ӱݑ^�%���d1Sט�5��{��z/��B�/ ����q$d���x_���+���'#��!�D���5�0�ϖ
'Q����8N�*O��C�Ѓ��;��y<$� ��@��� }CM�p>���À��l���h"3�O4�5�-(����+/0���hG2�ՙ��%��g:�*hUO��zd�RrP���ܻ�W[�&#�&0T��*c��H��NA���RN�����ruuC����PN�=��?|�מ�V̠��I�uJ���D���}9�ݗ'���7���h,i�ү�U��'�0��lR�� "�:����������+�x�3��y�?aप@4�ҁ�)@�Mִ��fÖ�	Bм��C��D�/Ty8���d	P߁9�S�[��,���l ��2���z|�S�|C����R�_���tA�H�`�!���2�	��X�����g���+�LZ�)����Tm�à�Te$	�sh��]���oݗ�����Ç:��A��9l����0�a+ȱ0tU6i1t��A�t���#@(QV8	4���A%��%���2���M	�, p �� ��j:9�E)W�3λ���hL�Z}�ރ1i�t���ġΏ���Mg9N(75�do?�Z�<��zM��K��Dd��<9�aYYAǪ�r��T29������A?��4v����7��r1	�5�X=����|uAҴ:�x]� +4�_��煍D7i�S����I�\l�8�׵2_��,�e��1��$C��?'r=1/$��?z-���r��|�+aܓ�P�C�.�X�k5���؄�Ƞf�גt����"��k�?XI�����B�}��ܑ>b�.��X������È�� ���Az�$'+#S9V+#_<}�UnHNBI(�ߔ��t�!�9�'#��ȚTeJ�E���#��tm�5ėGߐ���Sd]|Pa��3s���d3/��	����0t�M�J�\-hH�m��ܭ�d�볺��x�U��gZ���/�.��Y��0��������tHc�V��I���s��I�7�y�8X�@�*�6TJ5�\��&�d܈��Y���5��c�`��
<iiA�k8�a�FU���9�,���΁�;ݰ�>Gm���b)�̣w=�������\�Η���3�k<�E%���j���r.�^������{$ l�X��xY�9[���8��[��DL���5 ����4�ֽb{�FEF�k"c�vRKS�W$@V+��Y��3	r�X߱A|��U�B�H೒0$�Q'�G	-}�I�9	�"#���"ʞu�wMzX�s�E�Hb8l��Ű+������w?�o�NX��mȢY)b����C�~`<����q����>-�K�h��hE1�H�<��YW}�i~��K)�3ܥ���J���/|��r{�N�KT#��g<G��rq��=Tn�lm���H�c9>>�5��I!?�r(_}�9�AH���,t�=Zj��=kW��ɝ#y��=ݟN��7���j�*b]��,��o�%�{��'ߡ����,Qa�\�Z��/���H�L�.���j��I�	�q��V)*lt |��gr��+//.e۶m۶m�~;ږ ٶm۶m۶_k��Ź��V8�eH�,� ��5e�F";�T=�EaGVZ�4��s)4���c&1�~!��U��0lD���y(jX�$��,�(KFi����  mR5���` ����pW�;=��j-�7�`A� $f�:��\V4�63�N���mF�(�_gK=��T��,�E�������#��w?�[IKf��\�(�4���� c~�N��!<P �ǱO���VHL�od�� 0rQ�1��LH��&A?�4�D��즚&v��8��!1�LZ���){`��F$ t�H�,����� �T�� M � +�z\^�[da>�e������ky���H� �V2�Fz�5]��s�[X.'���c�7-f~0*"�C��3? ��ұPD ��$���aN9hL�P�d<<�d��5ZY�'�d���l�Bj�H��%ط,TT�܌oHnAb�j.����-�QV����2�{��S_��M�F��A"C6z�4=�yM�~�C��&����A�5�փ���1�vؐ�X�v�L��[��QY��W�X���y���
�p�?�ٔs�P�.9o�I����Z��t���gdwC���Pj?k�i�1��+�/�2�\U��#J�0�d�9�\G�A7���a ���W:�c���#?�s*?�����Ӌ'���n���i�Y�j1H�0� �eқ��/�A�o����{�3u8#�l�M����W'�L��5�UNxӔ���2�)��2�r����C�&�R�CIXߑ��F�Ʌ^k"�{���� ��@�\+�k�5�TK �@X�R�F��4�3�U��B��7�a`|�L\/2�ר.�n�����2�F[V�$�ڸ2���� 4�о��l���������L�/2��1C��>��WR�i8��1�H?w-k���3���<k�Ȋ%�J���OCBy,�e�r��f$_�#����w���;=�Z_c�
��_�1^&����F�� ����!�i)/3�x]�b$��~��J$~q�Ϯ)G�wdp�+^�P�r%��>�Z&�5?�A;�k�^%���d��d#�Z�?��W̤�����p��E_�q�ҵя���*�<��k\�ϟ�%lN9�
��5��rd��!���宪�s �Y�2F�4�.�m^�dـ��6���B��� .������׽��ï����^K�J����8������=����Z�x��c�^���1�n>�g �c-�yxi�J��R�T��@h�]:�$��X����B�M�Yd	��zT�N7�5G� ��|e~^YN�x����q;�&�(r[�ϲ���z\��kל�hk�S���p>�\&ӑ<���Ŭ,�dh�S�p�R���L��w>T�-���XZ�c*�/���v�����Y�x��x�=��{1#r�|�*�� ��d*:���y�¿����#���лF�8����X@�+�������'.�����A��q���1HT�>+W`��l6X��h�$]r�e�+�����º���\�_�����Ϫ�겪c)[.$�g��5�^������txp$����w��<"��Ǹ���*�Ģ���e�
c�,��~�ejm]
%����u��u�<v�'�0\��?�,Y�y&��X^�z���3��[$,����g&��X	��p�z����|��'rtx±���U�Ϯt����ø��YE�*aO�%�Y,��"�S}�c�����.���we۶m۶m�~;ږ ٶm۶m۶v�s�t]�"YK��I��@<h���q�4`S� ������z�mv[�\MLW_�ܛ'+ daD���� �5�s |VX �
�5�������V6L�a��.SY�2fi�:]4�UF9��Gz0���V�E��� zVt��)u�{\�W2�ٓ?��?�4Y�P��?���s�*����@C�ߓ�''N�i%���i7e0�74Xquu-O�<&H�zp��$[M�z�vbi5۔��]�'*�Es���4Ku���4.�C�~�)3+��.�ȃ@
�X  ��o��������C����e��g4��Y����7�x��2?C=4�����ɒ��s����?Py���wߦTY�ݑn���+�פF���dN��L�+������C����(ö3�c�(L~=z,�?���50��谯����et=�d���ND�"�x�}V7�72���o��OS��{,b�6�R��K���Cfq��G����:~�lJb��R׹Q�t}�'H,\���cf��[��|As���J���x���TH�������MҿUR:�� T ��x�Ƞ��:����_�~͌jx�\^^�h2����uO�#��$I�ԹM��T��:�aV[PxF��-ك*#TQ���1��q-T��>[_V�I� y����e��4Ao�=c����$�XC_�Ծ
A0� ��N��8�X-lJ���*63[d��||��R�}�,Z�����ɨ���D�f�}!���F�}�s��d9�} �-�M&#��s���?ۑ�5�>��k��4��=�lM��{z�+C0-?8�x��-��(�_�H̗��	�j3������N�6��m��<�uv颡��_i�,�pBb$��.��\_��C_�=&�͈� *��8!����X���T��Y�?�ȳ�"�~���#��B����K�������#�?����x�T"&��GR��h�c����b��Y�j�D�_���㆐x=����+���Wѿ������|9�2Q�ƃ���A�ƶ�,��8�W�3�\k�5F7�|��Sy��|u$�?��w��JC�o�N%�tlzs�Ս"�Wήɪ?`P=I�£�ӱ�Y�]�h�n�>�|�e����ܹ��P�:�����D�)��HX�?^?.�ƻR���1�:��5>�"��+x+�Mf��i[|iU�����tX�C�K�4�A7A�,5�^���?�L��/�B^�<��#J��r�o���ޡܽsJ�"�9��5��
	��A�rE7�K�G+VQ�l��uV �F%�~��o�K܌�C� h�!~޷d�,�P��l|z�8�D����w�Z[E��Y�����Bf�V���qzr=b��	�ób�{��4����\#K^|�ν~&��6�ZX?�!��n�'��)q9����m��C�����)�Y��Rs �S�	���T�JBf
Dث�5��׈�����~b#�2	1�>����9��Q׸���LI��Y�
�+���UP�Qf2�5kM��&�d�C��t�P�U3 �Q�@�-DV����ɩ	�5&
MҒ�Z�<q-���ai�|k�["
��#r�&�A�׆�/T�!A�$�grO�T�_�l�V�!F���c�k�c����p�ƺ�:8ܗ�?�P>�����ѡ�{�T2��ղ���r��a��3�o4c�u�{&u�{�U�a��ԡ��DMT ���������?;�w���Lu��t�9�}�R��_��{�S������{���:���`u/?TBc���[o�/}� v�����Cy���)���'�ȯ3����}ݿ�5��Y%�p$�{;2�������ӿ�{��~Wޤjl۶m۶m�oj� ۶m۶m��ϮE����,��04�������fۅ��΢�5 
Ȓ��,A�4F#R�����zp��]:]���1�r�� N�ݽ+�'���:20�Ʉr���rV�PFa���|�׷ ��"��C$�VJ9�b����l�!��j�!�I �w(͸�{ov��z��?�����Pe�F_R���˧2�C�*��s�j3_�2�yrz�}e�����E7�i
��ȝNz�[f"=L :�s��53؛�5�����MG��#��P��K���������d� ��
��� ���"�V�b/����d�a�~�AV�j}�{�;$E@� ���>?����ط1QJ�Њ ��=�q� 8�x��l~3���+=�-/^��u��U���ٚ��gOe�������N�g2��Ո����9�/7���y��\\^�$Ma���k���0d�� �X�`Ʃ0�D���6I���a��U:�Ha��}�޺���%,�&���^!�
�� �}S��)�u�N�j��`��s��Uh$A\�?��F��I�J�f&���g2Q�C���& '�ь��nViz�Ŋ�i�'%�o<:�bș`��ry�:�H��s#� ����� �o]�	�n��sï$M�#��J�G7:r��z/%?���\n�U@�HH
��������E1��"���L<����x�#���D�I�!�~�Y���U&4�Ƹo�]�/�L߳�
�˳����I,���X$2~�RzUS�;{r���	ڧ7 '
������AV�8���YB����k�YK�n�s)��g@q�%E��@��\%�U֞�?J;�����'��$��<�M�7��|��� jS0�R���⾟�y�L�'O'9{]��-O�{��C�
����X��3�{m���R�4�O˚�3K�F��j|�C�je�3ϟ��dͺ������x;���R\B���Y٩\h_m6b؃���8/��p���B��lR�B�ȠV'��cW2y~c�҆�sX阫�r��2��'F�8z��o��T��z��#j�x���OP�83�΀�3<�#�_�s*u]�P�����y-%���ִ����"חWRk������h�G�-����3V���Vٻ�f�c����$V#Թ�1 �i7����7��_����G+?��&�O��@��<�>���90gfn�s������^��;�x�j;��s�	�a��#ģ[���oY��G��}[G��Fװ�U� )C ��U��O���B�?�\@uDN٤�I1�,�g�+	����	�dki��{mi��fV��d����ڳY�	t�?�HMx��L�=5��VV�"�Dq@R��i�} �m�P�AFQ��|zO�"�D5@%��Ñ��kT`��������B����Vc �F�	�XP�	��>`��*6�۵�����9�a����ƛ>�Pf,t�<U� p���n�&qI��Ī�@� �%�߉ybDQEI%�"�ܸf$�]�(�RF�#��	�	c��D�D#�q�Jaq?[���=Or[���Y���@{�����z��+�����{�'�}������{��υ���Q�Sʪ�1��d���Ez���J��s�G�s�m����1��*�اC����|�{�cm-_}�S��}��z�`�h�����i������^�X���)��	����M7�ŗ�ˏ��Sy��!:@?�M�w�UP!u�c��ր���������٫s����;���#ٶm۶m۶��%@�m۶m۶�U�tLog ��>���X��r��.�c�l�a@N� S����X��%� e/Qi@� �����e�Yc��9������z~���f�m�L	n��N h��a��<уt�"8��˥ӑ����a<�CXUdN[zMp�����ށtC���^螣J�����ߖ?��#�^����HƋ��x,j�w��d��}qV���F���K�\@T�q�$�''rt|*g��2��H#0n�eP:`Z�6uu+�Lv_B��ii����f}0�~id�t�-�+2Fs�@"=a���� ?�����%2�A���4(`��j�$�~�IJ8�	��`e��t�&C���O��{����p �AO��H`A*  $�]�A�{�]�oP�Mf(ݙ���w�����`&�lK�:ͧrqq)gg��R�{���<y�_�����<��)Id�滹�J3 �Ϥ���!]'2�1�']DH�@�f��_�L�ק���_@�0�thy�P�TB��[	+�f�		�ɕ���8�X�B��������UV����ٹm�o�z���xӨ���&��0�]@� ? i�9�{�PIU@��^?�����r}3"��`�wA�g�d����q�h8��dN�$[��+��f�s��M~��H��y��iG��G1�q�"(�N�8_WYa �n�@��]���]�����RJÙqr��}�B�JfsV�+�ƹ��E��P����>��wh4�*��\H]��Y���� {G���g��k��Y-σ�"���H�?��/�h�	�xT��ˈ	@�d*�@�����*���e�맬V,�q)O�$��uc��ל�_BOQ�/t�m���R&<#�]�1*�kh��{Ж~�1 ��G.^��lYr��@YC�$n�Bf�X�~�5������΃���H����FxN��L.��g�����;9�%���(�g��
(���R���Ls��\��yz=3�Ld>�k�V]�M�3aC�>8��R'��'Դ��IG��C�~�n��ߕv	���G0��8e@�z�r����>���tW�F){�SƘ�>�Z��k99��NC���;\�KVϢci���$a��'���SV7]\\h_�C���>H2`��9�+�H���>����?>��w�Sk��8`��$�F���_oե�5C�L8 ��a2�:�����t(Gy��k<�u��������������Uq�є�P��VS?3�s�w�-[#��tU��I16u�	5��3�!�������V�Hi)�(�F�~��b#�V(��&��A�� ���d�P��y�EBɦJ�<?� c�����y�`.*�2�c��t�s��FW�P�þ���98�J���q�>�7 rp�ﳳ3�p��{;���I�KSP�k�Z��Ї%0)EV���tt,�D���Vs� i��ق����1]n��('H9M�����7so=�ĪQQ���r~vi�+�&=ָf��&�A���	�蔎+H���ʰ,�ס�J��f]�,#�d Ʀ����I����rq���
HĀ�)����=<I�諸L3�!�߸*��D���D�Kͼ@�x 2� ���Vr���`�8o�'�:�X��	�	x/�4
�L�$�~(����d���=�/o%�l�g�i�=`/�>��*�?@@�9-@��"(���+��C�NQx�ܩ���t9�=v�w���s�ǟ}���=g��g^�>����9�ݓw����+�q}��ހ�1�E�:�ˌ����L~�w�����_���������{���/�r�Пm:I�h�=��o$S���ޫ!�:7���@��_}_�m۶m۶�7�m	�m۶m۶m��6$}�� %A~��<�݌�f*q�+~I�7���a�C�ْ�_�O�t�MG^H�� �ɷr�;{҇���X�w�ꏨ#������ KsU=,�ɝ��j�7M�Í�mz���^=,�\f82�p��l�7�*~��<���=N&s���K�S:CΘ��88��ʃ�ޖ���!=���G�� 2�_���.5d�x=��L�'��'  0���},�z��s"~���Q�*)� ɟM�~v�I_X�z)NncM�V�5�p0������PR@i�&�e��nޣJ ��;�=�ӳ������y���8�#c��rf�C�"+M����<Ki�bfv�-���'KG�4(a��T-��s�e������ jw�ՆTXD�$�fB��8���B�&�0����O	���y���|�ӟɫ��%j�X�1��4������'���/i����H��I�ݶ���l����u�lbFrH�R�o����b>c��ׯ(�>�8���x<%(�ß��H ������#�p- tH�@�v��s����}��fB"�$@�u	`��wf�W��=��`�2�y����Z���R&�OT]�X��g2��E��v�R @$m::�Z46�H� ��;$(��l������ �0�{}^��ղ��o����^���TW怞�]�kɌsd�#\��/�����PM`�h&�aL��ţ	��O{rz���ypO@ 4�׉�ˉ���G^H
LR��ޑ��c����j�n4%l�$�XY$�K������ �*	�r|򖜼��Ls_}���<��/��g>�zGGsW��]�ؖ%�W�D���H��q!	+,
Z3������5���yB�*�9�`9�[��|$�>2�#�{ �Wڍ7��2I�2Տ������r����1���}�w�e�p5h�K�פ�,������:�W�
h��"�a_vOHsp��wW�M!�^<�����g/���@��Gߕ=�O�t�,/E��% S��QF�0����[]3���zR��9��O���͵����rt�Dױ@�%��!P�k]���O�? ����i��jJ�m	��<��^S��\׌T^&��·;����1X$]O���Ȱ/P-�h�ן�SH1��k��i�u�h��hL�	�=���%�����vt���"4~�ndU��Y�{�]�־�����D~����L�}�ϵ�!��e��IF@���H8��/��5����A$,`�����0�Yu��?��\��	��� !I)E[u�ϐ� ���xI�x$)Az���Z%$�e���!iP��*�+X�5�p�9@<!�\\��o��*t�/+��Cr�[l�+23wGE�~��A�WY�Y�$�D�.��o�򗳕�+H��e��e_�2Ǉ��s��^�f�h���*]WP	3�O$Ӊy��������8w�13���zt��d{��~X��PG?��n����Ʋ��j�rҨ0B��PN� �8���p����Lp�#Q�_cuy� �Bl6��.��D�
e	��%(@2,1�U�9K�R�mEE�!b1��pE.рK���&��� �����;]~�*�X�o�n��d����Jޚ�=���g?�z��U�XKA��U����� ����TSb����|��:�����e�X�EY��s/�	)DHjj���N����Sy�Ïd����Sc獵�>�X�"z��ܻ����>�����V&٦���y�ﱦJ�b�HP��+BKڀG�L�i��VW>�}'�9���J�����L�e.��g�c�a�������>�N`L����:�^��ttm<�7�&2��4���O]�R]�P�����b� �|�%��^��g�Ϳ�޶m۶m۶��%@�m۶m۶����_Nn���ʋ�>b��o�-�~���!u�❾4;mJ=y�L�ZC�o��@H?)3Qy�*�K��C[�%o�����!,_���|���> �H����,	�FzD���%9��l|[�O$]3�r� ⁷���I������|1nn"��l4p�fv!gm=�����~������O�����^M��W��uZ�%��u7��`v�fֆk4�e��a�?m��4>q� fb���꒩3#"C����s�Q�0 �F"+3#��?��s�9M����ï>�o��-A�1ɓ�\������y���τ'�"]����#��/~��>_UN��H �&�o D�^D9�h��t%j�Z��;0,�xKj4N�(�0c���2� }v6Sbȣ)}���e���~�O�/�D�f��%e6�� ��Z�s���	R���0��a{�l�gE,���-�^+�\�V�ua�hcJ��/C�����z�9	�ax�PLH � �h4���~�����sik��~ss��8%�3���ޞQ���������ٖ��;�ί�}܎,KH��o2<��A�'+���}A�)
iz�2�E�-@��]wD^B3�߿d_��no��!�2F�z �Q8(�F\9��xS�iMt�����䏊����� "����2�������<Kd6�QƢ٨K��E���)��$@�l-�5s�@�t�V�Z�A��q�AC�� �G�W|�O��wd�T��H�dݎ�ݖ��q%���[���a�T�R*&�p^�����U�Q�>�2����dn��)�bC���DL��)Ko���y�P'�])�L|� ���B���O���>���=���T����w���cY�����`Z�G�uPUڻ�{tG��'������@��\�}�\N�|+����;:�=���������]���Τ�ѹ�1��P�f����5�ï�޹+��m��g��@����}�����}�@v��������R��cuQѮRH�sj{_�ܓj�&ק:�h�׏�9�� r��%���hj���I/%������=�������j���[�9~��ӕ�h�m���K��[���ԛ����r�&����d��R��H�@��O(�f�n���g�ڗ�:׏��Ù�?�������щ���Dʭx�V�|*���>#���ZW:gH,���`��mHS��ѭKk{&����:������߬�0�v�씇�r)�|"��Lf7�2�qTk�u(�YDr3\�Md��p6��z�V��ՙ��J,a'����#��T�h;>�L_;/�r5�y]'��(��g2_N�Ά�^7�  p2����� E��eDa�F&�Hx�z�Q∺��7���_-�$�_$�$��՜�9Q�cK�R�吝\�%}�t~H&~Q��:SH�s�h4dvDK��G�y:Pv	}P�%L��\Z����s�f����е!��>�
fMi�@?#A�т1���~����Ti�3���<�9��=ɾ��nK�ݤ_
�À&A��*Fݍz$;�.	
�w��>��@��7���p�G�g��G_,�'a�����������D&
�3()Z����4���
2ː�����lm����D�e�%����C9;;�;w����/����$�%l*�q'�_��o�Qa{.���Z?��Y�a �D�N <��6�F#HAA/q$M����3��B�!��ٷg$���X�ZOL�IL:���C"����L$�kX�����ȴ�f%I"����|m���pg�J��-��;9�a��qݨp�}�����{��ldC��?��&����_�t��Qk��&��*x�uu>�`#4���n�d3<����)�����像>�=͕���\�p��E����Zvwu�ۑ����M{ӿ%т d#�?'̲�3�ׄ
2a3�����c)����X��=wB���*��Ȩ� ٔMٔMٔ���!@6eS6eS6�O^z�=� ���K�9:ޓ������}��$���ٷ�ӓ�;�d:�嫯���}���N&G���0����wߗ��ωӥ4~�9�C��	�֛��'P)��Ar|�X�޽KP���.�ߍ�H�tY���+���E�Sݫ��|�ɀ/�YVJ��ЏC("7�)�aJr"����T59��?�P���;���S#�K����F�d2��ˊ����UF�!��ѱ��d�l��QCĮ��*Rue��{XI�g.	�d%k�C5�Ղu�ϧ��\�ri���/6�V=�w�-~�\�����j=$���4��\ٿ��0҃z����VG��#`	6��ߌ�,�Ɯ"���m�S����)�"N�#gA�J��-��#�V˄��@���g/�9oGʖ�\�ҿ@�鰢���ӹ\�5n�C�`��n��^g�&ؗzÐ}�S<1Y&x��ky6H,��E��0E��՗�w��Z��$�n��� z�ƱX�ɜG��O�/�k@����C���'���4A<��4�L��@c��_`f,Kf� �c��1�N<f� KB���Va-����R}uO
E�� x�E�9k��{}ϐ,Ѻ���>#"�qO�cC�`<U�֩����Ǳ2��7��4{ԏ��KE�!�i��������H�]��BO�bCȣ���ړȯ�<K5��}(H�������D�ԛ�R��A׼��ݖ��=�ɎLu��w~�2���k�ʩ6A�ˑה���H�����A���Sy��+�����y���ֻ0	���H&�^*��T���?��/%+�d�����BYS�e�4v����"Uw���	Lϵ��mm�=�4�RߓK�^ŗ�VK��^����s��nd0�[��d�k�f})SH�r��m2[$hi����r ����<lU�o�et���Bd�\�ֻ�4���!�'�|��wrz>��ȣ��FZ���2�K:�$f2�I%� �"�L۫�M(u����b ~�L�b����+k�jW�m�t~;���S):7&��3m��>�����@�e���H���ʓ+Y�_��d�}r.��n�?��Lo���q){ !͓�kJ����ղ!�b[�:��/g�y���X�/�������N���wz�c!���s\g,�����������T��3�k�$ש��+��M!�������/er}E��j�E�{1It��XK�悤`�]&$Q1Gb~��Q� 1F� �y0��2���-AS��!L�A�Tm�Z�SX�0���(
˨�} Yc EF�7�X&[plh�kc`�\)�aM�f%�U�\{0��.`�i�/-� 4d{�	�\�g`]���:$��Ga�#g�u
9�iJ�"5ţ:���@`��t;M�`J���^*Q��7�n"J+		�,�3C"ҵ�C��b.�fU�����=I�L�#9y�\�єu����ϋ3�7jm�*���tb�_��U��b�@"�Xg��3(��XV(��j������a�v�ڀ�� �!͆��ߧ��d<r��L �4�x�=�td��ɺg�iIKKSe0�>c�%[ ����7W�lU��^�x�����nG���^�2A�`�)�o�y"�����Ԥ]�$H���/��&u�I�2�B�'�!�g^*(�GA����1G�3��SAn�G`�$��} ?P�����`��|�{�0�g2�?{2�Ė��" ���u�$��@T�أ����!}U$l ��d�f����Z���U�l6�97�<m�YU ��{���K�o?�"s������Ҙ���>I��m9�v�L�TPQ���\�J��amе��n���t~(F#��- &BFYP����>�`
�+P��۳�����?�Z�)��)��)�eC�lʦlʦlʟ�<�˫g������#Jp��������O>��;wI~Ĉ����ӳK2;�-��O	 O�"�U����A����w���w��թlooI��ԛ5�%�z Y�pfk�'�=҃�!���f>�"�/������^� �u��i�X�"H�A$7��S/���ƙF!7RP����-�c=���]	#fZ�����'���\^��)*������K-�N�g���X��/��ҪUe03����@3�4��s��Ӳn#�C��m���+H �b��H��Q"�,L.B��q����^Q� �"���q�uTH�۔��4�F�[� $ �#�y���׸�H)> g�NGr��&� ���C3<H��$����eI�XD��Lg�$<�`Q����R���Rb�㐾"U�!��m���cʳ��W�˓�ߚ1<��=�d�
��dy�\�7}ɴ� š�@Z��h�יAj]�KG����Lw�[P2�rkF��Fod] ���8҂�NG�39����( ��%@��/ڶ�ù����y�o�VY:V(/��6�]��dbD1xs�!3A��Xd�V2�4pֱ�[�Iy<�g�#z&� 4�&[�Gp6���φ,&��4�E�QA#V�����e�\�Z	�m^����O��0���F�if2p��A�+�%�`�\}�z�nc}%2�#���Aa�A����l��Rolk�h;�e4)%��u�����m�V���[ (�-�A�ĳִZ��<�9��@�<H��Y�I��Q9�7�=����T��������+y0�e-�$�����\���U���Oe��߈4ZR`��8_�mC8K�$@�^!�@�S_N/�d��k�lk=V�t���al�&M�U��H��H�@�/���F� �푡����2������7_\�g�e��q#[�D�.�2]��<�`~��x�@�O��V�ond��~2���X�̏;Lt����c�N��{�i�z2�O��ō�l:_�$R,�u���rsu��{+�|DߚB�{t�� �gѾ;�e���gW3i��Pr���V�KÇh�K�BD�G��2��� w}`9ϧ��A�v,c�ni5�of�����^�Q�i�s#��H�~{*'���8i
���~�0��b�9^�1��G;F�ΥҾ�yףǖTsi��R�'��`L�j㕤�6�`17�dj}F�\���d:�/���z����8�IR,$��2�慍qx�)���X���˜��WP�ÜCQ%�ڗ�ɍ�u����O� n"`tHi��2���,�l�C�B�񸷻%{����M'�NB�Y��"\� NH��-+�޹G�3�b�����;�2bk��3�e�uu�i��)=3z@�W�	�y0q�F�Z�H��"��L�j��t����=[�j@�1dC,�	3�\�,|�9Kbfk��m�V��_�Z�O�:��l~d38Hx������(�}J��t�������7k3Qw��4�Ƃ�$D#�K���5�'��ql���;�{�DC�^<_�hWP��	<3lª�7f�^�}3��J'5�0)׹DRu��v�|A ��	�ǡ����I�t�N��f���e�2�k@�\_]�`�D�۲X?�R1�9+��`0�A&@�^7=�<m�֙�'3F����߬�j_ �A��&_����������:�7dv}�sZ��]	I@�ݩ�A*!0"p���z�u_`?��� �#�P�T�rh���y�y�t+J��I(�Ԗ�۷;98>�����]�헜��.�F:�UH�n1���=7ƚ+�y��������Y�/���7�7Ӿ0B�%����b�=~Y2[��i�-����)��)���U6Ȧlʦlʦ�i�~�1 �����w����޹C�摐����7���k�j(}��|�����[��/>����D������o�� @؁���Ő�	�� I��ݒ�cF�� �c%_��
�n�;��5c�j���4�-���ڌxDV2<de��Õ�D�{(
�C!�$��Vi�|��zo�ן��$ h���/e���A�&��|W��`�zpM���B���K^ݐ ��o����3I1��f�U,
�ZI�@ɖfnJ%2���I�H5�`�5��7B��U�kQ*�{ �B��@nnn�`@�`E����&��~k�o#ND�-|f��0���)�%�>���B�xA��0��%0|3I���1y
٭�|_Y c�X{�x�ID���/y^c}K�A�F�-��(���z��#�{b`�`ȃ<Mm'cI�KJ0A���u�# f����j���rxzJ���T�� �#{��DF5��C$.}?\6�;��'�3o�~ 9�Q�.zR,R��c��k��h�a8Z�. L���H6$2fY�/���f��}1�z��C\3����j3��y�e:&*KA�.�f��@�>�*���!Ř��.9E�I��&Lz��xZ' �?�v?�4 ��^���5]��8��!��(��%�ɮ�u F!]K�}-��VH>-�_o��v�6��qn�q�ٽ���,0@����dI��n��lIt�f2��/�d��?G��!����@��B��u Vf�-�|�t ���K_�ڇjr�T��~��P�Ӆr�~M*�@�H^����Tǐ��(K�����������/�:��������X�;2_h�:�s�1�Gn}J���/EE,��D�9�չ@�{8��b�J�&��D^T�}K�y:����F�_\��gS��`�c!?��� �8�O��݅.ڧ�}��g�!������iꜽH'�UR�������.�ǲ��H�ty�_S��Y"2Z2X4��7����g����R��J:~Ƴ�rv1�z��q� �����l~Q�Mdr�ʫ��I��5������9�j��w:(�{��RX�W`Nr$hj0�T�Ծk��&���a�lĥ������!��0Vq/�aO6� ��b��F�L��%���3Ԙ��-Ț��-���u>�Ų�	����Np>Z"�&��Tm���Ί�������gs��H�)�rPL\��R�e�4NPǸo2{ ��" V҄|f�&:�§@2�1P�R'|ǜ��C��4$��L�(͜D%�f�w\���c����K��<�������Z�Δ�%�d��!���G(=[��mV�,B�k5Ao�'���\�{A�kg<�0��u�zwk�y^�+�kAuuZ-���RR�y�/g>����;�>k�5��ǯ���h�����ݣ4�2���G&����������S�}�G� ����s]�<�:XV)�@��Rb�Ș\�mVWm���u��n�6�w{' �����o2� kM�i�0��w|>��;Ͷ��&G����q/^�P��R�E��iS�@@�T��P��X&ڮ ���m��=��2�����d��k#d�&��K�����wlKt�mq��qV����u���+ُ�<�����RL�A��|�=a����72@@��n_W��#B,�ڇ��C��ܻ�4}{Bt�SXg�F�tOBb	�oN*��uE�2}&<?��̈rR�����s0���{�9���A�/Td�	��E�s��-9��@��ݗgϿ���6H��j;u�T�=t����w�2S�ˇ�C��";{��ÿ�w��?��72���<��y�����������ޑ����}���������e}�z���ٔMٔMٔ��!@6eS6eS6�OZ���3Ro�c�lo��{���'=�@>;}I��	6 + ���|����ۏޕw�y�l��?���+J��^����S����i"�����3
R�;���C����h�p�ߔ���-)_��|H�X���!��+��<|��������t¨Pe��7��	�A��D����\�x&77��'��]����^������������s �7}yk�V�C�,h��z��v:<�����'��fx+��X�S�+ �����Nh�@`�!p(��C���x��!!��z���O�23���,�:��A��m��C���/�*A� ��8�O&s�S#J�����h��jN�jD�;�zHG��`��Q��cE�>	� �сz�w���e;(!��j�Zj� ���O�!�5Nc�+ߐ�@��<�Rv�v�ײ�3m�}i��~�L��&�y�Q([��m�����;ȱN�!����m��zD��y�˫�km�5�Q@� @>H�#J�%�*��A��qȂ DTe�l��`@�
 �5x�4�A���/c���)u�:������@N a6�Ƕ�7$��L����zIX�#�7�z�IEU3 옥21�O��� `V���f�Z��H����>�SF_g� �c6I�a���Z_��{!�ԁ����J�DL�݀(B�-��b0��H_�<��I2Kd8�9n	I�D��H¼\��D�� ����C���֭���l���ń�"�o������X�|j�O��L�����~���Ӷlu�m������?���@Ʒ�GC�\�V�+F�O�c�N���;ڧs�\��ɩ��X��X��z������l*�v��;��q������;yz>�2��_'�#��,ks�H ��\���`.S��H��k$���4~{.�V�YM7�3���v<�I�q��?rͨ��,;���dL�@�_j�.�������J��B^��Ҩf�Ƿ�$v��e4�u�k�o�����Onk��B��!�YBkQ0��ˉ~V.iK��\� ��p��i�xf�n��
�#z����wY }�w���ݼ�,¹��Z��S�~\�ˊ ��1[���;��Q��\�Xs=Y�r�$�,�s�۳��:�x檶�@z+��ߠ�#8=K3	�A��L9�HPa���*!����~�z��`O9yq"��Ab������P����ar�;^�K.9(��n5���%��0�����j�a�ؐ+�W�����Qj�H�2�ꕐ�=�p�� 	��4��h����'̦�_H���Ø!�@�bs��հb�\-b�����^+.d$"S��3ϐ������yb}j5+a����������/�V]�U��Kf����4����"�x~K�f>)�T':������}�)U�uzp��p$;�]��y�4A�	I	+�ld�z���� ��:����!%��ũe+`O�/$�e$jx��!}�(�DrzN2&ֵJ�� сz�4�xd>"X;��� �A�h[�Y(����l�d4�ߤ{���P��V���
t�':o�@�}�����յ�u����K�H��9⾥��2>#I �����$:�����dI踆w�u>ֽhwg�rPأTtmC�(�d6��s~�zźN�y�"((]�|�ڍ	Hz�`�ѽk$�N*�^���
������Pv�r=c݃Nu�7��תWI��s�yQ�{]��~�q�&�N�{�(��3Թ')�}��x��*#�k�u������_f s�C ����f�/CnTiʎ�����2�~�R���!֩�/_�:�/��]�ӽ���@.ϯd<����lQ^���w��?��<|��r��[���P� G���k�{S��>�sš���J~��_�?��?l��7eS6eS��ʆ ٔMٔMٔ?}Y�� ��Bvw��i�
O x)<}�L�������sF��B��������������Zz�����i��,�!@�r���r0ɬF�t�t���*I�c�0Qo�8f�<@��\�����h��r��y�V��g��x���0d�g�0��34�4:M>u[m�:AZR���f�kLу��������ݽ����ό&���V�#�Z��+"�0s�*�GÑ$�%%T*�J�sZx�Ѐ����h�] 5+WRKvZaĈe�v�6��t�qP�a4�'�f�vs��kuY����c�l��䆔T������;�5|��d� "i!%sڊE�#[����}F��墙��އ�y��6�����^u䴥�	Rp凁�r1y0�1E�%m�h��r~~������9���l�Ç�	b�xqB�1��Gw��o��g��|��S��[}��������7�ć�PNB�]�R!���CR�
��ݭQ�.�>GけW��!<�:|��Z�#*��/M7�
�̙�J�f��zNҙ^�j�V�G����eMt��b�z���{�_$79�0���ŜM�,aN��!b<���N�f���&b7���DHZ���B��
�0(!A���䭂�H�he.�z8� z  !{���� ��<�+��e+�#��1�>ZD��K����~�	-v�q)*���2��%�ܤ��@�,�h�To��H�E-�~Qx���\��x�V_|�Rj�ki�:��|��w3gf��bd�1��%�s�� �>��A�u��?�g{B�	���E�C�c(��L��0o�x�|��u���4��4e$��J�-̌(9�~�6�`h	��G݆:?�)_L!�b��u>�������N�hӔEn�-En�x��k�Ϗ����AfQi���23���{�
��(K��	��3J�H��Y�T�ֹ�8cTs�<tr�6j�̅�Y���7@�@5da��~�}}��~A> f?m&�zO˂�T��WP
�dg�1U��H�uSx�������	>���w3���W�b	�����������될-�*�8������-K�Ԏ
O'�+S����^�z�a�`��rG{,&���;��湔�P,ۆY	���y:AF��X2�ټ����  �Ȁ��1��H��X��6�@db}������J�dlb-�7�.#��|�⤋ }:�p���4[�K����"� �������m:ק�k^��%������$�*���@06u?R����k�o)҄Y�p��,5=�bnf���cF(�!�7��'ؓVgK�z�XC�� �ͫ�d��0�A�IO�lmS�w���壎��8α��	�4�A�!��E��~��&}�>;a�P�P�#�'�E���^s�s�I��п�Sf��saĂH�V|f��'1��S������������(��t�5fF�2��dr��Zw''r��qY+�̡�~�=�>+�^���`���[��ٯx���yO>��cf�D0P������LNt�&�N��Y� �!]V��k�zo,�������2d/�[��5�v��~���@�-=�0�1�"���`8`{�{���u��u�$_c��n�g6��q��=>#��S��ɭՃ·��tPO X���g��u���b+;�wd{g_ڗ��Osz��f	�̆zo�G����ɳS��w���û�#�uߋ�"˼*p���/;;[����<���f~������8h�v������W�cS6eS6寨l�MٔMٔM���v�&�ق��6��P_iGȾ���W�^���5��a���X�ЅƁ��fK��H�F������'<�FD$H��N�"
�3  h (��h?Fu��|d���u#�Tk��@�M��������R��[H`@o�&��Z ��_��AX(??=�ϯ>��A� k��Lc��8lB�!o�)?�{D�)�{�{���c9:�+o�����O~,���g��/������ YJG�$ԯ4�h2#�p}kgO����� ��p2]v� 	`�9�[G��4B/	����z�3�06�8c?�8|"J|�mPa,Ea`��I� �o��4�p?`FeQJ�grDiRX �yb�XQ�G���x�1� �O9� �D9�l�����9bT3"ƙ�	������I�j�7�k��)��Tnn@�}K	���=a4e��n���$� �Ȇ7H�����i�oˇ�����|��WrzvJ�QˑMY�x���<3���l���1Z�T	,0��AdYD&�;]�W1Rd�&���Ch}�:����+�����Y}���=�z�@(_Gj�q��4�A�!���C �L�,"P��@ۉ��7 	���(�j�����K��w�Á8z�c ���s/�t�`�K�C�k�A�Sh潐<bW��d�j5��q�!����+�*R]����>D��e՘�A��ݚ\��ru>�f�_h��e�B'$r�X�2ѿ���h,O!ϯ3�ޗ
a��j�K����ѹh�F�b[�:�J�g�/|r�� ��ea�J��¶��7�fҐ�4�&�Y���������������Ů/KGF`<FuI��p]K�˲8oz B��}Q��z�)$��ƽf������+�a���$��>�2|Ν|\�k;I�̩#�.���(�֢�m�\@��*i	�yӯ�=E��W������D�]��E!�m�[�<���&C>�e��w�M"�ȱV̄A�>�J\'�I�!kHW7�6}#y����'��d�
ΫV? !�ۂ����we��0��$kB��d� ��4Q����kU��\3&$$�C�����&;�s2ư������sLVݽ�܏k3��6&9��'�4�5Uכ��Kk�)g�"�)�l�@�W�l(H]\����dg�'��G\�p���Vl��
R�5���踴� d)D�ļ�} g�1�£#$�%Ȧ��%��n�׵K� ��{֘9fRiS��&��Y	�����;�kbJ�էO�GH@x��@�1ÄȈ�K���j �z��@
oCdfޝ#�B��v��N�t�j��@�1�NM��;�|�c��lw[f�A�;3�;��?��� �x.��/�,7�wJ�Ӈ�Hns+9#��+c�2|2��$���@�I��a�r�������'����ơmO^����/�v:��S��	��9R��-�y�Z�����F�X/1�1�d�N0HC��728 ���o�kw��c}0
B�Y��R<�z��4�g��(�҂\����\D-��E�1�\+�"Mm'�;���"��)n@k�d<�F���U�d���6�A����u�r�=12J@����<���2O�WBP�8�0Z�m�W�W���u�~����ݻr�����~�l��5d� 3��۝=�������+�}��AHh���$^|�k"f���q�G!��9q_�6�9������vC#����MٔMٔM��)dS6eS6eS�,
�T������%�*;��� ;�(z"��`@И�u���̺��������!೽ӣT������  
`���`t�3X ��}�֌�A#h��kIz' #�F�ؒKOf�Ϻw�P�������0:� =#I������ȗ_~)�/Ox&>�C�m��!���ٺ�E�w���=y��C��!��?����W��<��2,����X�2��ǽ{w	N��R�Z�3 t����D'2*�X`Ƴ�}���P&����A�� Bd�^��t� w��6t�����RK��@M T�v��9:Mi��v(,Rr��<L@{�aJ��3�ƗÃC��}H�Ue8�33#��1+���[�,D�R��#X���K#&c#ض�wٟzz����յ�E��GO(	q��Y,͠��w���� 䃬��ے��+�i,{��g��wdo�X�灼������˷O�f�es(�U�"*A�n�`f<9G�̙��� c�,����dOd �ƣ�T�����v(L��wRX��A�-�o'+S��#�|�ݛ䕷��Z�<�� ��
��X�TM`���:�$Y��,e[���)',��_E�S"(33xꙻ��ٙ� +_K�{M.�w�sC�(�1��We^���bF"Z��j�{��|nr- |W���!Ȇ ���2���.���Ր��ґN��V꒒�3u�뵗������NHn2�ra�-�ec0j���g)�A�E g R!���%��<h8�,"��RA�#T"���'\���tҹ.���̝L��.��66QG���@F�R	���M���У]�3;	@ch`+p���vH4i�u�@�h�U_��B�=`��EZ�0w�������ħ���e@L2	�뛌ߠ7���{��2C�r2? <�ȜA��RS-Oطб��к	������0j?Li�������E��K���Jյ>��<�������}^Ws��g$���A
� {"_+�y�3(��+�zK��B�L�#1��\�Y�m�� G6]`�X���zi���Hh�gx�x�o��<�%�k��܍�#s�4ݰ�ď��\[	I�b�b�/h4b�2�c�x�IM��Ky�j*��P_{W�����Y��CK&�� Y@4fw�%��d��NfE[�Z���3�cJ/���g� ���OP9����X;�k������[M�ip-HFz�"��X�Z�����k%�K<�7�u��oh�}a�cY���:?9�'
�3˖dF2����;�x2��8��ӏ
�^�@3��ab��9�����u���^��ϐr��l��`��AI9��i��u� �ْ�Gw���rH��e�
�$�������9CFR���ܾ�
�yN��7�YEuiظ��O�f>�O`���xGz���;Z$W�i� r�}���*)�7���l}̙�׸?.�����,#�{�W���g����jȄXZ�
dY���$�H��/�G���V������$��S���8��/��-9�8�WF�������~�|�l��g���=��������ٖ�рO� &��p8��*I�9�^��ɋg�w�/ݭm��5��{Df�/���m�5�l�I���h#�`��t�t��^�R�i�)��)��)eC�lʦlʦlʟE���H��H�v�A�����#�U�n��jt���L�'�_�R=|L�� ��;��J�ݐ�l,�n� & D���R�ݢי= #�:��Zr��y��.:� !���u 6�O������ѝ���X�3��-*!��:��kz�M$��eog�v��Q� �!����&��<Ye8�J5 ������*�{�����L��!`��>5��	�gT9�sW���d8�w5D�!j�?���Y_�����ՈQ���(J�������N��M�0�O���"(�t��<d	�u���C�/c�����#�qvuM�.�W#2�+���LX}����)�� ��u_>���:;���s�"Y缯�tDid�l��2y�� WT)�B��$����O_=�v�+������w2���0�Ϊ�CMmn�v�e�D�Ti��r'<��Y2 ��*Q�*~ܓO?������O~�����Q��,���#0�S}�6��Xp���@�%+��r-Yf�� �K�<�g+��ef����e5d�j [bw��Hl ���AA�@�$�H����	�i�Q��2uKA& ���{��K�~��IǗ���J�"��-'k9-^�}�1jܴ��7~��|��!��Ѐw�S����W���G���_=Ai��*	�8�$X�s,P��K�Jw>ݩK1p��lI|��검2�T�VBf��k��y����}��!˅E##H��vn��0<��4���b�}w���2$�X�
@�E�u �njϻ�.f�4����$sF�6�VJ�9;�xK��OٚX������D(���VkK?���H � �D �YZx�gAj�D�����+,K(�b*MY&˅�����DC
���� ����:1㐂 ���Ώ���9 ��DF�˨�u��p�5Hg�`�Hp�,1]('�@��b�ݘ0�\k�Y�0��8wQ��z2��DfVM�� ;��R��%���`��y'$�l��̞���/���ÜͱJ.a�KfgX��ڂ����g���������[d?2,�Z'���[�� rzu)�o���#@B�lq8�<�� �J��Tn�Id���)�w2�e��y����$�r��pu-��	\:�๶C荶��]���5CbT�M�{D����O��=�8? x��<�+K�sic�1c���M�}���Y�;���1Iت���]�'����4�˳�6jz�m
���y�*��$�4���� ����,N�#�}}�P�?��m]��?�����szr��<V�!3]���>��!m��!#�ӗK]_������F�yw�G� �"�N��H3cu��ü��'7Fm~��)�4�U�\��UtN	A]�9g�Y!� f)_q�S(\73�}��x��H��ͧ/��i�|a8����<�(��� �y�޶���X8)7#뒹yGe.X�ȸ­�N�XI(�R͘a[p�όX�7�q�1}�ciI���1�}k���9��dL��{����,���>��LJx��:Ɛ���E��'�|&��O�^?~L�8���xL���i�^�ͽ<V���},�7al"cv���5��L�D�Xg"���ܑ�:=yA�,��އ{�꾽Ӫi�O���R_�\:��uwpt�~5�f����$v�^���5d:�^]_Rz��h1�x�c!�
yS�sS6eS6eS�:ʆ ٔMٔMٔ?�R�ʖD��h������9;ܗ���e>��6�&�-S=�=�������Z�!~�F$ �q���`��@j6���_�W �AT��V��i5�2����bm"m> �Fq���i�������/f2�x(K�'^��G��/�."�����������h,S��6"q ������x�6��Á���#�����O�����������i��
`b�P�}�}f��d������~�Z�~��Z@t3�r}g���DU��Yj[��\.[ @��n�ږ)�3P�J�2$h[D��� _��C����|O@x�C;�p��R�{�6��%��zQ�j!�M#��u ����F��e���/�ۉĐ'��:��anZ�e�5���`�IP��M
�#�L�R������͖d�3<\��dw������W���0�P�k���E���E�m�����z��d`�R����dJ�Nu��C��ht��<�������}`�6��s}/��gi*N$<0�kSp+�U%I�6�����kt�g�.d�s�lv�j����Y���Y�A��4ms�F�Q� @QIs�O��`���(��(��x�y㵫D�w�� ��A٩� 7F�C�*�1C)\����<C~(�L�/�Q�PS~�<e �����eB������w���,���m�����31���ˠ�k�`���@2$ �fN�?�0 ���{�5��w,K�~�I
�ކz%�l�B�Qֈ��d�W�P�j 94��VH2��3�G
M�$btw���^q@/�����G:�8aF��@��3�4���!�Zg�E6�  ��IDAT�ԫM�P y��w�|�=��NaT�uL����1
 �YS��|-'r���'��=z@-@� K�"<&B˞�l\T���(�l8�hx�B�|l<��̗ zA0��!���O�GV�$���gc�`�y�)�����L�`���M���2�x?+�r���(�x$� I�z> �)(�,Mi�d�k��@�g����˘ui�%�оȎ!���j��]��MnG�	++	�ދ1�Z��!��x��푹A�Ė���Ϯ���E��X�?�^<B�C��IB�>R�\Ihq*-r���J��	����csc�^��B�@�|n��������F��A*�ޞ|��#��x������s����r����E����� �؎�`i�$rf22�'��~���>�t<�����fm���^�w�Oe4�XF A�{��9f�T׼)		�wZ�����L�u����g�b]b B� ���׺:99����J�ϯ8&���1q\5,-�Au�0E�'"���}��k�ۡ`!����9;9����䪾��[k'���-��jʽ�/�Șu��;��sA�[�@��N�k2��H���ʙbA�'���%I���������2�\:B�t��Zy��ٸ�X_K6��eX� ��l���_F��l���C� o%dd$��@Ҳa���O@�@�����駟�g���}{<1���QC �ںW�~{\����.��7���
"Z���LY�ӹ����[�wpH�8�:�5,0R����f����~���D溯	u���{~$����2�����C= [
�1��yujc[2x�aUƺ/cf���z��)��)��)�eC�lʦlʦlʟM��'Rݫ�l:�ɨ/�nC��zH�ݖݝm��A-If2��0c�Fz���@����@��������T�)�B���A�D�L�aF�mwx i�Z2�c%����A-���.��ؒ�V�Ǉ����Ⱥ��Vn�C�0eV�P��L=�%K��<�F�)��D�/�(I���� �MN#sQ��ĳD����@l \��r��`��p�Q���{["�	�c=������ɇ}_<|@�\�kkOG� �7���uUkY0�/mŨ�i%3B�ObB��_&K��ptF ?�,�,��5$���BEDA������+sY��B��s �e<�%�	B�Z�$��.c�}���!�+Jϲz葍�g���rzm�I'-(m��@�S�6�H|�Su�孇{�_\\��ѡ�g(�H�iYAY �F�b2�I����8M(U�w�+?��H�y�]�k�O�c�m�:X�2�����_p�?;;�z��ς��"��!Æ,�-�`L��	��1(�L��D�єIX(Q�"�����w@�_p��֊�0�tM�h��3�`
�Q5[d[i�C��^������s�j8/��fve��DOf��@쇲~
R����4��h��ILp��,������f����g�N�)W_ ��u�F{�L�_ ���}��^eO�z!��_L�)�5!g��g���0��b�|2'a����h�G���U p�qZ �+a�s��cu��I��929���e�fׁ��ER2�/0~AWl�`�/!��`D7y�U���Q��B���@#�Y@�Cf,�<݄˜B��	(���� #�c�+�+��t�t:�l�b�֥f��J���#)%A[�3 S#\�Љ��T�n�W��3���sy&�����l'Y�o#p�ݱ�3�o��$������O�Ii��h3�1H��K#� xj.]�c���*i��������.�հj"@+�;�|>JW_��9菔LҒ���j0`/k���(F���(��N�-�d4�a�X��[['I�R�_M q`��|C�Ǧ)���(}��3�u��Ҙ��^$���K �-��7�L�t�=.����Hʖ��h���@�� �x�l1�7Ch � �J/����?�������|��od�?���v]g �+���%��?q�d�+1	6�s\�^&�����|����k�f�W���wvz�(����3�%�3�Hp^�K���� %W$���"xXM���2E~����?���ꂁo�$��L^�	������@��`F^�p�0	���  �y-_��72�dkg����������KA)51�'��L�4�2wcE�3/�<p���Ը��������֛j�z��\�)���yC��I�9��՘���?��A��nNA_IB_�̑x �����wػ�ώ�c�.\R��G���\�_c�dFT��v�5:�.�?�ar����k����	�lUC���}`I������'��,�K�=?t�W����6�/���V'3��'b���Ɲ���t;z�ʵ�Ļ��{k��h,M�o�9d�`�1��1*mۮ�@^r^���7�^wz=བ��P|��*����MٔMٔM��(dS6eS6eS�,J���ã���ř|)B��$��`�x��/7�$��ۖ��\�Ő�/�=���aF���Z�0�h��ه2��};t�f`���7��h��o�xN+�tf���~?��z� ���E)dA� �@��Q� M�c�� ʷ��:���Dijʛ,�"]����н��J��RF�1��N��L�[Ͷ��z��!�xH_�����׋�^ϧ�H�(Vu=06�&���Nj�2@V����Dfn+�l5��¯�h}���$K>s��6�{�=$6�ˊ�g���(�* �e�т,�ި�d!��B���	�ֿ��o�Y�#��t�^��A�� �Ф�׾|~�y\��q�Q�?Ud-��o�:ǟ JDN�"q������D	�+C�m�0�,d�ia��v��Cz�i���ɉ�dV� 6�������?�������W����������T_��_c߂n8Mz���>B&F�"��y Z������D�,�Az��W� �?H�8���$�C�`;��_�C�v��y!|.��r 2�� 0���
AG�[��*�����������WA����4QP�̴�^���zʇ��)H��,�J��2W���t��ڮ�y�RF
Ø�� D_�������:�#�B�y��H���:^�"�xA$/��b�p� A�| �J�F0���HA�#?���6KL���}Fr��K�.�F�}�E�V�:o d�f ��>�g�#�ޜ}��q��h��x��P�"�K�򢝉g�rN��"K�@RּcHRČ8�`�@�m��u��@.��<��T��dJz�~NI=�t̨(+�:������  J�1�I��L�u�2,���e+/ܫO�8#	sF�甗��6����	8�+�~��Ј`�+�d�3!�C�6��h����MJ�<�{8b3��|��!R�ְ:��p>:+C�&���s�x;�h���^�C�7k~����UvI�4q�eY_ko��kq�#1��W�:�__)��A�Է@z+��������2!���F�8����<8)�z'��2@�_���k�6q�{%\�о u�"z��q�d2�˞<|�X~�������ŋ���ŉ^'v`�=/�V(�Tq��k`~V%IF�C#�Mc��3��8_X�H����0N�R���;���O�W[���2��đ']�ݓb�G�Kn~3�[ �#��t��![���\��-��kx�/�������:y-(�!��ٵ�5u�c6��E�'H����i@�ܳ5hI���N&�/����ϥ�l��ѱ<v"]�jՊ�.��Q[��g�k7�@(��2���/%ܟ!K^<$�Şq���2��ӧrzz*�z����� ɘ9���;��	�<���<+�j����FF���`�B���!Q �7�E��+ք=��<�����ea�2w���w��>�H��-��!	�t�:N�%I{%�?=[_��j��U��5�	4m#�'��֯@����ڷ�6X�YG���t���A��\�Mm��qsp�������޽{�ju,�Fk׃.����!�ewk[v�vH���䧿���2Z&�G���_8�lʦlʦl�_\� ��)��)��'/y21�hϲ@f�1ʈ��9�Rd$4�`Qo8D4u$�1�=	ψ_~��j|���i��f� N��.�*��n%-EOD�;�cm:���Y�o02bɃ=��E�hr��SD�X�[i�ql��摬��>3��)���&SzZ�������H~q�^ɂ��p ���#�_xT��v��h�-]�\��}ppH��k�l�4B�^?�̤?��م$�m���ۃ�g�����5�Zd��I�N ���gp8_E���zF��Łm�ί�|�.r�u�)k7*��/ ��H�|�x6�
��B��B�d�ԣnIE�	�iݴ��3�o��F��/�U�����-A���>a�1r����fT�(v�������&8T�yB��Z=��M���m兒 ����HRe�cz�D�'�6����=�b����޾�>`�ȴn���)I+�� �D�F"=�� qÜQ��E'H��K%���C��xZ�ϭK����о��Xd;A�f���n��q�ݓ'����: �h~
 f�Hߤa06��(��|E.`[:c����B���<j�S�?0�&�yDi��Q�!�%N�(CD8���N ��r��9��}fڠ,�ב̨D�a�8F�=��y�$�}�2�Yr�Ձl�Li������ѪT	��*��Y v�����>%BP-=��2����y.��ܓ��I � ��[-z��\P��A���dN٣Qlq�4��C�b�3�y�`d3"lA��a��n�xM��S�p@C=��ӹ�y�`ޡ�e�Z�D�Ih�jX�Rr�\F��23����^Ч���e����J�Y���{�D�9�;r^ �v�=-)��~�KiQ9lc�T�o$�^A���s�+}Fw@.A�
e��}rd����/��%�@,��G̐o���[ ��`_�q��l	 p���|�+RMN)u"θk���|?@D��RX5��)��9�8Gl�4�5���u
��'��"(8�G����jU8��ݔ��I<לLbfd2�:[�5���[���o?����ind%s����=~x֠�9,NR�wa�U��b�/�|���Q@��.��͍:�!��y>���f��KΏ�&��|�0Շf�����t�C+p�,]&e�k�|��SF����\��ć'�tZm��a�D�����\��Z������ �B�[p:�X���"ˤ�m
@�I &����'�|́�h[��Mt��@E�~��=:�}I]׍{�ẗ{d�â����{�)��p��/pV�S�WM�}ي�]_���|��/u]�Z�c]ׇR�{��Nr�3�4L)ۈ��Y�FS��z�/���ļ�LI|����Çoq�}��W���2ӛ�M�����
�
��|m�*dP�y<L����0G�0o t�	3(�s�s]��}¹]�6�e�!�� ?�;}�J����螧ʌ��_$@�q��D&Y�ݹ^ KA�ʶ�]`FƾY8�Fd�����r||�d�����,��8X,��*��Y�>��>�����;:8��"�w��w�T�X��^6���^�/����Y�(�/����E��Q,x^��*^��/0� ��kz�����٫��$��ޖ|�O��w����to]�D�YGm�kv��y_Xי٨uYH�sz��a6[0A刺�y��^E�êW�B6eS6eS6�/�l�MٔMٔM����l��4���"�v+��.d��}���U=��bn�����<�y6d{y���!۽�~��`o�iĐu�2���~�A����Џ�f�1N�� +S�XVs=$'I`�ِ�
-j8
�<<� �����$�)kS��	hƳ9��x0\�Z��f����� m�0������ۡҢ��7 �!�f*=�����$?�����������*��}�D��8 5 n � �{KO_�$8�����X$"�3�j�(p�hI>�Ygh1�,�y�$�T�/)��ͦWz��$�p�e}ü��)��Lf��eD=�r$x%AP����E�Ҍ��M����`�,�T�/ } ��®IPـ��x*v
���������}~�4�M'��)����H�w&̙�#`�v�
Cfs>O��J����-�|�����^�������C?��եd�ݻw)}quuE"�;"����EZ�
t�������@>���7��w�F��8��Ғ-�M��3��� Xw&ˡk��A;����`�E����>�_k�0�Yg��ה.*�7~�ٚ������l�6�T�{�P+��̙��Fl��4��gx��	���&�*�ί�Hпf�6��t8��>S�3ZwI�J��#�?$�	t�S�����#e)�Y<2�z>��)/�zf�F}f\�<	�[f	�]!ɔ��18�0��1�#�}���d��d�YF����z��e^0�>4oz��4�-����mN�@,� �2]���0��ʢ�c8#�K�'YT%؍���l �*Z�5"�&+囜S����e��`�j��"k�XI�1�(�k� 2y��Ef� �K�WEf��jS���/�o^�d�,�/+l}��a&�̰)��~(4wv.�V:�#dw�z�;/�{ �����U��#� �|��Niv�GJ��U���*�������9;��9x�U!a_�?���������Ae)C�oYW��<|�e��e����\��K�оd����ЃY��v��إ�B�a�d�=���`�~�y?��3�I����^K�dٕ�vu���*K4z r������B3�����@ñ�0��꒩*Ed����^k���{������W�?~����Z��?q�Ɔ�A�K}ٽ�s;����r�s�W_}�*�o��F�Oϩ��u��s~�.���!����܁��&!�b�����:�U�*'#?.f�F��O2 s��T�:�޽/[����h,4��Gfk v}�! _����u��)�9�'��Q�6N5�L�E��;��i%�N��P!Tz<��6��������م|(�8FJ{f����G��G�(�������}ν_~�{�!a_�쐤���\�W�F���{Ť$#�3���W�\�H��0aaK�������oF��漌9a���g��[]�����\�}�롰1uP�[��	T������#|�����ުs��X_�B�N��=0�Q$�'�{��.�ne�Ԯ�2%}eyU�ؿ�^�{a�
� ���3�Ncy�L�6V��[�Iv�X�������Z�bFLLE�D�,��$D� Hd��������}�9���)�3w��G�����ɧ?���{�H��u[Ԏ���k�(22��!�p�L����>ԎX�a��;��h����������_ɦmڦmڦ� ۆ ٴM۴M۴?l���N��Z7y�n�M�W=\Ƚ{��
��ƫV� ���������P���o����t�6�w�%[[;�������J�_�r���P��hq@��C�܈Ji�����5T�5�� Fhm�=ʮ���fn��Sn�:��[��>ϩ*��ylVFP}�3��ӀQ���;���W���V� #B��� С,���`�ߘ~�n� j�rrE�,T����U۰:�G��b��j{�ᤴ�x=XX��s�}����<�!c�EӘ}�� ЅjJ�=��Y�%!����;��㇙i�z�ӟ��i+*_.����mV�n��2���b���<�5j|g�O��h���vovn���F�5,B"�|1̢v2���B����N�
���D���� J樴-rV�bN2Bn*3�D=���l��cFYs�nF�5������fc�� o 2�3�nBIq^��!���"��7 >���;88�XĵO�أ�,,���-��3���}l��+�0F#�q�
!o��tT���0Xhr�}��o�E�#�� ̄�o�pH�y�:�9 aPu�`.�[�GX��ߥ��X�����J�
�>3.���$�����a���jr(M��zP'DE�Ғ��P���z���SU���r^[�De Z3�s�r�����DX׬d7`?���M;$�� 7�w@E�։e"�wE�� `����_�i:2�T$KAi�~�7 f��W�x��X�y�O������O�$����r�冒��vb�"P��vU��J���Tڋ��:�<�����07�h�"����Z���A�{�.��0r�&,h��8���9�W�DV���	8�A��T��|q���wF�% N
��
�ͺ�V��=k,�Fh;����k5#F<�\	rLD6p�`]��v����u�gE`���$$��v%��y�p��0J�
�p��l�2�:��2|0FJ�
�zL��ӏ>䘟����N�G>T�@o��#}?��}׋Qwۑ���$�57��2�mSP�w�źr�܈I1B����B��gsQ�nWH7���+�;��(�v��c���<dfpM:������p�%�E���_~AU�!�^>��Ͽ�J����>�J}n3�k�`��~�����5N�����3R��
BSL���~B� H�No����� �A�EF��֬i��PŃ��s�	B�F�gɉ12��t�+�-ǅ�wwoG�I0XP|F�<K�;#��5ֵ��Ύ|��O��>�Go=��`�c9�����O����r��<�c6�B]��5�ss�*潹���l����1���۩A�6��Y��5u����Ȋa���R>�я��>���.�_�x���L�uk�S���[V��0�
?��^Zq�#���9��?|f����4m	�v���I��L��(,W$�^؇�x���.��5]�XK`�jj����h�#�|ߘ:�1�8>3�H`���6W��2[�gg�씵��Fۻ��+�˿�����\����̫5���-���J�T�8.f<���^��R�{�>W���y������k�������k�6m�6m�~pmC�lڦmڦm�U� k(?fy��5U g��Sۄ���ɔ #6>s}�t:��=����B��R��B�N�u�<����?���l�ʬ �PE��� �Q�ǪI�0��ӖJ<�4)��R�V9�y���Ga���Ym��dX<��1�Ya#9��e���,�y��Z l�C����U��,H��syy%o��9o�e:���z��H�{��Dup�&ȕ��R��������+V��*||�	�ڻi×+30�����M
�����+�6�$y��D�v��A�a�`0+H���O�sS���_�v�^��k/�?W:6�Ja�k^�  ��ˬ���\ �:�/}��?͊�G%m����  $r�����YI��"WY�e���|�}��;wLH�@
��j��hv eC�W���܆��'������>�5��,�潍�������+S�����Ju���xsb���P�oXxDPX���3|PLMn�� ����U8��X[}���fEg��zY܄�`�(�Ñ�%�,�%��z�u���b�kj����V�B�(4�[u �ne���vc�����#2<:V	�A�h8Tl�K�j�v P��^�nI����{��$��V%���$àl"^�eW���3?��Vtn���푓��đ�6��_��� �h���hG"
 ���^�W%�V��<kɈ�mQp�0�L����=Z@�9����E!0�� �˼��0\�����f Yǂ�E�y��xϱ�%�x�JC��̥��+-�!�<��hy!�cSX�mWa�� Ȼ�g:��uN�$����T���*2AH�#v�ǖ�'��"��A;��iD��� n��b 2ȕڈR|�q�a'���D�	Մ$$�w�G#f�Ք�J%���8�����h�ƈ!�g"��	�3����y���R�������ޗ�����s���V007����)�}���W�}��;��A�C-���N�w+D�r����Z �>�l���8��6oVAj�����a^VP���9��>͞e���r3fW��ȫ���x�`�:a�X���7����Tz��\����A��uC����ڝ/��1H8��\ ���r�%���9���`M#5�3*6���\z�����(]seK�s���;�@QO�a��7` �.l��,d@aH(Ȁ��a���\D�����ɇ~$w����p��庵%�<�����wtG>z[���c��8ձ���)����[|N�^�R`����U��pв��6�7|.D�w�Y)�s5��N ٚ�)S��Lf���nr}u�HD>��e�qP��]���c����fF�?�M��s�Z�%",�p�@}z� ��c+\q�,
w���i�'S�8�Լ惾)�@�����s�,�pC�9G{U����l#i#����HR��KZ��f�5 �?'�R���w=O(�#�s� '���9z�;�T;�����?�W���������72WL��c{������j���5�,([��0嚎��x���'�3������������������i��i��i?ض!@6m�6m�6��X�&��/c�הܸV��$�3�#���x͍N�a��lmo�Z�f�zr%'��d�"� ���nH����ryy-�ߜp��,t�|4�E#��i���
�	~� �Q�%�]�m��2_�{��UR&��<����t���i�z8O�᜶<�7�#���~�	6��$��v�����t��Uw�ø��Y�MQ@0����U���S=@&s� �aO�t�ղ�XA��I��,=&PYF%+�)�^��jxe彌�Kݮ}?� �Њ�l<`q���� ���n��!�s����S�Nk�%m%4+&K�2��4D�\��+o�+���:þ�\zқ�T�&�I�B"E��ǶX�1��.�>�CA��}yu�����=<::���H��$+�q	Ƨm�d�@\��?�I�3������� X��d���!ؽX�d5_�X\Ӛb���q ��%�w'��$\P�X��f��L�aʴj��1��|��q�� �#_����GdC��F\$����\$w<Ûقp%S[9�!<>���3!�FK*�|�S���&(G<D���σCR��-�A:��$2�l�b�O�5���,y0�Y�}y}�<��`(*�a�iZ%��ۘs0��]c����� 'z�u����g5����2z؟��X��t�yХu���bP��pցvdk�.�
�j&Z2��l˷@�5Em�k�!�!�6t*�`!0X�2�rK<�͓���@�08\��&�]^�%�F�TV���+6("Q vp� ?���ewf*/nL]��� �욹ś��Fx51�œ�ò�p`/��c�V��bD�'-#%\�H��(n#H5I �E��z/iǫ�=#�����,�`��ر��`�s��H��+�b�i;��II"�L`^�=�D!p�,�сg&�H��*���T�d�`W�=�N�z�L&W7a� 2�ܲ�J��+��"��.%�0N �U�'��-�!m���l���m�==/�����9P,��k��3.̅$@�>��tl^���=��ڄ;:�'��ȋr�)�|��<~L��e%y}�c x�l�CD�'!	4�?Ca�W�sD��p�,񬞔㙶n$#��b�F��c��5u�,�!�=��w�ۏ��1c
 �/��9՞[�����1���A������9XeIDJ��9�,drx�/�#��5�0������\���{P���;������~V�s'��K���*/x=�$��U�ǌ9j���1*#O�,�uZYz�Յ:n�:'3�n,;;ۜ�@V�y�*�B������z����ˠ�y2 #�����+wSf��[C�Y�X_-��,�v�Ṽѵ�gל_]���O�n�#���R�=qc݊���@1�)��t=����|�507j݄�����x6�J�E�]��XK��(u��(�Mmcꑆ���	T S�1�;�|^R��� Kak;�o?�:&wu>�t��k��Z�˱^��9=9���r�<�ãCf���@� S��O�D>��]�nӚR�G���^R5��_���������ڴM۴M۴j�L�i��i��G�j�PZ�V�/s�Hh�n}���M4�:�$aؑ��k�H��L7�H�������E��+�, ཮VT'ؿ/e\��
��m�\b��U�aUe�j��.�.���g���`��M,��4��R�	��mF qkQ � Y/,ˣ�£�z yق�Tt3*bXS��7��TD�-������9��H7�V�wΐ��A�@�i�1^��5�k�.A:ZUTrcѕu�F$��M �B����7@Z��u�F� �"S[�+��ϰf�F��*ǁ�Խ������5��B�8��4<F�eܞս����X�j�8>��ȫ�������S0PT(���ˣr�s�G娾�ի����KG��}�̃ȃ�,�����[��?�e��ǎ
#��F��Z��y$P�d�C}=�q�<�e&�N����Ņ��"��	l�z=�\�ng�0�iC����W����U���G~��x�����r����Pl �I�<���G�q5ù�l�Rq1R&n3��яMtsQ*�tI��=����fY4��;XŚ��N��b�C�Ԋ���>����^�  ��+��k�7��	����Ύ�z����_~)iw�߱�`eT�k�C=��F�B�1ޛ��0vKU"�W!�jlڐ`�0�U�@�Y�l���/�5q��zR\c� �lطU��B`6JKڅ�?��r��AFX_TNRk,���ߡ$�C�MҪ
Ti����,�b�:4FT:�ޡeVB"��+<���ġJ�J�832�0c��(�jy($%�\��������>�M��E�e�ķ,����X!Q�v"������4u��9J ��w�i	R�9����R,]E^�-��AA+�T�j��9U@���ͫd A�EIK��@��2���o��Ю�*�t�ߙN�8B�x���mǯ��Y;ѹ�ڀ��6q�"���Zn�A���L*S���Ę/Aj�+=&�x&"dDW�d>����6A:���������]�IV������s�����j�sm: �g�p��f1Ψ��5�1t-K%�P� ��#�vԳ�8n���p�k_By�ͅ� �x�?�q5Pv���4%9�5�|t���ޞHo$S}.Ⱥ�}��q�,ب�`���]�I�>HNZ1�Uk�ҫ	vn��U%�/)�<�� �$E��5��ω́ ˗�+*&1�������#��ڥJk�1�߹+G��$�LB):��z���yb�QX�1���eϔe��V#��H`��P�t2��@~ܿ�@>��y��w�Y���o~.Ϟ|+��+��k�.l�Rα(h1ugb�.,�������I�*J�$N'A��MyW�?�L=%�5Jx�A��_\��@H`�م�"�r�\bs�g��B�*��Fb>����yd���x(&��Z�u%���u<�@Hz�:�-�n��+�[��	A�x�&�kyfJ�k�Z���gc,!�c[�KG����}%�*~����|����O"�=�Vө,�3�k+�PRnm�9oB)>�ޑ�d��5��F��1��J�=�i+N����k��i��i���md�6m�6m��(}�K��v�VyA0I�# v�v��g��*����ä��{�t��^7q������a#���d�$+7���_b�M��t"]�T�I��Z�@T�e��ԦBh%���z����h�rzz*�і�t�	>B<�1E�"*��@<H��^O�C��DH^F;�P���d�j�I���.�H��_��'O���@��@��~#�w<�湡
r0��l:c@z�߿\���� �~�@7����Y hq\YlcU�d��U��F�_(�N��}P����yc���_k���h��;�E	7Ӎ�� `���|������[�5�7�^�Cdn��r��A�j/[�՘�ô�?>2r�R�<�@a��{���ɂ}:#k�C�iw�H��{@�Ή^�'Ͼ����!��zy1!���"�-�@�4Y�68P�@	� �+VR�=����|�����%�@
Q-����l֨ڈx� X�Z#�"D��7��̭?�1+�k�`(;�nNT���������2�*ب��TI�*�۷���w�����K/rY�K�Ab|�ĭ-A��3<X��� �Q�����v`�ͦ	�J���7��8�� c6I�@G�xM�����c�tEev �`����\N�/tnۖc+[����J
}��=�6�*��.	���ob��g:�x@���R��9�J��-�ȥ إ�]#�zm�YN��A��LCk�ggTo��� ��x���v��;F@`7��q]D�V0 �#���qo��J�#������ ��Fv
I3��U�G�V�6�yc#�X�,�*� ;��J����k�[a�U\��2��N���c�nqm��"[X��,�nWf��&V��R�;PFU1<�ٌ�< �u�KW�@<r˶ď���P��VaTa�T��/���w��q�L�aPb����!����ܜ�s������%��:!H6�����brǪΓ�0 �R�P��{+}�b4�`kD�H$h�:@}	[�����y����;o=�:�(Td��t��`�&�! @��7Ȣq[!�OU��s��]�1�ôa�Foz��D&Hi}^���5�K�5UuW紒�p�ϔ���J\�RU?z���ވ�E�ٹ�I:bPB�E��a޸�3sY��ȝ��J�k���<���~���:ewG�M�,0`�LY>3J��f�,+WP{�X8���l�ҘD�40g�����[� ���؀��S�&�OX�@U�����!�V�w�b����cI{����Y��z}~.������뺧���������'�nX�i���;]~-�tL��D%�0`����o��Ls�ዧ���;9��V�u�)y+�&�V���5-��k��95)��ٜ[�����M�wL:�F��<.I .�LS.���Qٽ��*��{P�&�؛af
<�`%u=�6B��՚v_f���>�:R/i��n�� 2��Qa�O(� юgG�>�e����+��j#r�*��R*둈ǵ��ҹ�js�W����7��_�R޼z��ejZLF B���Ws�O(�@�ɋgO���L�?��N�k�O>��}�=nڦmڦm��m�M۴M۴M��6T���=d��<З :t������]y��t3|O����7''iܻ/����������L��Wr����B0�����z�ZV�������&����]�u����m�������*��r��~^�� ��G�,�^cS���$l����n�ʿn"�w�>|s<�L���K9��H�̬�������T�j����Cd4�k D��7ή/��?��������7�2��X`���_�(�V
��H ��8(�$^�l�Wdj��)K�j��C{���r/x<	�M;�6�+S��qo
[��I���U�BͰf�g���2�U�PYXqY��DT�PY�K@�c�\,	"@x*�l�d1x�|N\�����1�Hx൨$F�3� �N%�����t���Urp���O�T��}`��5���\��mP�uM� � ��z ��v;$/�b���5 G��L�-�\�;�9����0�r�W�L�g��쌷���\���&3�Ƈ]EGǔ�h�w|�ʰk���Ca��`��ZUF*�g��f�ׇ�S����/6e��Nog{����q��WC�6�Q��;/bul�> ��1��ʂ�9���&���q
p�� 趸��A7���m�(��#!P�܋��▅�6��M�D^�Ғk���~���ܵ֯AX�_�^��9���h�:P!o�{��M��:m�L5c�7�	��,h�o�2�@1�Oa��뜑+���o�l��<�;�fT�S,Y�EMuL#�B��AEs%F� �G�/sIj�ω[����e�fN�����̪�礦��{i㠜���=�ƭ�@���U	�7e87*��K��'�7�7#rxx�_ق9�r;7&}��(�$5����
ų4�)����t�Y� ��T�.q�Rd�⴪��f����@��V|P5D��y��8o��d�wtC�z�*vB���Nr+�F�Y�Z�Z�`�g��x��}ȹ<���Ub0$U�s��^ X1b���5$s��s�O���{�w�c��Ot.�3����j3���>�0?E�d�P��*��֘�J��ȍ� H���z���=�
d5����P>z�]���G�2_LIҔ�B���~�����$+�uĬ�eR0��*��$���$p2�z�]]S�eJ$S�9f�5�)L���?�ɥ�
���zA��U˜���E4�uek��}9tD���ՙ̗>�@�����~�������9�k��Zxf�{x$��y_��t*��~'��J�%��-yc�im��[����b%�ze����6H ������
�2xN��eF�V��y�\�t�s̵r��'<�{݁>G�����~f�P�х>�^����y�k0��cV2�Hl��L�u �5e�0�d����������ޡɽ�o����Ҋd��',�,�
����%ׂqg�Yb9	Ţ\�[$�@�B�uU���y���1�L�ӕ+���*�v^�B&�B�s(��C�db�����`^��KZƢ_@��s�dr���%�����!(	�f����G�8c2���8��MHR�p��}ό���	�:˖�x�X_�:�)2W�9�u+87��X��ʓE��P�B	뜢X��/��0,�f\��<��8��F?�8��P��֧	-̊���C��i��i���jd�6m�6m���͋�,@\7��ܬF`3���'���|��'B;� yK7F ^ d@�>�M�']7fρJ7T�a3=����3�`���� �
/�C��9rFF�!7l]��cu_iV?�A����]��(�R_��?_7eE���d�z#'o.�0,v�hD��~�3y��)�ǻw���?���j����=9<ڧ-Hwܕ]ݜc#;������h��緜��O�w�����������~���Q=��\3LUvWť�t��r0�Uc��~��Fxv5����G�1�ӘU $וU��[�Z�N�v���,5&�' � ��n���ťnf���{*
�	� �T�6�}� � ��F&z�G�� �l  C�^��^�����W1���i8_j�z����{j �	A\���mG������Z�;7��l�I3�B�y�����G�ʙ�'H���'T+�W���	Jtu<�[z�WT�@%d!�A4T`��&��U�VG�1/�A�|c�$�o�?��@F�J" �6�Jj�׭��JC2��lb�C��iF�K�[Ϻ�*I$_�U݈��! ���rnP�[6f�B������Z%vC���b�r�J�ÕT��1�U��������,�*
���` $��]B��]a*��i���c�q�O���e�@�g7Ka*'��oV3�@]4���tw�z��M_���#��z�@e~@k�� t@H�����������F�UO��W��{`�1����અ���-p>�{U<]����[Ŝ`�y�2���@��wmU��9�nǀ��H�]G� |�Ŗ����ދm4+:��<��
�|ur5E��?1(�y� I�n�j\���=��a�!cä���-��=�הg��M�K\�P�,�pL���Т�,���h<ã��ކ�++��:1uD�?*�||d�M_�j3z�ê�4�ֲ4�eL����_����U��aF@�#�@�ҮeW�]�r���J��Z����u�E����Ь?;�Uљ�m�=�d�М�j07He!��9$4����,ǄUމٔ�+�.m���AF��"���>{��������~��cVS�fZq����řU�gg�m��IȠڼ.Z�B����ZM/���8�o�^ �(���7�v8&��odz~���P0�(|��v�����_w���Z-V�.�N�dP��HJF�3���%�&���2G��>ˏ�L�p;�Nb��o�ْ�*�]�W���?�GC��z�����/�3�ܽs(�|�|�}�k����8ޡrr<��t=��ܗߒo�=�\"}��pG�w�rz~&��Q,��,II��R��ĝ-�Sɋ�v`	�iG���c���,��6�%�~M	K�B��moo1�b�����sv����yio����$P��
ϒH���c*L9x~@�x��|��r~���Xm�J�v꼦�lڠ�5�\��]"�c�����m���H>x�=��?��ݹ'o=z_��ۼ��%C�>��O^�_~)��}�<�g�T�fik����+}6c,�=�Ѣ�9�0Rsɰq��˺���,_k�	��|�`Q�,��()�������gl������=8-����=��>���cg�q�v��t$HY1;�჻|fBq�ը���jW�X+`>m��^ήd�/�V�zDL95ȣ�1�7�����X���1UHd�M�D�| -8! ��io��2��$�ʆk{T(8���r���� �cPf)�#�nż����3��Ɣ�k������?6m�6m�~�mC�lڦmڦm��t7�ak���ؑnn>��y��-V�YE�p��j:��c���Q�YIX{�#�P�z�������\����3y����s��Zl�������7����3�n��5˴��v�j=T,�>+�m�b��M֐ (#��Z�.&���_P��* /^� 0ۉ���4 p��1�"�ܽ+{��aǴ3ܦ*�	����|1�R���;����Q���+99>�� ��Q�=��n�G[�ĺ�[��uC�pO05;���3��p�8�� ��ݰ�٪�+�{����sf���}���SDn������
�B�nN �lވW6^U���(�X:������a���ɏ%�2fR�ծ�	� ` �R$TB��na�3���
�
�1��[0 H[㎼��-�������?��g���^T����t:#�0�k�5�����lܒ!!p;����n���I2	U0��^�T��iq�YE{e��P��� ���(
�[ ����"�^�c1���BVd�q_��ʬf8jA U��h��@5)�%���x6�F/�8D_v <8\G�9Y v�þ��d��y\���}����lI2���X�	CS��X4,��7 '@�mP$ikp�/�#���ثe�o�=�2 ���.���[�V�!�Ԋ�����ˠ���ɱ<��[�wT�Z�lb�����x�~�w�ِ5�_Á�i�FE<τy�>�Q�[���B&KoY��W�7m𭁷F ��y��1K9#7rZ��'L �ZPu�����N��l"��kk�N�P��~�[n�}�*V��J�f�A��}T��3"�� ҆���5�o���~.Q��(��1W �[���-����ܢ�nC|q~8_��jO�VB�����5�d���A�@���ji�_�y��4�� �0C̭�[�q��SS�5,�����e��n�xn����Y]y^@"Y�\�p���=�[-v�@ڗ!���>,j�x�z��+�:?#�SCI�Rā1�˲4"/T��ۈ��)���lF�x |�C�ϖݓ��*�{��#@p<�i�(6_զ�QVL&7:uݞ�UD����) �s��j��
�2�����t�Y�塺�e%���ra�J섞�?������+�<}q!�׿���wX3Pi��~�h8���BW��]|��T�=w����Ze��q�
"���4�^��؉u�I�DT�u�,Y�f��{���%��^�}��<�ϑ��8�_�1ͦ{�����6U�X�!� 7�c��m���W�?�
��^��S_�x.��� ��cFRc��J��#����ە�ܗ��]����~;Ե�}9��CA
�X1��*T@����Lt��gUb$!Dz/r����.�cS�A�WG���,&+�Tp;�s�4n��v��;|lG�b}�u�k�2Pܿ���2��zS�ɹ+��'�t;�ٖ%�	�I�n�oN�����ܿw�k���eM���X@_
�r~~��=���K_E$I�]$?ˍ�҇�hmc�i2���钹%���p�~��wd�+Y�4��:���
��Fd���;������gzM����L'�c��P/�n��}]�ݹw�
j���+�X���&
nS7m�6m�6��6Ȧmڦmڦ�A[.��![JwP��?�H~����;���&o�\����m��\���72܄�f�k�F�|o����|��'��'_�W_}-��I��bXՉ�����lo���x�Mp�$�l6=)���E ���V΢�2�^�<ē�*W�Q����A�݈cC:ζ	� �o��hgG�tc~���	f�[n�У��x(�'o��?������������� Ȏ�2��B�X�a���]���H^x>����MP)6���#"�=FZخ�I�|q#���%ɗ����ُ�~�6��$GV�ܓ�Ɍ��k�~$ ��l�ܮ���n��}�iS0��24�aU-*g�k��S��"7 #@l橦���]�� 8���BZ�M�ȭ�
V�V�Wy��	I��f?,$G�|ݑ�|AeQ7p\��B%+� �<�v�8�lc�,�j'
��(��,Bj��	/HL�sZZ�B� bX<�@6�8Y��`xG�+����N�z�r��.lj�΢i���^H�/P�TPd����	���������=m�פ��Rz��^�O�E��7�Y1��0���a�����)*�7���}75 W|���Z*"V݇�ma���w/�0u{ ��{�%��-Fx� �a5����cS?���o���B~��_�Z�]�tn@��8_;Y�y�ಫ$"�u1-����@�O�؎;�{�$"�� �r9���*2;@���w`�"~Ϥ�-�1#?�� �g�J!e^<��lŨ�hH9!aY��ܘ�{R���[L�!��Pe�So���N���M���J\��XvKyC��c�1��Ŀ'65���}WN��~�ܑ[�`�.6O8���&�w�� �H�ډ��X��f�^`�3K���,�W(�`��y�׵�4�;ir���l��w��ʞ�mQ��r�����HK��>����P�y��jOx�d���bmaޞ�B+.(L���][i����
��ѯ�U�������!I�%I�,��j�R4fK�T�d��);~]%nӃ\�.d����+1�ľ+��;�_ -*���ڣ�Y��;÷�L�칏�W�r�������nqRϩ �ɜ�<P�F~�l��x���P�g��ť<y�\N���9�'!���`G������w/O�Ͼ����ɓ����S�YPѭ�YEV�|�熡�,�*���g @,��u�cH��}�X�����YU�3�\]����Z��2s_�>;��2n1����&�wUR��	���K9=}-�^?�)�P�EOV�e;n��*��-a-($n���
���ј�($���̑v}LME���l2���S��\��E��*	cͻ-�Ine���J1�d��a�'���tµ��穀n�e`M�����y6��ҵ�>�����g(X�y�^��l�h1;��u�
���cy}�������C����l.��N���������3f�wL��.r�*X\���-ǊykzVP0���t��2[/-���)�2+��.�dc!Pw^�b�ˣ��5U�U���ե)V�{��e.K#P�|�ɧ��?�s���!���椦����f����M۴M۴M����i��i��iT�����ރ��ɽ���BEH���7���3�d噁� ��w�����ql �� �;��b��[���\����C��Z���G6>�r#�Jp�v| ֺY���=��ba�B�!-k��BE|V9�.(Pnz�d.�5�.���҃���������޾l�����
!�V+~����W_��������'g'��`�1P���0���Tt�k�^�2&��L	 �#P���s<n��YasyHx�n������V��? �T�Y{�5?fpy&} zl��T֞��Q�GUp� aV�Ƅ4���B �`P��a�NSOTV�[�#�<S�Ǳ��������fy: ^f�T$* ��G�T��z��Я����;�>ұy-���2�/	��Bᶳ�B�a*��.��]Ç����>�!u�{�J��AcA�<X�t,��O�֍��D�������5�(���T��I �6Sڇ���������Z�V2.S� ܃\Pp�f�Ѳ�A�d6� S�Щ��e|�o@�ʳ ���P��q9���h	U$>�_�=�����V�7�!�w�̪i�w��բ%�Z#��]�n�kܿ�,"H��}�sD� �;&��)Ui��p�_�����/t��t!}�/q�P���(�{�s�ցd�eSӒJ�B�w���[݄�J��pP_𳭬G���[��ݚ �{> �;�sNN���iZCY/��M�� �#��rW4�,㜑A�a�=�!vC8�y�" �vnҞ'þ��;
@��7��k�7#/K'
��\s��[Ҡa�n��]����(.Ak��G �a�=ȏ�������屩�	�>�,�H�7�`�oB���{$#�:�F�GS8���d}4vnM�|�X��	A��CN���"�b�EU���I����u��9_��R��P^��0�=3"2b��lO`��j
,�F�\s�`�h,{��}�ĝ_�����bq��In�������J�F�B�U��<�!^�>(Pp�Y�.F��|�vк ��L�	�# >�m �rQ'�[��S~�٧�,9;Y��PM
{G(bA��K99��g��?l�:�9���_�u�>~��������c����`���

�Kp<\ok>�� ���-��;��1�}��;i���Oq"?v�� �}��ҲuEl_�� <��v8�fj��Q(9�|�0�Ra�b�+*ꐷan�����v�2;
SD�9@~��>�!�u=w�2B�!w&v	��C�
��pO����5����;�{�D��_[1H<6�+1Z�Ɨ�]QT��
�����Ċ7Ѕ�!�}����.'r��~0т�T��^������SR�b��C��)�Qr~1�o?���]�ֵp'�q]���w��z��sA"d2Ǻb��RFESW�٠7��ֱ�گ;;;|N�IF�Ү�>��j&o�Yxv��$֛K�Va从�-u���m�8���c�0f�9�Go��뵻��u����aOV���t�5ޑO>�D>��Oeo�@_�@x3����y����1�O@��� ��i��i?�!@6m�6m�6폦�Y�-j�э9|����X�����S���s�y��KV��f�i;a��#nfx�=G�p���1@ ��X��f%u-��n�vF�@(>??#�h�@�df���,6�P'�2 /T��<���U���L�%�~�P7���Kd�b �PH�BKh����֎���dgw�� �.bNB.;Á�y�ͷ�7���#�������5�.Yb��� w._G�s���8]�$��_GkV�]�������"� .������*㱉/��}�C%-
 [�#�����mr=c�w�F^D��h�G=V�"�v[7��Gp�B�6� \�~	���U�(�=��%O^,�7웊'��� ;�]��]��L�X�i��'fe�df?��um�ѵۡ��@�&<���B�>�V�zx_>|(�gW��ű̧K�-ҋ��O�S���B��ٯ�b=�@��O�/*���3P~]�	t�G~��yl���AX8�9�KZd����l����WW���\��b ׫��j{f[A�
�h쀍���2@d���x�Һ����6� ����.<�H��:
�e9�laRH���^ͥX�����7��+����Rc0�r���З��q�	���e�B!�s�A��=@��	�c�b�G8����F�	x��J����� ��k*# 4ϧ�2վ�ʹmgG�yE���u( ���BWc�T��q՞�S9���Z��Jl�c �H2أ]Xӂ��	��%V*�6(H�+������R#��@2������l�Kl�Y���(u�	<���iI���1ns9u
�cÕߏ�l���*�K������߫���]TAԦ�h	�2Ȯ�q��A��Xe*(�!�Q1�=֠�I�f$�����S"7ʊ�����Y��Bz��A<B�q;v. �I��'7�'��bs"	����}����"m�
����l�_0T����U!���UbjB^7W�F�Dk����T�xJ�����@���m���"�:��c
�
�P1��Q ����{��r\�2h-aέ�y��HGsG�=��l|�@c�5�� ��p����r�#�^�e#�БNlk��N�3��,�@��N��~$Q�Vf1T�K�I��
�^�Ղ*�m�� )XBv�Y���|�sO�1yu5��o�d:;g�j���T�𾏩6�ňS�wP|��s�-�F���T.�.I:Ž��cA�	2����s�:��5�*�!�����3/`7e>H2ޢQ�4K����if�%�{�F�o��@J��
Қ���>d���=�+7%�ѝ��ٵ�1�af����,���a �x�1/�5�}y���I҄�эJ	
��v��0�	�B��t̉��ޜ
_ڵUAi���r"�>{Ƭ6�z0?߹GדCf��@)��$��"�j�[>_�|z��(��R� �Ɋ�=��Ջ�K�Lf�y��p�%[:��=]�鵂-������vYl�	�W����s���������l8=\[ܗ�ވYXg�:ΰn����ׯu/��߹����Jt�q���w\����g8�\�''gT�9<<Ծ�b����d�ޥ��w������>���,���i޴M۴M۴\� ��i��i���m �<��o�m`ͣ��`��MZ������ى̮/�3q~.oN�P�%��u����C��ts���A_�@��fMG���F�J?�J7�$*.�ֺioo��m�`3���1��d� 	 <F#n軙�Ū   R1ڕ��}}�ǅ?EL��LX@t�����P'b��H7��z������?������S�) n:��;;���9�Ӂ�i�U}En�nǪE$@_��Ge܈vH�P��fN�d�@�=T(���y�˂dѺ�_��ot�|%���-sl�1_^K�^�y�HeJ�}"^���L$���;�n�b*��$����2%�v�O?��^�{�5�� i]���	����ai��1r'T�7~Ū�$�2�&�5ڑ�^yvM�aooGvw���H�*h��r��@�󖫘�_c��@ѠРG}�a%<��t��&������ h��L��Z��J�e��ec���$v%E�� 3lЫP���_�w�ͦs�����|����{�t<��0��!i���ʑ�`���Ƀ��cxW8����eEg�7r��}�{�nkI7�Ox�K���[�GB���c��WP��|��AAa9*A�ф�ڇ�H8 �qBd�Z���׆Ib��	���!��"os(p�����-� ����PG���-�����$d�h�o��Vm�?�Ĭ������㳬�Ȭ�,��Id�߸�µd��[�P-Bҧ ���8��J�H�X޸̀a�4Ǒ�qc�l�C7%�S(�y��Y�*����nX���O��f�e�悪��efH���"�7�쑄2��l�*'J�%���b�)nI���47VS7���+���V��+�����­ c�A�+I��9p�N�$'M1N���8�ݞ�y;�CHw��FAo�o)?�6O�>K<�#n-~��S���x��=��E!H�*����g�)��\�Hԣ� �Wb����%*�^|͖�J���Rdv���j�a�9�Ū"1�t�2���bR�T���*��Oh�%�_R��'���N 6x�o��I���+np�(X9�R���mɲ4q�9qB2�򛲔�/��汌�De�>:��$;��x)s}�e�%RԖ��̦�z!�'��]9�ŉ�?X��9���j�� �/�g ��(�����B��u^�ul�Ğ��o�p��\(ކ�6��k�R�UP��uJqdP�v=�f,���uL���p�.�g:�G8G�C;��&7k�������ޓL�\$'�<0�"�8H��,1��>g@����k�g�@O���Ç�>۱��q����f����xv���"��FMi����aj���AiM�� ���7�����'w����Z�M�rD��t�cA�W/gSiVV�p�������/���+^o\#��-$���=��QmA�(��uH%�[7��ʉ�k�^?���sy��y����3�k=̧$:9c4�΂�gv-/^��o��J��'&����G挞x��wx�����{ҕ#=ރ�����ދ(����b��r�f]���B;}�s�sŭ��M۴M۴M����i��i��i4����U|B�?_.�����/B<D��0�1Ň�IKY]Z0������u�Ob O����A���ġ�=yQ�� =��G�<6��S�ek4��WWJz��$@��X̗T_  !��x��0T)f/sC��3��nǰ`�j���F|�!������ z.�d*����_��oi_��M�3���
�$`΅��8l>2�.�~����V膊l}?�l��N�yG#8z����Y��V �����Z�ӎ	 U�p���6��}�v����^��[����"d�7�sy#�1��1n������R^�xL0��]	��A4-%�͓)q,{"b�8^��@$�[@r�N����G����l͍�ݻw���<�˫���T&������B����K��H��%��l�v
��%_�[���bf��Wrvq)��gT���2ж��=������-�\��mVs+j���ʆ��"93gP-��{X��t&���-� ��yCuS��p�)tI�\�2��RT� ��>� ~h����WeJ�:�pk\j�	=���	���w�+��G2HX��ݰ#���Of��Œה�Gl���b���[3������[/�S!���#�8km�X-^�Y�k�7Yl�=TW��BVj�ZFVO�Z��@�Q�V����n5�VvoVpAp+ׁ�
� -�"��v倩;�e����&�n��y\I�ϼ\;'?n[p��RӒ0>�|=��L��S D�iX�����+�������Z5�W@S��d@�������vB%�MI�R�5b�� {��"�_��'���r��9�+`TK��<7U������\�Ն�'�ف�0�5����Q���M�G���f�7i��-3��DK�}��$oi�v$����ꆈ�����W#Y8&�W�g�.9���
U�R!� �-@�)X�&(�ă���xzf���2��2%l\3�9 �� �eN
��J�������5�!\$�u��o}3撠"�L�HLr�2*#3��c�k���ڷ��>��cT	��p �%�Z�(�1ش�ej$I !����s^��ۮ�tH���������O���W��ﳸ㲬`ǘp�ʗK9׵B�z�Qxc��}3�MX}���K�{�V�*�\�:�0�9��mf�Y�En7�<����be֎����m#�m�B�XŹ����� {�>߃~�����v�|���_�U�T�-�zlk(`�
卐����X���B��}�<��j�J1��,6�j�l8钩�yp�'o��6�X�4>�w������UF�CN{���U᤻yEޚ;t����W��7x�t2��>���ч1ɫ|ɜ0���a#����H��`0����>��Һ6^-[���?���LF�;�{t ���|��EeF5�DX���ϒ���^?ձ9�/�������W�'1,t,��cKT_��BV��㋗��o;`!�荼G+-��A��~�-X��{ Kz<���i��TpM�&�����_WQ�`�>���WW|��i�mڦmڦ�`ۆ ٴM۴M۴?h� �`�7V��F�7R��*{S�RX,$��٘
��l � %��>�'Q96�O$��0<�!��	���:����'�����*���NY�������p��q�����e%d���Ol2�8���z��t� l�aG 6�+T6LĆ��A�����ψ�9�_����o��>��4��C7��C�_^�R7��y��-9;��}G�6D	`K�����3{�f��)�� +r;
^��,F����2����`�6��h�U���ܲb`	:�J�����WV�R��Jn�C�s�jb�WL{/+G�^pk�V�y��=}]$o^?�f�O�;�J*���q0�SMy�Q�@Xz��mMb?����ѝCnĿ��s��o~)דk����%XB����>U�Y[�欰��(�Z�a�eM�����8PD`�LF����1�����Z�RQb����� '��׏�T� �U}^�
d�ܜ{���c���H&V������!�>a����Y����4�LyM�[cI�=����� ��o��V$�4)ֹ��]ൊ_�P��sY��,�Aň��в!���K�dW}��$)�@s�)���LX!�T�.!�'6&�ц�@�J�cf@��k��+R���sD����s=Y�N��An4T^�-��u;� �}��k���[�<��p#��m��`_Sz�����"�l�X��P�n�r/���?g�� t&>T1߇����M�6�[hE��m�s#Y�[6^1-��;B�����"��읬�����ثu�'(<?�8����m��m>H�UĉU$��ĳ2�:�-��yޒ�w�Y��F�c�bV�7�����i��ʈ���}�Z��{�U�$�ݔٳ�x���p�2X��3�KbץA�<7��y��\��]���	��1��\B;�m�(��6����q����-��F�}W`b��b X�����S�89l�2�7���e^U��p����\-Pڽ�К� Acc�Ə)�q� k��v ��0��� ���H�bahz�f7Y։)n`ɷ���)���xd�WTZ�U;ۦ�����3cֺ~�|��A@�˿���Ӛ�l�0ΐK����ɩ\��!Lb�����K����m����q~~~nV�z����(�ә$V��1�e{_��f��&F�Q�B�h�`(]���#r �!���<�e%˸��l;�vL��֦P)� �����Z5ba��g��2�øc�)���qeC�VX$��^@�D]��)��v-�gBa� �-[ŝ�=ڮ�c�Ġ6d� ��pG��2f�q���{�t«���7�|�(�x��|��Ⱥ���l9�������$�3��r&��ﰼ�37c�2׸V ��9�����*�wܻX�޹w_m��i��HI��J�U�~���޺��ʋ����ou�2�>�&�y�9*+ܧ+�ߗ�����R���kS�� ��ߑ�C�#�"(�A�b��5����\Y!�:�c���~���U�|��Q�̾��������W�i��i��i?ض!@6m�6m�6��PZ!�<5k�D�*z('@8>�'�=���/�|"�k���)fSY�g�\3��ރ�T��f�8�}�s�{&6�u)��n$��e{�-k���W�����f�
�-'��҂�Q9��t�uCϑO5J��ǭ�7����W�V$�O���B��Ƿ��-��� 9xy��������O~�f9d��̣o6�x"Z��n�*�uS�&W ��n0a�u���
P�$QJ����˅~޸ͤ0k��̡�X����To�X��T��v	�M�����@�hv%q�,���u@�h����- �����;���|���^	��6��ױ�C�Z�5
��I~�H���d�zy�n*�ᖞOW7� ���f�҅��#^qi� ��N�� ����4���xA��N�ɳ����2�����%	�c��	`��_}��C����y���C�����{�$�$Y��gח�#\�Ir� �4���������(W�j��򠄊���%���h��	�
�جL���{��a�Y�{-T�|��$����ȃ��4֮���&�m� p�5����i+�[���\`	�p�ͨTyY��k<$���0��������b�Ѿ�efmU� �`mE[��k�cm��U��(P������%8��`kƱ��×D?խ �a/C�DbV<����'��.N�JI?`�r�2;f'Դ~�2�db�m�xc&< �p?0 5�� N"*�\���
��	#bP=<��,�����ALG��D5�1�H��@4����R)=_�AoW�������,�>v�3�Q� D.mn�<S5f�GeYb��J���"�m�cB���ז�D2�	�EX�^G�9�lX�b��	"g���<�iڪC���FҪ����MZ�>�V~�E�����D����Y�����N�H�}�1�[�wB�u^[�,D��_ސQ��Wn��z��n6vLq�>��`YP��P��9�e�
(jǣ���F���L���Z���V�͟fud�0��F�'����\��9����	��,i�:���8ul�y�yD-�:fQ$������L���qXIF�����ç�c�=ˇ�j�[������T-�= ����7K�6W�b���d��HBE�����~��֟�3���t�������ݕw�y��)���lMR�;�ɾ� 9�+�E�������	��^&A��b����+�<�[�{�x�c�M��ƳyS�����i��g���#Gw����� ?V�I���b�Y� �3��ȼu,��jq��",��0��;�5�ņEe6X	CC8��gKZI޹����%�6W�t��|��\�vuPS��1��k�&a��\��4��8>c>�c/�0����i�ԍ�A���uU��$����#g�t����\~���p�����A*c]}���3jX��ׯ8N<P�3��H�w�^�F {}���ء�@W�7�)�(��̎-r�T�X�!ϭ����X�vu=}"���g������Xת(`Y�ʁ��ѵh��
�?�-[ۉ�o��1�,g9}��=\[��㑩��:`c�Q���}y~�|d�a=�3������O�m�~�~���b�u�ZGQ���ڴM۴M����i��i��i��y[�H0,�͝��[E�H7R��n��ȋ��R7�덶�^֥�~��=n�稺�׺��e�"�:��i� +��r�>�fG` ���Ќry��ǁ1@k�P3�<n��H�kIa���el\�M�!xm��a��H�QH��wAi�Ү˕�]���h�����B���A~�ӟ��c�/�EY��F���Sa�{%m7�v3:�����>��S��u��Q�o�� ʚ�Upq0�`t--E"�:��p�`�؈� �Bȷ����Mu���JV|�V�6 MӶ�����K��_��{��q@����D7��k�.�z�8��Z{�sG,��ce�!�B�i6/~�6�`;`��
TCUS,=�3�M��ܹs$G���ֈ�2 > B��U�@'��%+tae���S�sx��م\_]�8#V@ش�b�'��$@T:�Ƞ�Tid	."��t�+n��I�m�Tc�\Q��V�Z��=^�:dw��zVr�W�Zޅ��� �0����XY�q2�C�=���_�P6[V����OY��h���+ia�ؚ��A��-7�;0P	�]R������b��)`�b���j8�p$�+�g���`����N�lt��N�����½f�r�6k+����n#�ĭ�
������@��T����1���*W(���m�ĭ���|,������E�6��YŎ~�M\�xжkԘ� �AP��
O<��f
��m�"��q�5�J�s~<X��-������s �J��>NB�����,�*'0�ĔiTm��0'�t�R�� �B�ZYx�ߓ�%�_���K{+����]��G���[�zh;�?��ܼ�}�����	�1n�7���6X�k:yg��Wm�|A�̗'t�+��V��U�,-$�����b�G	�)e����x�{CM�A9srfW���^�
�Ǩ�AbI-��_�|Y^MB21���{�fI�3;��1�xc��ceV����`[�ݤh-�jGnh�%��7�i�����d&3ɴ�i�+.(�ij�e�4�j U�U�Y9��o�x/f�t����Y Ii�x���"<ܯ_w����c�MUDE�>HF�}�K�uM�6����*�,��ͫ�J�����+�?��}ZƓY����ccMz�B�Hok�ii�9���l�l�g�=no�p�-�NW��Þ�=�a��/K�����M�A1�Af��K�ت�̴`D���	�$r� u7�JG5؏���l�s�����uBR*7 � �qW�\�*��53n"w<Pm"�{k�����'�JԊR�P�D�b��wߕ�>�������C�-Y�8��)2� ��X�\_� ao���c���3Y��u�����U�g5���!i��V �1�����"���h���a�OSf��QK74��po�#�8�,0[�B�z)X��b�Z��W�+9�3y�����BQE�����-��q^p}���c�VѮ+�=%���U��@��@�ˍ�CcN	�9�%���*3���[=�|_ɳg��?��|��c�ݸ�Q��2�I4�:���_w�n���$��#��L���K�{]��Iv[�>�?������wY45����J�ێ�����ԝ��$y���D��w�Ϳ��76uVMkZӚִ��� MkZӚִ߈�2W�$* p6WXD��Uz���CY�E(*�`ˀJTT��~�8=����jI+���=	��p?P��]\��-��R�(A	����5Ԅ���9:>a`����A�c�~��wu�_����C������� h�2۝V�%� 
w[qB�H���Ɋ��a�m�mˏ~�C��?�S��_�%A�����-�F�c�����l�\���rtAu�r1_������ˋgGn!����<�	��� ���vvٯ�~D�������n�j`t3� �"�b��3���-�w�ͦK�n��� @|0/��ˌLw6rT@_}Tx�&''�Ӄ�bw�-��q��ΰ� �RHd���Ui <���W��@%ni r�ռ�ྡ��x��Η�rs��N�/���r��}.���1�/H$�)����gr����Ne��(,r��X�kF�Y�j9����z(+��w< =�{ a@~,�7S��G,���l>uc�T˲��5�Տ�3�4�
Q���}{����Raė�Z�^T�Z4��~��#���,�I�u0<�)�bҜ$�q)��aY֠{!�
_���!����4���X���DA* ���3(��$@Z��U� Q3�2�Pj <�NT��C�i� ��Mp!i��T �����#]�a�cć���;�� [�!�gRu�s�"8�Z��x��{ZU<>f�-ՆR!\���v@z��A@̟�P�����2L<��?�}/KS�ĵWT�5��"Ckj���$!H�5֧�cY=�PA�âQ}_l���������!�b
�0��`V�z�Ǧ���;J���}���-��6\��1�bT+ZȻm�k߬	f;���UU��>���5!#,�ze�ɏu��^����?�<�EY�*��׏	%�ۤ&��	P���Y:iފ��aD�u�N�?>��z����T�\*iWy�lj<1u3�+f��ZoA)��0l찍!��/T�-��n1���kJ�MUSzr++�*,A���Ͷ~�ږ��_!��:7�w}hk��C+�L�*����*I�2�=��?"���zkk[��yʏݝ}�/�s�͝�����'��#�����W�@R���LC�A
yI �E��K�aҰ\��Nx��u�7�1�G�+}~vX����D�5 ���'��#������B����tOX<�}�W�3�r7��#?�Zy$a*��@����/?�Ѯ<{��}n��^���ba�4�u���k�g����1�-�dt�
���8X@%-S��
H�#y�ֈF�Vv��&F:�k��@M�,�H��Ɔ��*�U�\Ǎ��i�ތ����l�+C6�;����s��Vդ�Ĵꄊy���z2��D��R=Gi�mC���SG<P\�a붳��ݟ|��\�NS���Q�r���������g}$��'Ҋ:��ye�t��/�y�*cf�<�ۻn_P8b6�n�Am����_<eF
�����v�<���m��C7�FT��ܟ��K^��Q�U_§S^�r����K���7HӚִ����� iZӚִ���[i��q�be`�-�..����]��X���u���E,�d�;�0v�4n�G��d>��ci[�y����=��xą+?{n����t�DBe��-G�Wr������Ç+�;na9v���!+��X���PhFQy��ԶW���n��qҒ�,�[��죟����������>��߹/w�ߓ�ф� $`�E�����s��B`Y���ߐ[{��?ϙU��M�gK.va��$Z������ՂZ�]FV�_)ȸY��*�ļ��4�no ����8���+�E����Z�!*��A>Fi�|? |h�1�!Xx����(9��7Z�_�Y-KY�s�E�<A�%�b�oq8��}����Ev�>l��ȝ��s�0���ĉ���Tn�:$����n�y
���ޗ(ݹ:fe*T��ʘ�1��U�@`��DZ���9�{P���m���G�K��������$ �P�y���j�g��s��a*IIۀ��X������a�C�C%�,Ԗ��>�U!�5��������ze���3[�7�㴿��A�UX�0��&H$��
PKk��Z�����Xa~���Z~	���8#��Y`Z\���# v���?�C�F+0�5��;�f-f��8]�X���J�|���*�2����j/T�
|ͪ�u��}���,Sp<��V)����
�b�@��� �Օ�R�s�OR�q�y�TVE�<�~�qW)��C�7���}�_�6o�4@�tQ]PL�4	S�����3�*e˫ ��+����HցD�i��}/H�������_�`u��gU4��CU��8�R�	�Pf��9��㕊�:Wh#�(j��)�����#�b�X�,��a���R�$�?��\2�%q�Mi`�'�"Y�w4<�p^�bmI�ZBf����A=�<��
�}jD�~��p��.����bz�Uo����E�J�l�
#Z�2OR�
�0PZ�r�qep4+�qM�*��3:i�sUY��ΐr��.�Ɛd8-���Z�e"I���	�z[��l\$ՠ�K�)�e�dF��`{8��K�c�<�dU'����mq������}Zr �}Խ;����=y��Sεx��cZ���lw,�g���TaVJ]m��S�-grtrL����ۡ͢�������yA�l�:�T���{>ޒm���E�d>�,,���=�?��l"����\�8<@��{vw�|�2���P����n�뮽�B�(b}��z-����\l6r����?P�>z���<��/�C��`����_��cy���T���D266aU�P�b��?'��eD2�*�og�}@���S���/��v�G�6r��9�9�o#
ǆk�.�:�sG�Ab/�����C�Ȯ��=ڠ��b�M�%lE]�y�s��ͻ����'�������=7/��$h�r��� @��B��n��ma�*>B��'�jaFR��B��Kf��`	;���7G�<��VΛ� cqRK�:rf��Z��G7�哑;c7G�%Q�IӚִ�5�5HӚִ�5��ۀ�I$C1VQ0�p6�a��|o�0T{4����d�K1Bے��t��z��`��!�,�Vsx��\ء����B�Gc�
��L�6���!�y{kG��WnQ5&&U��ޮ����-֡FA��N��Ih}R�W�?6�4�B�g"�? �d�t�P��my=�'�?���˿�?��?��?&!���C��R�n�l	�D�Э���_c`�t:�����|�{�7�������j=��.�{,AL$�ZQ���w��Lq���7J���(Tp�.����ZY=xA�]�"�y�{��ﴃI۴�H[ꅽ�|�.���@���~�j�D�~�k��"CX�LNO�Hn G�eU��P�\"�٭�[`��Kzrs��{�,w��"�(�/ڟ�:�h���#Apvz!?���IhM@���>�ޒ�k�s�}��w���?�������?����ry>�j4�j��g���r�Ln)�����c��;[�U�h-7헼M����ȪXby����*Rk#��$4~��Tdk܅�V[���EX����5��'-7���Y�`��\�oV0����ri��rX
V�V_���6��?�Fԥ� i	U�u�;ъ�%�SU*��D@3�˱V�G����J� ��@�(jARЧ]1d�|�i��ܷJk��{6p����V짚�`�l�b�Mؔ���}u�'�0��c�w��u北���`Fr�+�`��7uAH0ZC�c��swN�y��64~��9���lf��d���[�[y�ـA�To��G�[�� ���Ã�̰�Ⱥ(,���	 ǖ���l�ձ�'�ݡ�P|T���y``�m��&ѡ�X��**B�X�w�R��i�F�Ǝ���^��>��&�@y�U�>��4��W��~�+�*�2/Jtܾ�����W�i(��1�$�3 �P�&J #�q�{F����*�rGHv1W�E *�y�Q��<�^�� �}ވل���.U1.T��)�R�����]j�� u�{,�-����sAWU�x�$�Ӕ�B%��j�1([Ϭ� j�%���F��Z�s�=F���)�I��IiE �>�d�Hǀ�A������F��n���M�y�rW�w�d����rSm���>�1���H�X��Ҡ� c�rkp�!L~2�H�C�F$�+�/Ar�bQm-1��xE������RՒqJ���ŕ\]]� sU�:=���AF��X0u�d�;����rjԦ)�̖�{^B�K��gjL�l`ݠR/��d������x���I<������T8`�P�"S�Ý!���XXn��� :�5Y�Z�jC	�<�Z*,s�v��/+&n�6�-��0e6��f}�$<6�U��^��%�$b2�jI���w�� )��.�������˼�Ϣʺ�6f��?�"*�2�C@C9���jA8|��|�{ߓ��rz�F�3���E>$�q.�7n���@U�����#ͬr��n����C�os����]?��d���K#>"S#�ͺq��j|���d\e�U'��y�������KӚִ�5�5HӚִ�5�7�e�)��4
%[.��䔋��[{��ke^��J�O��Xڝ6��rN����n��-V�TЯ2����Ͼ��7Gr�P��g�d��lV�X��l�BA,�Q(zv:v��'�6�����gl��.�Ym�����Q�4Њ�U���#�p
[m���n�-[87y�䓙|��|��'���=��翐�O��q���Y�2�N\\��g �&�~ǻ�<���V3v��<z���ߐ��]9~���	���ci��0i���.��oN�.�0��z��E|i /�cmޣ�]B��ȂPC	��"AP�Jf�C�iQC�I��n ��;����?%���$�V���YQ ����`�>.ߜ�����U��7�_��A��Fa8�����j;���k���w��ruy�>7r����;�'�!�j{�&x��E-w����/��Y-
���Ϟ2���ϟ��յt�Cy������ߓ����߸�\ȢX��I�q��V]*8{`q�Z������&8�C����J�c�A�aZ_G ��׉8|�L��+��J[�pU� ��Y�5��K%hQS��U@A\[d��U���R�@�-�p  ������+��0phB��T���qf� yD�HXO!�<`~G"eT�� %m��l��������fZ(��!��lh�SYqUz�{ Z��:���������P�$밺�_Ty��X�9��QӔ*�����QE��}��RR�PaJ��u����5X��ľ���Z�d�6�B�\T�kE$�T=�4u�n>�����W�*?�*����'1@�H�p㸩|2;�Mr�	�� �W'xŌW�� *+Ñu����Qm�jl��lyn�͒-�Ǧ�݀B���}�c��*C��ޘ{���r��p��2�Wɯ�ш�C)7-μ+_���P�K�[��WJ�P���HS[�*M�
,�=d6Ѭ����	����?�>���H���Y�T�a�7R%��ف�1�,`ڮ��TI����%*2�	�CK9�~���z�V�ڄ|IP#��/� ���^d�)"���R_�2=�$L�!V��P�/T[X0�[d��R���W������
�>F+�P푼�}�	U�͒�ߗ�vQ���HZ�NJ�KH�NRm�@�C�����l*�{��:���+�DL��S������!![O U�AGU��T��G�������
J��
*l�N/���Ǉ�c�|�8��>`BKL��_��]J
�g�/��;�;��#���n�p��H��.Ip'��{l�y|��莹Ȼ^�-A���$72����ҝ�O�<�e��_��|��ߦu(�sPݝ^^ȹ�+�~�dK��<���;~�z�ϬR,�$A
�f	�K7ϭ����,���n��,��z�$��S�g��2�B��BX�';6��Xt/M�y��&�:�5�k9���<X���F�B�[�s��L��i�'F���!�3 ���"٘ɹ�g��G?����#���#ޣ�� �h���}a�bA�H�$�8+�4�J�*�<�t����,��� t^7U΢|���tڜ���]�>ha�Z��񍛻����e܊?sW���R���/N����{%MkZӚִ��� MkZӚִ߈v3Ik[}���S(t\�PaxW�r!
K+Q��r�-�4o4����q>�2�q:�v��Sy��K���?��ϟɒ�0�,`4JV�B	VA���2�M�b���OX�x�J�w���|����7oܢ��!�����肘Ѕ��x�V���L�\�s�2�����$>>��#y�ɧ����r3x�VNg3*a���0Q4�M�)�^���o�ʻ�E����[�]��l2'P��Od�к�-�Q�ز0v�u�C���4�4@ۃ�
_���%�b*jZ
�TU�E1>3r�e�|V��-�	@��i�����K�4 �`31�)�@a8�o�$���m�����sƅ��c��ppxW�w��)q��J�ޑ����mw5��?h3��~��o3 t�Du��[��K�u��5���b$�������������s�3�oߖ�]���q �Zd��,�5�<N���6#�WJH�$���U��{�vN �QY�	˨�4 ���	S[�ބCU�b�0�H�ᡅ�󲪔d�zP� �@je4+����ŵ�
tˇ����$	�Ɓ}WX[�h�Hh�
v^kNm�rw���MY[_��DɌ�!������Y t��/<�����B�xl��h�n����ֿǁ�����Pke�z�Ȥ��1��*T�8f��e�<���)
��Oߔ���u؏�Ѭ_�,l�HD�N@VYE�0����]�?b��؍���?5χvDP��(4�[T�/�ѷU�A�J$��iS�l��o( h�S�`~Z�)=HR��(РRF��^i�����,h�5a��p�HY�3O�DaM�辆ܗU�$8-��u��Z���ܠNGsB��=ғ�|�C�=�o�������J	�0
�{���T� ����ʍX$ߣ�$�&t(]�6^�V̦+��v?~��y�#��Xm���+2�`g��k?4�:q��̾i}���ϬT��\�@�S%m�*��al��ge�W%��LnP������/����c�ES�^�5Qmd�`&m�v�~%/Z�aDjw���+_�lQ�B	g��[Dz��N�f<H�(���5O]����r�����d��$
T)�d��['jŜ$��b w�\
Y!�vlY6%+��/�LE��~��~l�#�\�)��x�@�v�}�mqi�| ��:��v��TR��/��C9<���6H([��EU�^����ݜftz����Bfˑ;�r��R�?|������}�_���{��o�p��^�ʛ��$���pp	t}�~��/�]�ɵ��_�d<����P�n.���K99=��ՕdP}���9T6���ܶq���������ܔn� �B(�AT�c ����l��� �vH|�zJ#B~�!�����;��t%7�ȂY�f3wχ۷�����ͭR�	�D�]�҂-X$�a?1��w-�*��\&�k7�}*�}����?�ׯ_�c9�"� y �d�����ۿ굈�3��<����^oPv\��<�NY�T���85"%�+-D�HBq]�fun���O��y��L����ܐx��?�g��/f�O�x�������?��5�iMk�o}k��5�iMkگ�a��	s�xC��|&���;�Vn� ���ì���˪< &A��>L�YX.\]\ȹ[�>��K��O?�Ϟ�̼��Ȝ�բ'0���y���"H!ըƻ]�/>��VQ���b��^���*�����6-��H�"�X��]�d�3f@,ݢ�׿�����O?�˫-{ �V �s<�+�t��p��̲��D̃� � #���rN_���]*,��o��X�~@�E#�N�M �-��ݝ]H����}��V�Ӳ+�jX�Ю��T�EX�hE<�樲f��<�E����J���-r~xo {�r�����V���V]=w�P�TVE���l*�%�3���LF�k.��?�Gb
�訄���^����B�n�+�0�uF�@A�0� β��	,���� VT��|�̍'SS��t	.���
� v$h�B�Ƀ��|*	f�nq�� ��(<`�S1���,�	�<�9Q ے�V��>Lm���W+ڞ��"q�v	�K�����+
t�l�P���Z�̌�M�bY�*v�WDjsU���%��g���
�G�����h����i�p�o��O[/�)b�s�t�Y/�y��)���p���81���l�4���\��H�u�PAM����?G�/��Y��T<�!�� q��<�J	uL�mw�B������	=f�P�3H�4b@C�=)��/U=y��0
��/�4#j	��8Rɫ��XE�}�m�s8�*��	��!��&�����y{+H�<���Zê�9�@|U:�8��%��(-�@�j�]�+���؁�W��}v+�m�X1��>4eDd� �t���P�\Py��2�����N�����ʬ�d����b�G=J���8�j�� xޓ���}����2�8F���
,h<0����������K�*<S:���%PJ�h�=Sx�����}�WZ-�wj��t�I.����*^�Zl���rh�_�y��r��S�$!�A����M��(5ˈd�U���:T�2�ǡ&��H��2e�;�P�7De��Ia[�7l�bw��Bѫ�|�:�A���]�I����(���2"�f�*�aIB30�+�~+-8
��TbZ���~�?��,<_@<hx�Jrt	 ����A�`k���j�.@���дA���/|)
lv>���}g�3�Թ :o���혪(gI"�O� ��p??����Sy�w��ʘh��F�N��q�^�����DU8�������V�{���/����3Z�~�?���?��n�x���'��}g(''GB��پ�����L�_|,��ΟĠPX���r|��C��ᱛ��iӤ�+e���k�-gt�=�cf��<���ij���DJ�q?m��j�c�u(,8�r��P�,�����s��L��W9�����c&sͭ
�k7�8�5 �|��Q{Þ�����}�w{Z�� A�N�7wp��!T���������<{��͏F����G��7W�X-9�r7����f�YAT"n.7�%��dEP��n澳��7�]��<T��yL�"�5�	�w�x�M_����񨪂������_�{�g��5�GӚִ�� iZӚִ��F���M݂l0ܢ�Q�������\��F2���RA��c�%�<[	�V'Vs 7��[`O����PB, ��r�L�K s8��9S[����{��������l%��r��.-^�~)�A�rk{G�O����߳��/ۻC��PA�Ĭ� ���\�����ZF7c ���!� !`7���+�uR�cO�2������0߄Aݡ돱�"�����-�=�C�&��ѯחs��F_�V�����L*T}�cH�&)�������y@1<�����ϕ��G�;����ۥUV�� �w1��Er)���{}��啝� �G��,�E�]UI�,@� 0�rkQ	\eTh�N}��r��V�m��Ĕ뗙;Ox�jw��ݾ��u���V�t*'�7\pk�HD��QyV�X L\-F��z�;�<� �2�Ϥ݋%�2�����R���w|��~�xq��~����1����>-��*J�|s�yˁ�ނ���G��Q� +0T���vKE�~ 6+�~��JC_tN�����8�i :�`��<�iM�+�K5t��x��ǰY����1�S�PJo������E�Jn����@�8���x�����/Z�c]�
&���o "�A�K�����Б��%!��u��8� a��"Q#��|*i`�S��?���5��x�*v��K_�f�оK-D��(Cb��%8�@�i��fLp�y7ˌ�# ����=.٘��		GXo�ᯕ��%�@�#̵r>Pb`1_�<�6쭪0�+���b!
fdX&IX���KP�m��*5�<p�PA���*$2�X���3�*��Ŷ`=#*��=�vH�^X��ЈU��՚} 29'(��-�`1�x\̦��B���$�h��Q@`�.�hp�e���	X �_'?P����B�M��H�=�'���ٱ���)�9܇��5��>3� f"d��R"$W ꑀ�NJ^���d��	J��w�f�����Y�1��2%���8α\1���B\5�a�#�B�*�#�?������g	�j�Kn/5���dFD��j6(�@�#�!q�u�S(�M�	�O�\A=�)A�{�W!��#�(fr��=��0p_Ԛu������bL��A"'a�&�Ğ��ep`lE�~��C�E��7�5�A�t4r���M�n�nn��a���'�$��ޛp�Ӝ��V�z�
�0D��5�\�
V��[�ṕ`�����)���#���a�m�}�����	(Z�L�e0�ɝ{$/�̜/r�/�������Q��H���z%���ZI((q���}J Xb��8m:2��D���
3�w��>:�߁�h��h�� ��VF�o�8pc�߽�g��ŵ<y�ǻ��G���'"���2X��t��맟~"�;���mnu��@����'YLR��4[|>�8s����k�S�Vsޟb�r�qE.�m�1�>�wd{0tc�$��|/Z���B�$E�zK�Y+��}�E �b�+��|U��8�\� �zU�"�Y6�\��t�_���9�˕��Lr��n�������U���s�Yx�۲厫�9B��07�Ǔ�g ����Ky��9?��
n��(I�|������x���@�O�HZ��حP��
�����{����#���d��I9�m�?���`�N�7�#��}��������'R�/��?����σ"|���w�}C~4�iMk��Pk��5�iMkگ��:�fu.���\�������ə��=���"�+���#��S�Q �;na�� *,\w��g�P���v�]�3�OI�dd�,|Pd �G�#ȋ�[;r5:��sB�����f���_ɕ{���<�V�-��Ky�����n�?�����\]Ծ��;^���J�i���-�?8 �xqv)��SYe��,d��#}X?�~�Ogr�ǊB�z߱�Ӡ����h��kP�������\+Y�� Z��-�H�� T�FV:�=�I
�Ry��js��JЪ��d�N@�
RT���ר�e0}P0�vE�xEP �q���kd
�����?-IQL_� S@O|:8-���`�N�z�g��lO4�=b�2�!ʺ�w����dU�" �0ߪ��A�N&S��n�]�"��0�b�G�LÇ�����|��rS,+!��"��ʅ6f�� �>��y��$�l�C0��$��Œ���^�i��y�廡�����l��Ei���斅@�v:f����c����+�c#T���k@����3�L��D���sBг�U|��͜��Dh�U���:��¤�-ͱ�4����a��~(��XW��F��5۰��<��m�V�v� <s���U������c+��w��N"BÖ���݇�8�֙+��e-~l9> ۮ�"SO��f��WȔ�kR߆��1uW��?�z�+q����k���WrD�oU���V���o�T��"���������(,R�T��Y�&P��-���[��Υ���@e=�0�O�^Y.ŋO�Hs-���\��u�F����jj�<�ʷ��rǪ`���7x��S�yֶp�exF��`%�G6�N"{�`�2Ӿ`N
H�H�!�����UYg��N*0K.���2�2�,��)Ə����H�qD�����*kS��3J�w�����J��aTվn�Tj�UU~����+�J���Ƙ¸+k{&Ux����Vi!��PQ����K�:�byFU�~�vAM�`�a_��Z�_��X���H�����uCb%���{��ڦ��#��iV��r$�bZY(5H�n�ϥ4�<T�/f����L�U[B퉢	m/F�n�W�39n�0S��m ��~��ԤUH���rߋ�(Ɛ/Q,H_Ȼc����;���(-!��U|����V�p��">��P�En���;�"!����{�ݞ�yԝ��p��ŪS��)���ʏ�P��k���$��v��,���<�A�b����O��-��)�Y�D�~�v3��$�*g+�Ωڋ�������G=7gE�d���`,n�bN�G��H�@h!	�lPm�S�9�W�c�Xp�ȗ/���ͯNO�eJe����M�r�ד��?�X�J�o�'��]_��|���y9�\̸]X�������+>g{ݔJ��fנp`���x�t���k�2��Pdҡl������{���>t�{��KWH@�.��;G�������pஃi����"*��]ݻ�Ή�㝔ex%MkZӚִߩ� MkZӚִ_{����bn��s�F����:���z�Z���X�:��t�_�˹l���������ܖ�[����i/��ƭ������-���cV̢���r�.�P B-V�j6-dVKV�,��6�n��wd�־ܾ{_nȹ[@Bpv5���3�(k�:9;'�E�e����3Y D�&T��Q��,hA�~�m���]����_��}�H ��4e~��;�e���Ⱦ�>J#���A]]����	�nv[� ���3?�󓴭�6�/���@��� �5L�I]�����e���M('���-4[$��m*����/?60ZA�����#�w�ӽ�n@���%����W��dE5< x� ���|.T'w�$+��^�k�ͳ���䇷T�m+����mɠ�a�#�ǳ�-rt�]ڶ�$��I�rc�M���(�� Ђ<cb��lO߶:��v#���W�xk$ bK%����쏐 #�Ͷ[�Z�/ �� � 
�1��q�#�w�������K���B��C���$D=�\��բ�PX+��@��F�:��i���Q�#�<���W�Q�l��F�=���Dk�pML`_�&�Lyc�~>��,��o��fC�X����@Q\��{P��kp؏+f���d]T�2'�z�ϐ�|�J��[t��"�W�>��MR�7���e�?��B�cQm�U�Ǣ�Afk���u�{� �)�w08ܬ~������w�!��le�"RE�� ��u�F�
��LY����(Hti�?���2�h�%x�b��رX���Ws��R՟��v��6���;(˷�;^/à4�e`G$%�8�|��H=�r�E��?�����kL�C�.��۹jm��Mb#�<�U��jI��@�}`K�3��WJ��Y�ZEy�''� �P6��^��U�&!7H���������
9ۛ��]+�l�*}2PyF�Qm��jq�Il>�^6�O���a��
5�C�C!�j�ҔV$��OI�!ו�*2Ǣ���"U+ER'���cYz��l�j�����2�@���|����[��r����PA�"���2�4�A�C��Nm*1r����2A�J^��
�\+w��@m�"#�CܻB�mĜ	E �aV�X�8Ω �%��P�.��v�����:����#}�)q]jE��/�ZB�2h��?���'�������eEKG�������c<��Gc�K�/Q��&�c�l�OJ4������7#�*G���^��aǄ��݊9@��Czp^i-��\joWY�G������y@Bpn0Y?���-���bn�o~�G�
�W���-W��9�g�՗��rpp�EFg�T�����>8W����\i�lUJo�e��7�/!�@mD[�|!�܍�Y��<���N��7��g�=v��
cG �KJ�?nߑ?�P����}�aa� Ȩnĳ8W�-���]� ���6���Gų��V��h����'ϯ��?�/^HӚִ�5�w�5HӚִ�5�7��6m�u@��U���F���-�8C8x��r���:mq�4�����ۻ��8==e:	|fwwG���\������RVnщ��"��[<�R��B`�-X�%na����������y�'W��r~q%�W׬�,�����na�%<ls���r��>��͔L:�[жܱqH۫�Ͼ�/�=���J�Áܻ�$����d�}b6�� ��>99q��I�	^�ܢ^���� �^gn�[`nme�t�&>��,~�n��f�4�M�u_%��T��P��(1�=ڴ�awP�N
*�%mE)-�6:��2;��۰�1o���\,�zT��T� �=R���L�!C�Q��} @��'�����VN�"W�}Zo�ʥ.��/Zśs,�Lo�ڝ��|�l ѭv�Κ@�;���h���s���6�yP�jX[�O���b���ڧx2� 9�� �5h�"��g�)�Z�(�wr�1��m���5?��0Gh�		��kw��n_��v���JU��Y�y(fM���s���0nb�r�� ���)-���6l�J#@,K���FAX���f��{P�Nن�@D(��ƨ�.�����/�U��c,���~xX���Z	u�^S�܀U(�JEF�V}�5�$m$ ��@��4,
�6�^O"]g@�jU�
 �a���"�'�)��5l#�G�z���
�2�lt�'Ml�����}�e����>yK1{M�_�:cB���� ���d���?o��_���'�`IL�GI r�|�E����W�+2�y���wh3��OTWڃ��O~�?�|�pc; s��� ��'��*�4w�6hyn���$I����5�[�����x?�4��,����SZ��j ��L�������=�Pc�_�6�叟Y#�X�(#Q��2���U�P̀k+�D�'f�I-?6#�*#��E�~M-�֤&�C
��P����ĪTI¡R�'q�'Q�S��h�{NY��>+v�-�Z�PZ�5�z#�I?�$��$߸(������R��<�Y.!��7���,=�:�A?n\	B��GέD��!���=``p��A��!�n�i�MǖT�o������{���c�B��M{T"��\'��9)��Ԋi;�E�"��t�q �9��!����Yl�jk:��J�����i{8�#U[)Y�V�x&�*jYXv��$2K����<��4�����#���~&��p2puq)�?���KY�&nNv*�I w���ŵ�'���ٙ���?@�`���nHK�TUjP�%�|�~�`¸@@�'8�C2�LX��1�'�T8�p�W�'�D� a�|#ky�t���a���c=87�A�,T�(��	�h�����MW&q�&�ˉ,�_�ί�.62aN����y�)�O����OA$�WTrt�ԡ�,�+����Xz�_M��v�Q?��Q��n�$�=�]�(����j�ͻ�C���U�bU���`L"��[�ln�ꮝjk�[}��{�������?ZIӚִ�5�w�5HӚִ�5���&W�B�����别�V�#[�$-�@�s�`�G�\��X�Ut� ��:E�eEˠ� <�Q����"�f<&��tVT����B��ʶV�#���/3���r���o��"S'��Xd�l�˃�e6���+�)�4y_������H��Nΰz\T�aa�r� ��ř��)rq5R�(|v{K	�3��f^������/_I�M��j���^�&x[����_�>q��ފ��=w� o�=�j��%�F�D-�@!� ꙽�=.�gG�4�ཝ��&'XBoy�'�z�u�PL�(**yЏXC��û� ��b@�����[����*z�hHuH���  ��N�C"�?�2_���x'�`�X�G�^��fz�k��V[������j{[Ɍ~o�*Q��AH"&��͌@ ��v�2�n�ߒ�-Zh�<���X��QD
�dՊ�#�����'B��mŦ� @*D��,=��ux��u��AFC��
�\�)���K���|):*1D�Y Y�� �T;he4*��J h����B	��r����pk��DT���J�� D�
qUrl,�"
�J?�g�,� &Yu��^��"J�&��(�Ҝ��pe��ll7�$S��Z v3��{}�>sB�׳�@jh&G���
jk,�>��F�ۃ�F��M�?΍�2��iI0��n�0/ss7����<N��PC쑗���ԛj|��,�7�i����Q�e���}x���A����X��"�e�F���< ���PO����{���1�_�7dhQ��A4T ��R�$r�o��D�vjRcClC�q�D 8�{	�?&-KE��A�О�Z+���,��ja�Y1)�m��,�� kWAF c
_+B�Y��=�AJ,t"�[ض))Q��Oڂ�u�:�;���e�	�G��@$o�e*=�U�lY�]�_!ټu�ǢZ�$�Z- ���Y��_ڎ��l*UU�A��=^5俷2R{C�Wh>
�7��!j}�網"�I^�Hb�h箋�@m~g�dT�?32Ƈ�{R��S��V#��mA�3��M8�VZ-d~=a���z,g�ތ�xG�F�J����f�=�`����s�Ү<�Ʒ����x�:���TZ�2Mb����}I?�x���� �;|��w����ruq�yL�]ji��$b�*�+\�w�$Q(4d���V�v�i�D�R���V����ŕ|��s�P���9�gO���hű�.���$2,���\�^���94�ܟ7���G&O&��伿�sT�.R�7���E�8�U�"X����l9�^2��<���s>n۬ϖYe
�L�E���Vg�ڒ���i�:Df
n� �W�!����@����5q��dU'��̞j���"�������X�R���W�T�W|l|�������V��6��'5buT� ��?�_���a�{{w$�scǍM�e�)��<�V�޻�d/�^O�ִ�5�iMk��5�iMkگ��:�p�$(?|��}{�����Z�;�jp̥{�½��kd�J��r��|�X|v���J	NÏ������1�3�v� �ݢ�����Q��l�|���;�L����⣑<^.�o�h7�����R�N����J�'�/����tqv��F�0;�.�w�oIok@�/�s�X"bA9v�6��)�u#�p��JX\�n�� A��C���'r�� ��-�Q����o���h� (7KR;�4������qn��\�N���
�HE��Ef ��w�J�Ch嶈f����0�p��+��&oU@CE�E1��6 `�U�V�1.����x< ���Y_	`N�܇����YP�$q��F~ж���Ɛ ;�[H�O�2�ip2���*�2�NH�tz�:ez3��Х� d��DuU@���-5�%�D\7���ª��ZP�Rg{����E��E�5�Xڝ��f<���;�M_��<��c]\)�l��\�����rE ��Җ��*c �3�Fմ�^�nT�s�P_�m�(!PW�યW�Ѐ��-P��>��T�b� ���p�Y3p���7[x:�>;��c�}VY��A�J����	�ʲ'P%�>��FsJ��Z�"���њ����F�Ti=��)	��V�c���t���Ϣ��oG�m�`W�-�@r�� iR)�o"��}Y޹�My�R�HI�X��dm�T�UY禍�>�s�o���� �\%Z9���7��+�4{$�}��kP�r��<�����T�|5p�����OL�P�d�AmQ�gLd� T�����f0-�˷��cJf������F6S�������p?���$!U?����Y��`6��W�N�z-x,��U�J��q�����=�Q������T6	%��ڎ������E�.a�2�ᨺ��<�s'�����P�	�r���Vu��C�4UH���F���{�G�����T^z��[���nz��T��竚��>p�_ϟ��X~��%�L>����R����}G�����ܾs ]�?~s$���J3>��U��v������\NIR�8o��u/��%o�yS���)P7ƴ�q�+�N�^�;���������={�w,�/�ݘ��Ҟ�9�P21^��'��,XI��f��-��Q�l2�����>���3*dQ�B�<df,V�7��/(��s���?,d:_�JB7���E^��v�/��-�+��
��=_: }��w5v���|�s��,2M0?����q��}ߛ��SՔ*s�q-E!�Q;�U �p�gy�~R2`6��/���ky���������X�2�����OW��|���J�eľ���
����>�y��'"��{�W�����|���v�c�����g(X1G��.��8����������TA���M�iMkZӚ�;��iMkZӚ�koGn1Z�d�%�����ߒ��e�ߛ�S����B�.��X.$	k �?��T�K_`�����%B�ѭ��;r��Cٻu����_��J��@�Pv�z2�od�w:R�E��AJOd���9C�a�pqqN�����\\�e��!�����6Q�v_Qpq�E_��������@��T�^^��ə�(��c_p<��^��j$דkI���i�Gb�6Fފ�Uwn�>^\�x|-�r�
q\#�$��ҵm�B�:,�9UP8ti�Ŀ�T����[ȃ<:;=�E��J�W�< 遺 EEK������"�l����	H�p���Z-! ��eĒ 	�z4��̍���	��8��AÞ�Xz��ou�y����.=�A;�Z�A���
Y�N��/��@��m��c����	�Z ��{C~g��g�8���n��7T�`� �(a��Y�0D��h��`���ˣ��+����V��\���x=�! �4�>�M��- |}���ޠ'���Z��k�y'��l.�<c�+[P��VXu	@*�r��pͺ�A��u�G�D����i�~���<������D�
q�r�;~��^[eY�D�:Kf�$�`Y�/T-�*{fq�[��ݖ���6Jz\ZՌ.�u�]�r x'qt�Jr���� �<_����+��\oW)��kT#ABPԬq���c�"�&6��p#G�64B"����-��a'���c 9�i=t�N��Q >����������ëR�>��>��t�>��w�u����<��>&�M`g=�~f�
��E-����3�d^�&6�iA�/���t��nˑ��c��k%�7�~A}�E`�R$�p���d���I������`M��8���Vx9��m��krc��Qۄ�J�>'�M-��ro���Vzh5��Œ�Yu`��5����M��R��5	GO`m��ek�+�?��Fh����y4�3d�~�f�d�Y�m�W�g�;h��PuUm(���(5����x.�u �j'�Y'Q�J+�R�R2h��9��ٿX���7|~B���K�H�=#a{	�`�7��b����~�����W�=x ۻ{T-����"���*���r��s����|�=o�B�@�!����E��G;���~����Wru~A(UUPU��m�>��*��(� ٛ�]碘�s�ؘڝM��|�y�Q����|і����#��;ߕ����99������o�0[�VV����<�+�~�k���,R���_���IY����g>�IUF�)�}���z,͑q'��|�$|k!CI� �I��8-,�\�,@D�:��P��)���L��_ȯ !6��*·�&����(��d��U&^�Tx���mŅWA��~&�� {	�?J>bSqʕ�l>��͍'�޷n��وM1ɑK*@Vn�u���k��q_����ʲ��bi���O��4���/���|�����4�iMkZ�~gZC�4�iMkZ�~�-[��xS�HX��9T���oqq������y���\OX�H˕$��Ց��r��<z�r��\�C��/T:#��`�P�y��cbvq���br#��B��~m?0~��X���{g8�G0�q^,� �H��'�e<�r����X�̖��b"�4j�����A[�G���+'���J�~��b��_�������Lfn�B�P�yx��i�4�5_i�9�È};��AgEa�a���a g�r�%���� %�qR�[���X��{P��M2T�RA"f%U�2���\-� pg>�9��u��X1Pu!��'��Bu��ԋ ��eYn@������Ξ����'G�O���������
+�@���FnB��M�0����~-frzr)?��G�����2P�(A���lN���5X5~i� �ԋ������oYey�@,
@�g��w:
�.I�Ta��C�B�ha �aj��!1T�4xx����:<�G����Mond����;�ﶺ5@����o1pG�O�p����â�O�F~x;�Z�0�
,CC��r��{�0VA�5x� b�Ω.����Y�ЉW�A6@0#2 ��nZ �=��8F���^T��!#Е&�z�4�T06}n|h+��mhyL��V�6Q^e#���x�X���"�J�(n���$w򕯮V2g�2)9���L>T�j���W��9e�&��T���A�p���L� ���K�j���*���2  3�8���T�#`>�=(�ד�X�/$Kl[� �!��6̟�(4i���g̈ԶD>�"��Tb!���"�{���!�U-o+1*�1�'��6m�QF5c�>�$���8L,�=������z�#J6l�
U:Q�#Jڤv<k�He�l	���$}P�Wۦ��?��8TrL�s���bE;M�����^�r�������}����{A���ڦe���vII<U��d-���ȍ "��	T/G�Ĳ@��js�1������Қ�	-h�vt$0��g�pg�OX+Hpo���#j�e�uS����P����tӾ,�f��q��_|�9�b(�
���=�f �W ���ʪ��~px[n߻#����|��؏d8����wN����˗,���I�֫���b^1_��s���v�.<s \#}�o��VOZ ܗ�U��!�)}F�VY$���Ҳǐ�F����L��R��(��9�C��ϼV'e�.n&2w��"�תn���'�n���cy��ﺹܙ�9�'O_�G�-��o�} ���G���ߗ{�<���}�l�˳�_ʗ�.Ͼ��D�MFU�挕�wX�b�b>�r����y�9�9W[Ű�Aḁ*׹�ψ��[fx��X�����@�VT���q�6T���(~��Fh@'���#;;��G(��F#Y��o+��1�6��Q���cNl�_��֜���w�r�{�5N���|&o�Ne�)�i76��>���W�LF�n����r||,ggg�{>�[b���?���_�_��6��z�+MkZӚִߩ� MkZӚִ_k{����������[%܆�]����������؞�˅t�Y��n�!'��?dP"����O��!��{�/��y��{��5+��U.ݖ[$9� 
���K�j�d��"���E� B��,{��=��m/I;��P�n1vqu%��	��P�k?/���	��2���-�w��\П�9��_����-�\�E���<P}�m��
}��3���=��n�7��GGnQ� #0?Y���XeN���=)r���c� @�y0'U
@��ѭ6Ac�\�ɲ픢,"�S�Wb��0O.������{(dOP�
��$"ؘ��ӹ�{�s���b rj��+���V��y6R �=�+y���o�b1|&���%��3K
�� i��ϵ������͖2v�~����|�R.�/��ݷy����n܅q�ci����h_}ѣ�D(X1� >7���8F�' ����#*�rT^�!��K��
���y�~ _'t�Ԗܒ{���*&�-U���M	.i�lb
��*
�e� ��|����`A0������S�/��{O<�0��]Œ ��}�j�!�&��Cg�� ASi(�����$���S݄
S�&�V��*���n��@���l��̲�*;71m�Z���.z���k�oLS���Ӹ�&�9s���B|���� ܀��^�A��}&[�h�T�W��8�k�jg���vGIVT(����mw�}v����˂�#��U$��i��ɬ��[�F����`���� �H�a�|���ˎ��h��jqZ��f}�sPH�,"���l`�����q�	UiJ���)*%Bs ;��4���v/��]�
}��}[� ���ަcw�BJ���ZѤvR��"U�|���$��(����}�!⢖PU�·iٱI��Tٔ���i�u~	��O�����N���'��J�>�	
o����PqY[��\�<��J��q�DvhYAm��}֏oޞM�/��ϓ��rD$����[Q��ܢ{?I��2��##��0���Yna�Q���R�-��I�{��&�kB4��6yf�U���� �Wy0�#��u7��V�Cձ4Ϝ�B�>�ٸ{K��6"*� b�,AW	("�-2���ы��:(��T���w����[���|���q����F����+77��O~$�?��ʅA�͗���?��n
D�J<�fn>�r��)��:���3�����X>>9rs����/XH�|i�y��c��=�	��ēԅ������"��gD.��K��g����cO�9/X��l���ø^����&�P�zk�|��d>	@}�3Er�������G�S~�[ߒ[��P(��c.x��������)�w�<�]�;��o���WkK��j�N�OA)�1���1�l��E�7T�Жj^�'x�g�@��gB�h&��ΉɎ1��űv�1s^��#�۫{�[x��%
&p^�Np��e��hF��_��U��$"#BV��%����v���ɋ9��ABCe��#7ߢZ�]ϙ�P�zn�������Z0d��{�E��j}��������-wGٖ�5�iMk��Tk��5�iMk�oD����A� j���  �P���~y�-~���=���U��n�r��6Ɂ���$B�s�lo�b��5n{���n����9z%�+Vb����-�Q��ΣG�]t�"!�[X^]�K��u��g�(�ݟ�����'����[-,�8FS����� F��9V��[��c��A�x[!4���tR�|"Y���q�֕�[�V�"\���m�{�6	���T�ޜ2�U��m���i���v���ޅ�&��XX(�֠*�L�A �h8x&���g���f����T[�^'`�:�M��e�$P����j��<����#��+`	6)��} ʕ���-�W�Z-������G���/�IT�� W�B8�~7ΧV�̏�M3#Ӊ{���`�OBd
@ ����/Ǭe�i�vS�	|�7�6�4��%���u�1U)"�A�bl����h�W�P3Q�����Bza��Dm���^iy+m��pKvvvh�¼��~%`��v���)%��-u31��n�4; ��	����X�8��׭������bm�TW[���]� Ȁ��J��|��Q.�nʃ�T=X��x�Rr@Vue�� �8��Em���\dP5���m�v���* �]�p�T(aT�yW1U�d����*۽���k�JxB<��5`}_b|Veed\���"T�jZZm�E��s v���*y�����j��8Q���
��#U��s���#�yYf�`�bz?T�$ �ǇZ��\A�,�����c��<�X���c��e��8�"O���	�o�WO~@��H� tU��e E�Q�VL���[[i��M;**��B�7UP�w��� B���+���00���/��l��o�L]���C򓬉��o��Q�5(PS�k̫�0V�͍g���$��}#ش��1��^}]z˰��'�����ͪ&K�c1��ʥ�P������4�J/<�<q��FF�����cX|__`���İZb妞[�c�R�r=."0P����Hd����G6.H��J
(�68)Ӗ۷��~��O��?���>����C:���B��^��Ǐ�/��/�o��=���z��Ҏ��NAo��+X�Z&�@w���/�����\~��K���o�륛W��J8��Y�>�SU��t�7��R>�0�i1s>��7����ӧ���|#	l�M��
��� � ����;t�%ؖb,��2t�y�_;�Բ�mc��.Ș'��Ź"Y\�~�->B���;�>���鴘�R�x�Z�,�;��l&�Ղ��$�U��^^��%k�1Z]�o����P(��ڈ�����B��V�}�P{r��*Q�X��wڎ9W�q�02�l~����^�rs��%wN���:S$��B���S�h�	�q������\��ɬ*ݜ��ȉ
PD���K̯K�奝�b�=.���� ����˧�/�UdŰ3��Ay�]�o��?��>����D�ִ�5�i��!@�ִ�5�i�1-r�BNH �Vٖ+������a%Ij��Duv�� ��-������k�A�y%9,�`�����@�v�����x�Bn�7�&7S9?=���[��s_�f`���r�>,�ۿ�?~,/^Q��i��O�E5d�����fm�ב�-��ګ�74� %R��;������HC�W�D �F���{�{�z����*���F~��`����bq�X��YG;��v'��D�ԬV/X����o�in�;����=%�m#�(~Ob��"#S�y(' ���q:���h ��P��Z/�rq��Zn�|���������� ��V�jE�U��d�H�Y9�^�Q�Y-�Z��	��8Z����ᢹk��^ep	����P� �*bh����7���j�����
A��e?��j��*s����i��4����I��l)7��rq�ZNߞ�";��GP!gh��.����"�� ���@�������w��`�]����\^M��Z��S�R�j����0Vۣ���
~~��i�\�B�G�g�o����7H 4�X3/�=(2Ux������G�/��Ã3�mhXy s �kc� \I�v�ڥ�L�%��YV�W��`����3T\��n	nu��V���A�������ZA�5b�����6��2���zD�~D���+ :{"�U� 5q��Z�o��TY�K��b`�K�V��������	P� LOt�y ����@WT��x�$�Y
'5��Y*|���Oh��Z��3^9��=WKw����,���4���@t���gO�`t���\+�9'�pk�T����]��J�j�������,�:��n���$��������~K˕\�`(H^&]U�d�kO��2ظ&�����8a��;R[���1�����~n�c���<^\���R[N��h��n�$�D
�ڈH�5ꯣ(��W�F�"����������l�)ux]��)��W:OЗ��*��*��YY�I3�2xuT�L��l�Sm)ɾI�>�M�E�t���9������5f�UE��E���z��y7Y��/o)�Y.O����ccz[1*x����,��1�� �p<E�J>$@�����_�ñ��-����w������/�K��_�B���$qߟ���
!`;usu!������_�$O��5�3P@����Z�RU��� �b��4��MO��X<{�T>��sf��O��vD���T��\i��;A��{�z�X�G��JL&#���h�>��3��.Q���]қ�~�g�%[�vܞ�;ڡ;���=ڣB��q���x�#�x/�Z���e�����O��7���ѱ����o����ƽkܐ����ߗ4��ùL��9�7���h^mI���\��П�n����U�BF��b���-3&�g�Cw��9�TB��x�7�?�{�X��g��kAeU2�p�']7�xs��=�!�MmG�!��vs��Kܻ�H�n��M˺s{Jf�������UV�s������,����u)7o`MY^�g��e����@I�y�w�ei�dE5ʮg������n���Se��>���7-	Ҷ���m�?h-Ҷ���mm��h1�!D���=:��[�aю|�u��j_	����|%׳)�؉`1����j&�U�cI�n
���L�	�	�^,RnQ�����,?�P~�|�o܂zI)��٩�M�Z_�2���K�b�i��Zf77�P��5 8 �ѧ�5+~��"�t8�s1��6�����d���`%q٧�A����U�X�#À^ҁ�yoh��H��p�L��߾z-��T>��#��?���{���_��wg�X���ꬴ"��M���
"���tY}_��~^d��	�$�i���R�^�MH�c�o�r�
�4�3g@
Z�U�^b@V@��U �< PY��Zm�R`I�d%�V�vWX������bt�}��KΟ��\����'���,$ (�~���%��� Vc���>��Vm�� h[.
��j�q,�K;��/����q}�Jɳ�� "����V4��I&���=l��
!���O���8S#9:��s� *ګ���l��4@5mi�:�O��XFFz�U�Vm��r�#�_��D���!�e(l4U[l���a��U`�`S�mu��QV���5�Sg�(!� sQn�6Teu��	�hH4��v��j��[YQ]U���FT)����^�5��d�X�^Z��Nc��e��J������8nT���N�����a�-�<	�L�0�v#);	��c��g?2���=��3�:�[�,>��l(.��ym�W:Ueo�"�6�ݹB��s�AG[R�|Y�U��U��UH��{ų�FWɂ�v�z���<,#�W-{2�$<���-9�1��3VDn�_oa�A���;Am3��+mZ�nUh�W�عW]�[��o����c䃾�P���
�A�9̓+���A���|�wm��P]a�}�Tvx��1���I7�p|�=��&��N�&?j2�R+>o��0伪�&���IS�Jz�z"��ҷs�JH%:A6VF���d�?^QD�/#+
˧����<��5ɴ�\��E�W�a?���TK��fx�zu�4yA�^/�R�q�� ������w�*���֘y�������G�ӟ��=cw���

`�	��իW���>����RfP�ƪ$XZ���Hn|W*�A0��Wxo��>-��0�;o�Eů��(Ӏr<[e�?��r>��:�l�S����c~�?������N�������[9�����̽ueR�1A�_=�{A��"�"W�Q����nB�����]w��2��-�J�0_�b��\^��w����jӃ�]9<�u�\���ў;�����Y�t���j���z%�s*5d>���
����(��1ԟ��>�*�g<�A�I���Z�6S��S��V��wH�t%=���~��;/�#8N�����c ��e�^���~9޻r�lp�w���O�6pϐ��>#�Ҏ㟨�l�0�����˞�x.�
r�#�o���5�ݣ/�����9C�����X�#��O�7���r�:�k�0��e��?�_��go�����mmk���H��ֶ���/�4C��А��x��;���ZVn�cT��tXn�rz����ZfjC�3Ѡ�b#qp�oT��M��ѣ�n��/Y�p+���G}�r��9*Ȱx}����y)�[t^\^��-���D�%� ��N(Xl�Q_x����&� ��f�S���Ś] ��"����״2@xe�t� 	J���Gy���P���_�֒f���P��<�W{^o�p�@��}Z4���J.����ؽn���������r���!� j��^�i�U��ƑV�Ӛ'�l������B07Z]�E/��J=�#�`}5sh@���D+��]�Se��&�r�����*�<^�/V䁟9� ��`�c�.��?��ĭ������p��a�����0�qj�BA��*;�N�V�[dFC���������s��y�*���1�a��B���\�{�U�j��}����w��������[�oY	��L�t����9+��8 ;y>!��'g��*NF�
�W�U&���0bBDAɍ�o0K�jе���@�{K`���o�ԩ�
�p�H��/���D�~.�Uu�"���f�rɇ~W��j[9����U$Xv�'s4G$������"յq#74Dp��~��n3 0YmC��[(H@u`<�2G�P&��f�x�4��"�-^�B���i-�!%Ѹv�
�Y��v��/�@n\�$�%�y�3��� �˓A`$D�P�eM�b��l�
 �2"����V)�p_ZZ�Zm�oU�ɂ�,�r��b!��=%t��� 
���K 14�(�6�n����I�/���Ӓ&�Hz`=#�p6��}h}&R�n#m�6�C^�
���Y�%{}�����OoʢP��:��]�ޯYR%v�eU7@�Ƶ�̂<�� ��v=5��l7n�Ce�3�`��5��25�$��.sU �9�m������ ���ùoD�Wr�ލ������84Ǆ�(=7����
}@�#��ĈE��D��$7-��9T㔼���I�~(��Q�%��~��fQP)�uǘD�=y�@~�����hL�J��~�; p����	�{A���b�}����o��J^<}&��g�y��Z튘�%�B��	�MS5�@�8�-�4����w�JJ�?x�Hޞ��
j�M);�1�E��LK䲭��'O��?�������g_~�{����$�������; �K��P�'�΂ͦg��j��AA���_����i8tמ��x�rǾ��/�޽�/� �J��c������e2³n#�_�����{�/��;����y/y���1���T載"5Oyͱ�dЗ�
�i%���/�V��,ɨz�c�:Kyp�9��܂�T?r��9����@I���oX��z��;�y��ȗ�8=F�m�;6��c��*���l��^�*, r�|��Ov�y�ޙ5��=�^��-��f��W�O tz�ݭ�缐T��.������G1����BNݻ�r�QP,V�G�=�ˠʪ�Z����~�ꥴ�mmk[�~��%@�ֶ���m��E��-ª�b���ř<�-�o߼�U���r���F�>�����vP����Rî[������t���|)�o����%�f7Wna9���CO2�h���h(?�я	��Wky��BE��}Ն @AP!N�����=	{���[�Aq��;6�o����t�@��`oأZ��
@�R �b�|���EJ묎�'}�#�t2b�uU�a�xs9�w(�=~(��LXٟ"�7�Hi��(�1w�+7�M�;���Vm
r���0OV�����0�ڬ	�n6]���k� 5�ͭx� 5��� TWn�{�J�z;T�h@}a�y���u[��kkNHY���*�>~�X����K�q��vyyI����62��#�tbX/��dH��~�F��ځ�����(�4v��%]7�+y�⥼|�Vmmj�1a%?T&��͙i@;�҈���R��ua�RLP���Zm=�S������?p��R������D�dR[�Ѫ�k���+#���{ޟ�y������·+��a9�t�Y- �-��+��nL𪨶�h���Y��dH_�O�e���T>\u����X1巋�g�&fICB#������@��A�ՖF�*��?A� H�B�7_	_6,��X0��RK��P�26��nsy��Q��S���9V
�{K������ TIfi�C�#���v-v�|fP�
!�
P��֨+#ЗV{�� 4CX��X�yBE��74%KA�<4p�RƪV�@���ZIȪ�BI|��*�ͦR ���#8� �|O(�\�*������R4���{�z�k��6��2���ϯ�B'��,�����2�2b| :s���F/6{����ϓ��=�w��!C���m��� m��ɍX��O|�۬��F�/��x�QC�;�T���Yj���+#Dj5��AE���D>w ��'��������(���PAU�L1[Ԝ� i���RDj"�זe�p>����]U[�0�vR��i��s��]�#�;�c�h�I���'�LM����������/!{���;U�Q,@����2������L�}�T��ǯ���?���~�l��(Ѓk߸w�#9��4�x_�:9P;��k�(J��P-H���gI�o�s��9�w$���*��E/'�p]>?�rtr߽����2��r/�[͍\��GE�������I���ݩ\\������c`?�]��A�L�QՁ��~5P)w�i6��ʽ�#y������ ����IX�����1,w
����v3�ۼ,-D�W���C���^��JJ�DƵ@%[U�[���
=fdlV6& .����š߯��-�w���U��^�Ѣl]ԡ�w�η
7W�ݾ�L&��l�*VBU��P���'B���`�֩�O@yU!��@-�e*3���w8���%ǉ��
�����rYvvv8?kR�Bf�N�?n\�������⥛<��mmk[����n-Ҷ���mm��kWg���W_����t�.oX�`Q4w�uTV�R��L��/�b�-$�@�n�z��썤��^�rZ-�r>�����-�&�>�QYή%�:)���O��$u�O?��|���\�3�չi!��{���C"h}��=��-�f��]ȳ�H������������uǀ dg��c)�B./od�\�<�\���m	2������rYԁ�X8"�2g>G���h$�����	�.VkV���^($)c�"��������.+Z��{}S~d5��_���,Y�7(&X�ӷ{M1MTZ�� �e0�s1>�E����{n��ye�W�T�'e� ��|�X�4 6�t AS��``��/YE
� �Jg�\��Jф ��Q��UX��	LEO+��9�I2%*��VQ��fw��+H��B���d�\r,�p7�V9�UF�$�!~ ��� 90"���=h�������� ,ŰD�k�Q���Z�������徭�M��$�u��sWif@�C~΍  ��IDAT1h80�ᓐ�����ͥ�� ے��AzV���k���[�V��-��y��kEC���� e�r[ކ����-����k�.���؂պo�����l���I��J���.�S��Z�R���T5Y�������RVO��
��iV�{���y�T��Ez�T0�}���+t�+�&�*�ʪ(M!�-B�?~�B��1��&F������>�BU�H��lk��(��ΜP�+��=�Y�J�m����� l=g�-�}!M�����o�4r7�SbVq ��:�(��*hy#P��~ �.��.�W�q5!�ǭdV��o�>F���������9��<O��U����J~��B���5A���Gv��{�������9�`_��=�L)��.j��*�ʭj�YP��u����$+cZ8��6K��! a��?G�G�D	d��A�5B�A�
0��󤕿�t���CV��Tl$~-�I(�l�y���4+6%I��9'e���]���g�ġfLy�.��CC�쀠&DK,ς�Y�E����m�@,��;�A(� $ 1���t���AWn�.�ջS���Ky��o�ݻ�����&�>tN5Э�W���p�����|NU 
�\�iA�Y[����g�r3����C����ss��������+�z΅�֟q��[��^A�9$g��2�,���y���������}�ƽSA偢�ã��&H"(*�KK���Ck�H�f`�yՍ���
Uy0���9	��PB��q�e�,3�7��Dlb*���Ӣh�����?��#�v#fv�*l\K����0�=]?t�
EA���6\��_�~���(�UJU�4D>[��,U�{=J8Ҵ���>p-�;u��v�R8�`u�+.Ƌ�%^�JU��Z��ݡ�3�v��ڣ�7ĉ����T�(7u��K�b-g��y��,ݻ�ms��b�\�Xza��5A�̎���;�?e��ֶ���m?�� mk[��ֶ������5�ޢT�����-J2v�^/�����>9{)��f��Et�-�F�-�"0�L���������o�~-�=�P>��y���[����g�e:�� ��4 �(��ݑ��O��}����O>q�����?+Tg�[X�H�X�� ?(5>��99��㺹��l�\��y|XXơ\����7P��Tr`ш� x.��93K@�<�\��]\rabED	�L*M�� ��b �p���B���	$�4���ť�PQ�>[H�U�[p �0�ؽ�� ��?m�f^X�z��qiPg��کD���	}����i�
� TeǛ�<z|�߃����/H 5���2A�w�s�*-B�[� dCx�;.���"���-/���c8�c�-(M@�L�c��ۓ�pD!4`�� �f p���ɾN���;��Z� Ƽss'4@ ?��6�����P`��R5����G������J�rK0��)��;�zyr��b���Z�!��e�`���Ǟ�m��N� ny���&~!|I@ׂ�	��pK,'�,� �(q��騚 `�����pA����Z���B˭�72�rv�ĸ��=�5O�����種��͓	h P�d[�����7���bK^�jO�
���}�vg��E[���$�t��U�{`�<�I�M	T�$n|�Bg:��L��"Gվ��W���9����mL4NB���Z�P!��~�.��cy������%F�A�Ȟ;Y%b�n�y'�"��%�^�	��lVٿi��ki�+%�$�ji?�<��8�*3Hv�e}]q�)?�ꙥ�_��7�yPgq�ܰ��h�m�5� 8�� OS`)p�93T@ %m9
˛�y~~�6��|�$�o\�wr+xN�������ʂ�V`���T�Y��=!j�U�ZHa�1�pg���J���d\�yUJXS��g���sA�>�,���i�8F���y������r��" T���@E��~�y�����C[#���y�0��b���吏b��e���kPD�vK��VI��Z� C����:�Q�1�*��偩6�靮�2�8��������M^�zC��=w�̧7|�@a*v�L��
:��# o�� ���x�H�E��}Qx�Um�P��y��jT�w�n�,]��VkԳ����%�����a� ydD �S���l����T��>��1�bP�N ���|)�=q�n��>�Qd�Zϩt�
�c��,Wr9p��Z96 �1�UwY��X�{���!�ˠ� ~�"�0���ʬĴ�p�^�ג�"
�O���o�4���>����}�7�g~F�T�|��i��eW�] <��j�I^<��ȐI�3���Z�ǹ����_4qt}I����e�c�������}��|�}�r����*�C�c�BZe������»0
o`e
"�F��C����[��'����- ���z�&n�C��̢0�b�Z�ɳ ����헓���mmk���H��ֶ���/ߨL(��j�����s.v=|�����<�ܢ-�~�K{���=�����J��9�,���w{����������,�3�q��{��	x>{���9}'�����}�<���ᛯ���k�m=<��E'Ș�x$'Ǉ����z-<������O>��b%��g���w���[��9�;��c�E'<��݁�ˏ����{���2uǳr��[����G�&n��K�pw�V�cV�#��e���@�PvC�2���>uJ�EX�g_~�N�ˋ��T��>�
�8���U��h_r�0�*)&��Gg�I�Րg���>�"�ɘ^�E��AX�#�$,2Z,��؎��eg��]�ٜ�"�n�Ͱ�fv�E7���TT�,  �(�j@���xǍ�#׷����k	Qd2���Bםk�̆Rvw�<6TbD�� w��?췦3�z��x��5�tz�����bn9QW���LF;r|p(����gY�q<�ݗ��OHx�*����}�}�ْ���w�jg1r���	�@��G�LI��� �P勊R|�t�)��͞H��1G4@��ۑ;>�5�p�"�Y���l)GG���$6�3�"��P[.�~�v
2}�^��X��w�$EPq��i��h�!�
��_|˩0�o��H�l��}�����-'�  ��m���V�� �V��@��LT��0>B�ӣz��,?�eSU�p恻�`�v;8��9��~��ti0��C�Q5`����/T��	������/� :���TE6�Az�Vm� /m�
�B�6���W�X&}7N4A^�*-�i�¬ wӀ\���>C�/-h�(U�>�^���2�' �����8��UF��-��Whe}dY%a�.�Pj{,�fན�^�6e��>0YI^uЁ����Zwy��������j��Y]=��6�H��x�$>M�~k������1ǽ�!���C�Vn�YB�Z��`�u�>�l�B2��SY��Y��/�h½a�Ȥ"Q�M���,H�0��첐ID����$P0���	BO<�%s�l.`�.��
vrP ��L�{�Kp��$�pP��Q`"�Em�(����+T�A�ą� t4H<�g�Z��38/��NL�a~>R;!��(֐h4��`�̝��*�A���蓮�4�,�X�@2U���(�s�Q=Qf�}���{�U�c'�gh�gr���yn�� �����={_���r� i���n��ʽ�|���駟28zg"�=��]�W����\\���&������")st-�p7��O����9+�����	�>O�aܥ��`4���R�g�^�g��D�/�:�Kt��u�wwn��L�qߍM��6\���R�{F�����o��5\�,����J�[iA��..���E����{�Χz�r^��s�/z�@z�r'�ۃ�{�#��o./��䉞�����1�ҕ̆�9�� o{�oB�0�{�L�{݅{�\�|G8�Z�*8�����Q�!��\U�bN��}R�!ռhc��wl��A��2�\�}�&����ucٳ�^��=�cw�q�u����5��w���*-X���p-�P$�i�H�^?�>�
�J+�K�3��
VY,OHT����t�������S��}��P���3'�Z�� F�/��JK�w�u��J�"�I���XU@V=�������ֶ���m?�� mk[��ֶ���jZ��Y,�2���-X�����n8<�e�B�}1��4��B)D�bU�Qȡ��s'"�D[(�??=c�9���>���ëg��aQeyrr"G�T[��o��GǇ<ƫ�y���|�e�*T�=���LgS� D��+�݂�`���ݢ2Q���}�b�d59�7X�*n�M����aG=z��y���-��b(�lX�^OM��I� \@�^�ӌ��B!�� ��:Y�&�j�( h�3 )V�Z }/k ��k�#(�c(� t�-���,i�R��D�`FTM'��  �P�,b�o�5�b:�s�_o��=>>������✤�):��%�����1o8X�E:�HQ1pҝ_�S+"q�<�����0��@�22@K1؟�:p�����������zL�ƌ�ڙzr<B�j������߰��Saz����̀;��; 0�AE5@�(�H�����F嬒$
X��AՖ5��K����v�R�W��g�W�F�!o�+�I����&ܵ��ٖV˸�Fu7?�)�5�Ѭ�������`l3�Y��x�2$*IJu.Gl =�/fǕ��1_	�~�\
UQ��^iJa��EfJ�0�3|�u$�<
/W��	{60��+��g��>�Q�ո�Jʳ�כfwD$L� ¡J7�� m���1�ʁ�T�Q�͕?��=���x`��0!o%䭩�p�T	L��YED�� \�܇��HĂ���j�9*�x��.��S�y��
#U�T�y7�IDQ�c�T�6lܟCm��%��kU�z��aR�;��m�F6��6*w3@��b�^+�LE�dGL��D�Ve��MUŹ���Ɯ�Yiݕ�vs�|ܗ�K��/A����ךo��ڙ���m������>���Zu�AUezr�$Y;Q�����[���#���<��g��Y�62u���(Ǒd�r*��m���ـ��+!�yW�6�j"�?|^Je3)T2Z�<
 fP�z]2�:`��̬r��1q�9��o���j���c:�ˋ/�����Ϝ �\���+�8;���sϮ�ข�ڬ7��%-@��f��:��ZE%�I��/��q� �l>H��'����hx�W�Φ}�c�g���J��{��;ja��@�~7�G撁�)7ґn��&��vIz7�U��k8�zT���|�� �GXd��a��QZ(x�*��+��}��y�{"�_���u����*� �u�T�Г�R��H@P�!�q���3~�Aˊ�T�*��
���������$��+9,$y�|�s����hׅ��u���ғբ
,��ΰG��?G�A7'E�nH�'`�c�W���)�t>��lb7���4�矪�ݵ��<d�K���Qm������ק暴Ƶ��ݽ]��'	�")߉��̞������g�hJ��ֶ����Z�mmk[������z�^ a�� ���q�Q�>���Zd=�A�|I+��>�"WWr|r�<Ky������?�)��5�J�ͮO����2�_p��Lz��3�X��~��ee��չ�V������w�1����Z�L�ܸE/�����D�ݷn��l;����b�(��,w�t� C2�#�P	�bo�`_vw
b>�=!�_��%XVQ��Ƃ{8LX,.�={B��pK�h�~B?N&#�+Q�mἕ��\� +�I1|����+V�#�wħiT{	���p���>׬P�mOX�����D�g 2��R��y�|%UH"��,���?�w�_ɋ�˻ӷn,C���w�������K��ֲY�2�WlV���� @��'�;u.	,7�]��-'O����ɓ'rr��Lv��f>�o��������O*< �vb��#d���Ƈ_c����B�E��YNAI���(yL94�N�ᵲr���:D1@����.�O��{]U�b��Añ̗�`d`W a�����j���g  �@�S���p_�VT���[�2.*i��Bm<oOp�����L�mE�����TU����P��gPqYl�k�*�:�ZE����@{�U��r܇"���Sy]	�<���\j���o%

��n��*�.+�cUF�s��%Ub��6sBm�Ă�3�S�{�<ܸ��Q߂rӺ�_��<Q5��:jb��d�6�}���ژY6�l�2�6�)
R�����v�?JJ��<�]ԤT������d]��a�(!W���R�nb���[�J)�9^��QVE}#GH�J������|�-��c�P�{�d������V�G:�unf&X���bdGQ���M�|O�0��?�U�q��;o�Mdj�V��l�?��q�4H�:g��������7/0ClvTaM����T��*������\�`r�a`��*7|NILL�S�	��E�^��lDu�P�et��y�w��F'e2m�#�{:�}�?7)l�^��$�9'>ӄ�ja�H�!@���������������A���Ź����w���\X����������i/5��s��3�sH���  �D�N���Jr���Ϻ�w��g�'��@����1��*Udk�!�m�:˲X�f(�x�NTd��B+L�^�.������\	�m�EV( ��=�P�s��2j%�r%B(�B~��d$Xh�G�I��u�k������jK:�,P�W����a?D�z��L)a�ҪL=�{8����פ{�D(}B�����κ�U'e?�����a���!йSZKmS'j=%k1%^+�J��P�QX[��<T2�`��#w�fFE�$l<}���k ;޽�����.C�hR*��^HU��hG����ue�K{Ջ�)	;�獆;,�	{Kq���a�B(���z>��D�G��u�mmk[���o-Ҷ���mm��i��Z&�+0!�ǢR���Z�����ɽ{��'cy��+%�x�.v��+�[F=.jv��}���P������ �j��zX4]_-������OX!�l,V5Ȼ���^;�Cn"r<.�(���^$A7��n���uh� ��3�ٙ��V���|�\���"��`eT��ݱ�$�vd8����P&�]�r�B��3� ��#�`#��\*8�S;�N���1K{�.��	�̖3Zi,'8j�8GH�>�n���P�[X�(�i3*��m�2fR����m�y�#O;�ɳY�x�l��8V,�1�����hk����?ړ��wjy�6t�s(�n|ї� +��-٫7����\�_�:�H�|RE
�V[ fn�<�Ϙ���98��'�����{{��@��o����Ç�D[a�\`Y�� H��PQ�*�XGe���ݰ��k�}�L+&�5�¬���A��K�%B��JF���^]��1_n�r�|C{6�~>G�&%
��j��7_��ql��M�#�`xV�z�È�p�GY5��Z\Zn����藺"]�m�8�ɠ&;��j������lP�p�ݟ��2Q�������L�Uuk58�eW(k�M�6�v�F�GM�׃�$U����E�����$����ؓ���ZtiI�4��#R��>4�����j���J�(�o9&��~�����z,*�fJӒ	��8��h���fiĩ)KhMCp����/�@Tv���sn*l����W�k:���q������EI�-� �KWr�⬙��`�F@pi�*XD���f�����]�c�D���)��5穑d�Cե��i^ ZiM��X��!�Lb�+ƕU�ea��tnY'�/�u��|�[ x��m�UU�D����q�-W}8@;K�|��%��ی!��3�l:�VVnS[��_o��CgfK��=��j>�Z|���x摨��m%G*�9�\T��k�" C�y8���`a���+�b�^�R�v3r[��S��P�F41�R޹g���s�L�!�����r.�ٍ=�E����
�s,5C��d�Jܹ��h���%T���7e�,<�6�u�U�7#ͫ���T��c�tĽ#�8�������sJ�
�"SkJ�vı��x"�s��D����u��	�_ ��U�՝5T��Y-yQ�%헌�����FIx<:�K2�;�W�l
i��'�I52��"^c��YU�NDa���b��fiNKF<�(Y���PR�rvp�u�ߓ����<�x,x%$D�㊾�q���T�I��2d���X�I�4���P���2����	rd�;,����"�g}��*���s�r�K�� M���u7����x�VVPZ���3_k�u�����e�TVm3R�V�-�%���H���*ZUl���;xw
T��8��mmk[�~�%@�ֶ���mU���-�؇�7 ͽ���w,F�_� HI/�5¥aOe�#��Ç���wr}}�����=�xw�V�"�H72���³
9>:���{Lu����;9}�N�ܣ�?R ���:�A�d$'��`E�O�s��)@��d���3�+I/�4��舠�C1����X:�xs��j!���=�/<y,;n�����>IB�P� �7��I�"�륬�KV�1w}��}�!�X�L�1doo_޾}+��Hq�ڨӣb �r�4��r8�@�r�O� dĆ���Q���M�����4k��L¿�\�*��A/���;X�������3G��S⃮��*@�eaM��� ����[��A|��O�l�3KQ[&5+�}A'��N��6&
���Ɯ��_���9vs}���T��X���J^�� w`喹��>�B%��U���X�Yup/�1�&|���b�F�%� �`��=�j{��5�/� Rt�����N��[Z�i�C� �<�~��y�N2ؖK�Rn���fyU�C�m%8=�+�a�4A��y���ʇ�7 X���ڤ4�GВ����]O�� ��y,�3�FGCܩ&q��9�����U�sT"��BF��(��� �?XrjaU��sO��w�-��vX��R��y�.`��U�UM4�VLeY+f l�Y
Zm��>g��U8�J{�Y�k��*�4��V��C囤^��l%�V,6��*1�;��i���$�����`1��bE7Fk)��qKA�Rg~D�yh +�m�4`�=>��� 0jp�qy���SY5J"��ǏU�Ed92~�p��MP�ɤ�"R��x+�e�N��,v�f7�8V��/��l�,��q�&�k��y�����$�<y巯yI1'�vd�_��{"��
��I���&��[�!�1�q,h\���'�{;v	��٘eU}N�@��'��
Zm%<v&�j�0��Oi���'6��H��e����U� ��jK��yՙ���� �U���~��ܗ��;H�)d�����@��|���T�G\��:ޛ��R�x�u�9�;����؏g	����`<��{n#?j�l1UJ��g*�m 9�aގ�;�{�eZ[.gsZ��EF��7T���m��{{{|�b�?�#���ڪ���F�Qf�����>Xna�^`{�c�{���n\a��7��e2e8ޕ�T��^�<�!U)��Qaj
R �E���T���ى����	-	0��nJiU��A�����u��]'�H����z.�Dv�:*�b��D����҃��*��z(����1X�E#�L���x��{L�������#�T)l�V$A�^�:���h��9�خ���u�FV��Zh3��}�v������z���e1��{8�b���s%�z�v���M���D�vF��}$��ե�;�ǿ���?�g�|�D>�ꥴ�mmk[�~��%@�ֶ���mU�}u ��f%��d�����d(!A|���B��@%���`��Q-v����\]�l��	�G�}vv&��W��w��{Od��O�{y� 	�{�'�j�2,./V�}�����O����`�#/^���??��w�r���?E|�HJ�	U=��� {$�#�ф�u��-n�v'r��D������>Ar/�w��~������V  �g���b���]�lf5���A2�_Q!~xp���!�t���ПQ���	���>H����W�9Q��-��ޘU�]+V�2?$[ӻ�Ei�hZ%��n�C]�\d�������O<�F����@N�1Wc�\���FF�U�ˍ��[,/d�XЖs#- @@j%�� ?v�#.��GI�w:*K5�v�3 �� TvR�Z�x��������~���h8}��a�_�Ǒ� �t.{3�;T�@�K���]i ��r
i�����A����Jk�s�ܣ�����;����.<�}�����޺��AR(�Mk�D-/�j;�����3IP��-��
�W@7
�-�\��9� �WA�L�s�j� �3C`?G2� ����F���JI�@�8ì"�T8��aU{�7T�������`���n��f�:��G���U&��WC��
P�1����5�cVu��y�[V	��7��SU%f��2�W̾������ji�G>L���e���q�r�c�\�U5@�%�_S��a�����X0�YG��_A7ͫPR*U��1C�0IێWYp�����p\��+<�����j��a�����Bj��W�IU)�.'W�'ނ�a��&�,��g�t�����'�jĈ�B<_�&���v��f'�T �mu�X�<	s���}�d���c�J��g�4�e$��~qmG�3��C��Ej��t�hZ�mɥ�A!RI�N�Vvk��aI�OIWQ@�j�n��s��b+�3;*�&��h��*f_��W�ٙ��{���4  �]S��+��05���W����E�����P�	���X��rG�)�*�������ʍ�r���hW��5��X�O {;���Ѩς<�V G������?��wTy�x������^���z��K����Uq�Y�(��k6��O0�ݝ*�c�w�b���n���ؕ��QMrh�"z�u\��������w���L	Q����j�(��bT��[^����	���P4DɈ�|�󒷻��������Ɠ�{_p�n_��{wdaM2�9iy�rޖ��P���c���w��,�������:$�b���[�������J|���_�E�o�o�t���,�-I����V���V�����(��$����z9��BU��#H��,�wE���[
>��u���t�`	5I�{2R@Fa����uz�}oH��b��ʽ[�:��=�S�č�L�(ݶ{��DP���߽^R+��ֶ���m?�� mk[��ֶ���w��&�HH��B����L��g ����T��

~Η�״z�'2�ݕ]��hV��7$EP�}��X?y"�G������s����!��bN ��*�@+�=~(��m���B�ƽ{'���[y�~V\��B?|(G�r~y&�o޹��H>~�#��eu�[��+��ۗ�Z,��H���Z��k�w�?�ٔ : ���ߒՆ9���r��7���#����ׄw|C�M�2a (6�l������_��ُc[���A*�Ն�}Eu�3�	놐�K���qL�k.��E�QDMU	n1Z �rCP��.3�͛�T�?&7���_G;#Zm<z�t��#�����n,Sy����x��-���r~3sǵf�g*�B�D�ͺ>7�lt�	U7�{G�W L�dI���QA�r�3t܂Տ���s����C��"��>�����ɏ���_�|J���We��kˊ��b�PA�c�����XF��� �����L,� �������������Y�9�	�Bb՗IWC�i��K�Pވ�$I'�״f)6�'��X����@3T�V=��A�X�v;[0�4+*���i�+8���픖����GU�"�j�W����`����$�f�����徍�(O�*�ͺ'�~��z@�`t�!�I�Uc�F��*�W�u\�X ��`�*xM�(6+=H�-p?���Nž�,�ÓVi�~�Y$�;���ow*���VP(��י��->�Y>X�V(n�S4H���H�E�E�\�t %վ��"(�ܠ\o(& �s���4�#���N���󊊛�4�0��
���C��s͗}��� ْ{�A��v�j�!�a=g�*^����O�ċ��*�߆�7U%���2������j~>�g '1�Q���k�f�%Ձf�l��«��3q��[�&���j6��� uO:� ���J�E;gUO��ۭL�Zb6E�
%��!������Q�0U�X��:S]؅g�Į^�6O��g��] �&in6h�)C;Ȝ���W�c��@sKI�'�_�
@�bо�1�ڐ	����CиYf��6��H@4����j~\N��ag����W�;����ٯ S|0:�n|�~C�����(S�N�gLa��Po$��F�Fk0�w�G2_͕���h��u��Z����=��|J7�,�u5ݳ���*S�|ϽJ��G���tC�9���5I�6-2���+�]�����t��	-Gq�s#�~��c��#��}�^��|AVJ�AnR G{rrx #����sJ��y���X�0Al���C�%�@~�8�u<���lƐõp� �z}��B8��X�O���N�VK��vK<r�gw��}G�5��"��ϋ;���W!}��h���~s1*�0Y�V��#��t��x8v�j#y�	�� �%�(Knf�/�lܻ2���������3^�''G��r��Ҷ���mm�a�� i[��ֶ��E۽Gǔ�òh8��d2&�Qde�Au%B�ӴCp���
&�Ak��}�O˫�x����$  �.���>|�m~��o�x�?8�%U�?&����.���͒ʈ�[�\�u�S��;���'?���>��9"�����������_��-ً��?�{'���W�÷߰����=9:�*��e��b9��^��~��B>��KZ@�>	}+�W/���ŕ[�?��'��̔�n֬�[�֚?��Xs �B��&���8o��!pꎥ+`
�-���t���y�/�7�kκz��-ѫw�}ج���\}��q��]�7�qZP��A��C \�o�������������O~$����pDN�����ɫ�]Le�ʸxf�|�ͩ�ZI�@=����Q���佼zAǰ��g�k���]����ȇ}@�Nd��8V�'���w�}'��{���%����<_Xh�(��HI�X�D���V���]4l����>K�oqDP��n���� ;Pm
���ژ��H�+мE�k�
Ʀ�Q+�:D��Z�LoqZP�[P2�`L�UE���J����Č�/��!��#�q�ݲeb��fr�<~��Uay���`��J6%JAbE�!e-q��FE�e��xk�U�1UL�j<� V���a���=!���`=�v��t(� ����Ǹt�s>��}oYI/�J�$��`p�Z״���ĉ�z��Q�7����y�BLEBd3�w��װ�����z;'�!�Y���+4/�W�W�,���&��y f!�JJ���^P�^�!WTeQ�>�77��%�s�����BV��R��"Oll�=9g�������kO���>+1zR� |�,�&�e�Qme������(Wuȭ��(�����諥*�|��;�]�y�-��hk�|�؀~�������i�쟠����уj��s�x�_�ݖ߷;���-x�ra��hr�#���kh{�y=Ȭ�s-2U���8��)_*O�p�����J!3�yZ2?ۀ=^h�1Z̙�
��q�y���{]ޏi�Wfj_Y�<���o<�p�vF�3B���4����M�I(P��<�=Q��s%VŖ��}��z���f5�E�de��{n4'�}=yO�L=�C D�YD�E(s'��{�����{?������,`�Bv:S���5&%�i���s}��FQI�E	n�Ȩ�3���z3��Ps7���X�L�u�o��HY����#��7&�����0�+��x@e� cH��Ђ�*,9͖.N4?��t#�*���I��`癌x/�3��jjv�+�ލF����z���3�۟�����y����	~D�luWErWr��l���]�$����ƽ�^]^�=���x�qD��L\�ź���v�#��M��Ѯ�;����kd�4Ԓ���������mmk[�~��%@�ֶ���m�6�E5[%㝱�P/t�� �"�~���f��.��4��~O� ������%�^_]��/,�2
��m�;��Z E�7�3����tby��\��I�-�w�"�q�#98ؓ�{'��}.����X��rr���w��<*ܢx@���!�n��WW`��]����Z��/PBv����^�o~��?~[�w`�7u�}yq��u�N�� 躥�ĝ��,V$B�Ht0�H7�J�d����G��wW$@|�+�L=A����-�sZ�Xѓ�>�v;Xlr�r��_ۏy�%� �6륁k�-��s_���y���3[^���ty*�߼e�������cy�����$������|��<{�L����F:�8w�X�\^˛wod�Y�^�+Cd�dVϞ��]O��kڍ��+���;�G�J���=t�ܿ_vF;����<_ ��z������_�/��+�h�,�q 6�k��v$0���@"��5r�r`��R�`<{���4On��D�@:���t�ſ�|8����Y�<�~����������W$*���XoԿ��݊Zx���Wɀ���:��:�#Eގу���r��7j��}̯\�!���}��'Ch�c���jZ�1 �KO(T��I&TV�ݬT׃V_vU�t$ü�F¹y�\#�'6@_���6��W�x5�m�����k%�)0�����=�u����X�܁��@�@f#R:��F��T��\���h4\�B�*#Y�p	UqV
��Xs�`)�lo�U�� of?����p{uvd�	P��T$�3&/�\���w;mr�����C�42P���e<'�m�r��Uƥ�� ѡ�- n����u��'��k�7l������HYu0�=�D�@�j'�d4ľ���Y�&��a&ET��{2�;��X�:U�͖��	I��u�dY�k��̟���0�ܹ�J(�Hk����{$A�S�����F@�W�6�B�g����VNU9�	�����qc���E��x0Q}�1j��yRQ԰�%�`٤�IM]0�%��'��z.��Fj�%�����jk���^��cՍ:�7��+�j�	|�6���Y���u�b�ةȕ4��$%�K��F$���Ij�	~�c�=c�M�2������ݗl�2��ƭ�m���n�U�6�{�X-�.Q4�p�����fz�����tG��E*2z�rq��x7�9�y[�����;��:����p.��#�O�g�j����y�p#���_B̦�5���l#����b t�[��dc��8��q�p���c��Ľ�*N���C���=ئ*��5��%:"�H�;&Z[�f��-�fz��\�cB_¢l��a�b!��0?GE��E�D�`�~�y�Q5 ���L���x�d�����b�y��)��}���w����n]'����i�%�k�}Eɕ?U�w����w0��o� �gg2tc%]7wM��]�Ay3O8Ǘ�#��h���]�߼�IG�ۑ��nl���)ZH��ֶ���[K���mmk[���-] ��P��5�,�h �o�4i�`s��d��@�*������*��Y)huQj�0��ݝ	�C���w;�Xt�ϫ�Ky��ˎ[T�iÄe�s�y�:�b:���"��痗����$��[������\O����V� ~�֊F�jFAE��7n�6^N��>����]8tHU��3��(#�S��bN5�t�p��p;Cyp����P�0��^�`��tzC VX����T� ����lJ�����k,`��C�!S��.LA��0�����}0�1������O �i�2U����A�s��$B��o�f�;�a�Sw~O��-��@����Η>@{�����tb��m�-4���������j6�f<��y]]]��;�i��d����X@~=z�H�?z(����v��Ͻ�1���qCu�
�տ��|���$? L�v	�M�7υ*�(� f�e�L[Z�,������E��ďC�>�̋�W�j�x��\�*�(���J�Op^e�` ��yI��^�M��n�,K���p��r�0
 �4Ң�"������NFm�"��m�A3+�O̪�g4�?xPH`�a��.�o����j�3D��p_E��V!��w�YI� �3P�Ԟ�9T�^	����e��}��V�[>R�A�TfĚ�]�VR�%I�ت�E�|p^��
Ǵ&T<i�<X\!c\V�)0���+�1V�Cm���6��Bavw>�^{�2{���\��̤6�'Oy��0Q �VX Cm�]q����T�B�a=��5�ǅVE��������J�ZF�F���a�>܇�7ǖ�ި>�lJkB.wݒ��3�G�ub+�N���l�Y��F�
*�D�Ĩr��,e�y�݆��)u� �l����*��_>�$TR-��e�D��>�um�?�4��[���p��X�	haHOr�܂��G���� %m�E�Wh	ß��*؆<9l�t���I�D��W�'�]'e���c^gb̖�*��Z�[��(���8�HI�@����D5Rd+�]� /�G�G���דǖ(Y��ׅ�g����4?�"V���gpaM��D��T���h����{gJɕ	f^�]c(F�3s�P��3�\]�_�w���\�z��p �v&P��wa5	�.������|� WͫI����p=_�ҽw�i(�z;5��h�i��g��f���0�/^���{�
6$c�Hz>���~-_|��-<�{,}�;�v]x&nJ%�@t�=��m֝�(cTA\��֌����ɕh�6���U���ʌ?���3������|����wI����]�?k�U��a����Y.rqs�����=��׹{W�k���Grt��ʞ��y���`�&������Bl�����̳Z�mmk[�~�%@�ֶ���mU-��$���;��
Kk��ѿ�K��E-�d�ʆ���^	�[�B�u�kw�G�{owO�JA; 4��sZ3������8g:�"�rlGE��QU�*Q�
�6���en�3��������
V0�WKy���m ��w{<���3�jM�&��$��r|o_N��}����.���@.�?��.����ײ�-�Wp0��<y�D<zH�����y�F93�lTh��X_/i!P�}���)p�i��12e�9��KI�1��Ǫ���F�"��j�H� �5������*�*̒&�hv���W�W׆b!ݾR�`u�&���T���+������|�ɏ�}(������yJ�.����$*G���}Y��Њ�- 2/߼���o��P>�� m@��X��;;c�/����7��Fá�������_�Z���ky����%�M����K���a!�m60�w�k}�7s?��Ze�"]����db�r�ȗVR������z�� Cej҉j0݃���7p�8����r
|�LnZ� ���JuE���Aa�Ζ���V>A 6�"�>��@2�C�˪& <(�h�[���(���?�0P�x�Z���U@Q4·$D�W¯��%�cp����u: �4�q��b��ʪ����{iEV�_4��dU����U�]����l-��ھ��}���Z�����@�#)�כ�O�Duſ?���Plh�oNBF|`���
�y+>[E��`k�T���S��޽n���@k�I��h�hC�J	�n�!*DG�f�@Y�cΫp�Z�<G���`}�c�U�$�����P�o���M���m��4R*�3'E�g��>�+8��?=�r�yb��>IC^O��F
��NY�*�*R2�IP�m��24�?�ꩩ��	a�S8$�e��<�� �d��[u5@��*M��ׄ��@04I�f)�'u��*�I��j�A�Bi�,+�5�Z���4w��*�(o������Ƽ�m���^Z��w�a�.���KfY4 xH��3�%t�wPչ&$��}N�dD"u|g)-�=$��s!�
��&4�]��7:7��EG�~�9U��O2D�u��Ǐe��J�������J,���w��k/!�۱>�v�e�w"���
�L�*�F1m����������avr~�2~�A	�>����˹{ֲX�jn���*yK���nLC@��g�r~!�#9={�y̜ʨv�j�\�o��3�<��S�q,'�,11�Pz^������B~���Խ����p�Cp��|�mΓj�}ۓ$42��QlVZxo�}k����+�;��d�Ղ��G V\�^�y�~/
�|V���Y������������/>_;i}O�՚4UU��6�\���>����N�Ƀ���u %������z��5��?�G�b&��|��λ��~�˰�;�KZ$mk[��ֶtk	����mmk�_]���5@�
��v5 >����tN��ٰ���Ħ`�A���>�V=�~�	��p����[_^Iy�A��{Mƴ�XBiqs�
���{2t�~�������d0����[O��U,� ��I 0>�s0&.�����Lz����nA�k�I?H҉eoo�^,t����O>a�y��l\L�C9::�-옖�2X���}&�ْj�ǻ��W>��v:}��Bf�%k�UO��T�7Pb��H��U�g�)R����۝�ڝ�x2�+�seVE"$�8.�o
����Ad��� K��~L�DR�� 7� J`_��A��j)?Pr�?�Fa����C��Ve�8>
�'�d�\�L�Y$P���ep��Q환e�o8nx{c�y;$�s˷�>�_��W�o����tn�စ;���f�@z|�G%�4rb����0�1JB�DH(H�]��D���Q6?k �Q�W(�
�OuǱZ���Ra�c�On�.�`��ξ,n^q�0O� �$�W�3J�ݾ����e�=�,I�#����/8IR��I7�A�` �=`{Xٽ�e����"#{\�����.^]�"2�d�ǝ��~��{d�@v�R���舌xϟ�����ꧪZQ��]�-�̤=�x�{)I�(5��B+"�D���Ǚ����:��Y=F�m7d om�d�ɯ�Q����5�kWœ~�'�o)ρ/�j!�٘*J�}'�l�Z7�哷�
*�/���v{�|��Y�ʡ���BU@�?aaYIX+�H~X�'Q��=��X��x`y-Jਏ��+p?��BM��r�_=6%L�~[��k@�L=�E�I5h�:�k�+������F;a��,�>+�o��a%u��<P����5r��E,�I���^��n��B_��^)a&/��q�͆hj�M��@T�������M-�4{�׏�k���-�}i�#	��!��c��u����e��0R2[O�+��?'u?`��N�����nq�)j�m6W֩J|I3.�aZ�6�U$$�|ٿ���}a�P�J�'�-�^1p*O$�@f����� e����_;״�ù�̫=��C���b���v{vNrI���|.��+7�W_����x-�~��{��`m�����P�����ڞ�%x��Tj7(�@�����o�ey���Ϟ�yХ쯏i���3�lO�М��fئ���z���3�&,�~ǽ�L'P�%������Q�n�vpxH���oQ����K7����5W� �5��=Ȯ+���j#�n���dq��"�����b*uз�����sf�@����	�W8v�f�.+����.����'��Cy��;����5ъ.�|P���*�^�"U���ȧ8#\����`�i������ϊ;?k�i�I�$�*z�����H��t>�F0���88��y��2Kk������������3�<9v?���{}(���I>��_���"e��2���s�ƛo�9�+���x@�t����,�mo����=7Z���_��k]�Z׺��nҵ�u�k]�q0E����@!8��|,@�h�-�J�}�jT�cш�-TY�%�ݤ�E��/r/f7�N��?���[�^\��� ь��-��ѣG\o��f~+��%��� �pus-�a_��!Ȕx���ۆ[|��o��E2j�]R�[�0�.J����%�$,ޠ<�t�WW�hY���y[����DA�9@��֘��Ӟ�<�l���DQP���	tѮj6W0�~�}�	L�?���z ����i���B�*�؇ؼ߽�rlU�u :�zP�o UR��Z�*�'#��ؗ�fe�O oTuS]�"i�9U��3�+P�y{+/N��`��}YI2�L�g��M9:>��]Q/c����&1P 	|�A~�YE��Det��0+y�ȍ�Jn��I�a��&'����S����믿f�H��a���U�@�`��RG&�]�-,>`pvH� #7y%����;vC���-�C�A;�A�0tlX�J�1����ޞ<q?�q�1��)L̞J4l�b��juV�V�Ъ���ܡz���x��Wb�ڵ��r&���DZJ�{a_3X"�u;�ZĘ�AԖG�Z5�J�aQ�3����M��&���woM���{��$�*�4\�ר4ԚD������/(�a'�％�*&�?�m�k��*H�:��3$t�0�AiZN�j�d�rf�<��(�mP��^ �1��� ����@��f��]��:��:�"2�ӦP�ҧ4�6�ji���w�emx<��;���.V�'h���l	˭ ��f����'$�������^���uTf
�H�&�A~�f�'͹l�����U;��+w8�MA1G��@�'!��J�/�� �UQ��]��o����.#��[(9��׬�����VU�\�ϧ%����yo{ž�5a�8�Α(^*#���r;P[H�1�{�)�<��I)�%ޖ+h�U��-�<�VP\����=?�ǡ��ա�>�k9����>��V`!T��yu����k%F���W����^��J2�5F�����zi�?aa��&����-���fu�I��V �&�����aΓ�?���g��9 -E'C��\0��x��y�I��J8�z�wi9���&CU�G2���T�� �q`��,W37Hv�<p����6އ��TJo�q����r����C*�@�,����ibwk^7P���j�9v�~�q��L˫��E�^]��n�-G�T}n�n���vd{o[~��_�o�'QĢ��Ⱦ�<VE(
t`��ip�|%�})�sJ�^�Lwvn�N[Q�g�9/��@�:T���WM�D�>�+a�yw�� �����>�s�7e$P�(��Y7�W^������r���t_����T��տ�K�ş�R��6�+,ը�1�s��E�1����F��n����}�NG�����F����~=qo���������t�k]�Z�~��#@�ֵ�u�k���ݰ��Ǭ�W��S��+ҍ�og���#���}M��Z�z ���Y��c���!��� ���{@��@�1�L�`�����Q݈/�I��c�������x���r{;wߗTv��ۨ.��� �s�h���h�`!A�HC~����,KVD�ӔU��0���	@b�;���s3�fB�c�������q��ܔ�hPC��Ox�f�v�v�T\����ld|h,HV�n
Y���`�g6�Oh�6�q���hu��_�6H=���!��7j#��V��I 8�i�,�.Ci��G�U�(	BK�`h��B�@Q����4����$d���?��;�		�H5@b����
�ihma�nPjXm��/�x��VK}>;{A{�� ^��ʋg'r��	�#�-���+�+�7��Sc�d\������l�RT�Ar�a�@���� TeA��L���9r��j���'[�m;Ǜ:�!�p]*�̳_���X^��~Z�( �F�@(�V�y�x����&Ȕ6@PGTem'�Ϡ���Il�U謀^+	�c���ܲ�RR�T�K�!k-;��lr	#Po�S�v[�3�n����ʤl��=(�
s�@ef-�j;JjUF`@-�ನ�Q��D��x�d��o�{Gn�m�/Qh�zF��+�¦ھ&����:�)͖N��2��[hH�w�"a�B�K���,�P�^(Sg�_�j�h�<Q��r������*�+��o*:L���e��)m�"wݻk�	�Nޤ�3s����(��K% C���T ���>W� yjƾ�?�C�yL⚐�c��������~y�{��o�Ӽ���T�T���_�~��-j�ھ̓��M���x��k���k�M<h^E�d{TM>O[�D�E%iJX�,uϢ����������Cύ��jZ��QɄUP�&�[��V��!����ʍ� �U!�5�öY��6�ɋ\�Ԙ�!^�׿Vi��C���_ ����T��~�����)��{��{�	��%sj��\��Gk0L�9��s#��Y��.�n2�I��fP9��?� (�V�� 3�"����ô���F����Y��2*�y9�T� ��
��ݑ_����gT��:�s�١�c!�{�b�\�5q�a�~�U�q�,k��J����K�>E(�}�>�|dU�|��=����M�Sr�kzgoK�3��J�}�����#;�{?WWW2ws�
֦}�����+͗)�	(N��=r礧�(R�
��&��f����s(�xM����)m+��(T�Fd��,��Г �T�!q��=w���H�}���[�"�&3��I�1-"f�e���Ӳ��^���;��|�����h�s�mVbS�iw�׶d��}t�ޡ��?����/d�}>梸Ƞ��ǘ�-b�o�TȰЈ�S�D^.�݃����w}��S�k7��YP��k]�Z׺��mҵ�u�k]�Q�x�����Z&��!� =�6���"���ݗ�r!n�uG/F�h� 8 V��lZ$�X̮hck�^?����ō�&c�h}����?�� ���k���t��j�"�����v!�=���7 6��k�y��	 ��΀��x<�M���V����l��\�n$��s�*J 	���2���x�8������r{}-O�<e%�_���w�}O���
3uٓ��lJ���U�QH`�Mc�V��#P����Y��	�����
����v�3 ���E}��X�Zȧ��X,�|U�5�����65k*��� _|O���i���q�J�Pŵ{���'�8�Tm�?|�~%�����t�o4�f � ����\B����x�T���ɓ'E}���@VěO{��kO�H��H�E9��j�<�V�|�)��MH���gx�ׇM���[�Uɋ���d������I5T��ڦ���zMeOU)��Ph5�G�$&yUR��`+���~f`K���� hC@xb�m����x}��k�	Tz(��s#��L^y<�Y�l���	�W;x�U]ݪto�T�T�Ym58L�m8�j�J�&�Y�Mv@M~��z�H	V�9�4T����U�׶X�^;$�>P�����B_OK-��`}0��ᯩB�͓0�>��_�t}����r]��� ?_�KjrF�6�Z�Ϡ����Zq�@��I����֐@	,K���y���)���0l��&?����/�J��Q <�*��K38̦)W��ɘ`y�0��

;.oGUg�Mм��(s�8���<����i5OL���GQ�$w��Lll14�H �(�һ�hh�i��i!W�v]`_�+�ϑ h��vp�{E�f�F"�[��@�Pm�|����[��Z��i�@��*S�:�$�xV^�����H"�V�j��_�\	�>�ם-��z=T�VhE3ּ��?��z+4�4W����0Và����_�dF>H� ��3�U[�B�|>u CaY������T"���L�{�|�Z�̇NN_���\�����6��;ȿ@H8��R�5�!P[���;���{8���p��eeF5'2�0�+�@���#�C���l�Y�,+X[�lOM�w�@��qXc�ݳ�:�Ԛs7gB��`b֤U�����fY:��l�Œ����d���e����~	U�x �`���^N�^��t}��h��-��
�b���&���6�Z��nN�9^X���,!j�x^����iO3A��;��΋�;�E|`���h�5i	��藡�XR��*
H����_�c�V��a*��޿X�TQc�������<}vzW��g����z�Ï������!��6A-Ö�G�A8��7����E��F��k�A�f᠗��{�O�����n�Z׺ֵ��D[G�t�k]�Z��U5���`@L0_�'ak���c.$7n�w};s�7��^�G�{2s���,*�^]sѺ���y^���s����,碯�.�^��PR_V\���
��]�"XJ�Jb,8zp��"mwoW��Ƀ���}S%�?5*���Ɋ�W�\_\\��ǏYٶY��"\�8�M&O�<c�h�K9><��o�V���ɷ�~%/�_���ry�J���e��h�	*a���k*��l�L�ļХP�����
(��O�b��3�.T�`e��P ����%s&
�ku��!UN���Y-����>�mU AY@@DX=�b�-T ���
*_�;;i�Ϯeu����r���-�߬��6�<"8��n4�p.�+��P�?��p]���^�g��$�@<a��x�%r�� @�Bx���{ 7��=�.ii�y7�n_�|50������#R@k����[vB�P�lAF���XJڌ�� �`qC��Z�E �AD�A`l��{y�܋c��i���&2PZ�>8\Q��jo��|��j1f��j���p����*�p�R��*�5T6���ٕ�+�r�$����UM��?����Ɣ	���9\�bF�]���̰}���U���U���@m�²��׏�W��|��J	Ci��5\3!������J����� �?��;�~�l�5�t�ر�s\��tC��+�J�߈Z����,����_�A����m�ڤT$]�\�7��$�"���� s+��԰=�z߳^��
�Z�fW���ؽ��L��0���4?Bn����
�j�"�P���+YO�RϬ�(@j�?d��,$v���#i�ʱ��!M+@w]b삀/����ߧ�3�8�$`�{p����j$j��{�'7�0X�$uP�f�-L�$�ģ2�L𤃞c�� h�%^TET,�C���y�ā>������pu^]z����@{8\fI��ŕ'=��)���?��0�ۏ������Q��,����g�RӬ��x�����P�~aM�����^Ʉ9�]'8������q�T��Ɨۏ� Qe �ZE��B	G�#|�=?U2��lgO a>��E���9�s��6~���K����z�ꏭ�V\Dn'���7��խ,s��d�͍0��0��g�H%(cΑ`C��G���2 mx^,��q���X�?�ǸWS�Q�enh�,-^��Y!P��%^�緶�ʫ޴ǟQx�Pu�'d����*U9UV)K�Ƚ��m��h��P#��G��q�m8o]�yJ��yʦ�x�Ǯ_0^�eQ[�i?'j���TZ@���L���6=��3W�{�̈�2u�`�IA��Z2?��ī=�0��A����'n�{|t@B�����1k�o/{}s)��Z�ᾲ)62��=`�rO�É���e��l�'W܉��X[�ٌڂ��P?���{�*ݸρ2���+��/T3�G$<0&0��1�v���c��;����^tr�=�}'A��u�k]��O�u7��u�k]�ڏ�2�����DK�	�[������껳�+�)�����w�ʳg/��� I����[,���S��EZl~p��-rE��g�r�꾌�S.���B���[\e��9C:=ڗ�lF�gdn,�_�i 0f{�'���ek{G�޽{$+�@%��G�h_ Фh*aU钒�9}�\�맟ʩ�������������"�g~$n�&�ړ{���?���,_~�|���rx{(��AT���WYaV:%��=V�����. h�}^�s��a5d��}w (��n���������T�m6U s�r���W�b3DT��0��+ ���=U?x}��j�R&���v`Pb:�!Q6[�d;�24���|�KTFn<�o>�B����w ���Qw���l���P��ab!��ߺ~��=�%6�o�3څXހsba�b<� ��0P� ��/�K� �ɊU؅;�!=�QUIb�8�mY}�d �R�&w_��?l7�P���{�,E��\/�(�퀲M*K� vw����L���������D���f&���*�
晔���:��Ӗ	�&�]���tc.m��	X�dmDfM��U� �Q�J���n�d�R��>�A��̖~e�
�b�2� ��Y�d��^Y�2�Zyy�-
�T�Ӫ�}^;��pРZ!pj�Z]�ʉ(�j����Wq?A����[X�Jv�����f��3T�ՕϨ��#�O� �����4��֫��i�pem/lSeCIB���_���Y�������6=�f��<!/B��� ;,dh�U�=ɻ���d�$|���I��L�wx�aT3�Hr�/�Q�lrr�)E��Q���f����ޫ&�?�c��U��ꥷ'��,���`�]�uO�hoǅ�JN��@3V,g ��7$�pn�|�=$/��A�g��%Al��@� �!�����7�ښAB��Hl�83\�>ͤ��Dm���˔6>~��Lo�'$�-��p�0�ףo�W_�JB�7˻��M�8
�`�m����l�BS�x��Z���F�s�:����m)��d��ȶ���U=R��l��bͫ�x�{�l����>�H�����Yp�D�Q�@d]P�>�w��窄�����J��>��O�7 ��>�I�B��	��BQ��@m�r-A��:�].L�!���`w[���(���=��r}{�=�@;�7T=����,n�og�܍�'rt\ȑ���P��6R�g��X��:[����$�j����ː��:q}������ �'�'z>T��@��xU$�ї 4� +�J	Ǿ����)�}�pIi�;O@��CޏT����ǈu��a���+�uoϝǓ�gr���en�*w..�.���7��'�Yn44�]�a���C٪ps�-Z�b<�g��>�R{6�%���BU=�r����Lӆ�B��|�J�������CZ�wh0���D��1���s������[������#�5,�e{Y���T�%w�f�|���n.�����]�Z��*�W7)�37���NO..�f�Q�!MN���������x�@�}�]�;8"Ѹ�����qϼ�|��W���3>+0����|j�{VE�9�y72D��W#���;�{A4��^<��b�n��H�ֵ�u�k?�� ]�Z׺ֵ��,\ �m:"�u��v�»�`uvqA0o ��-��d���؈[�.��{�}9
��yk,3�Z?yy&�ѐ6X(��R`;�l �;;�2@����������%) � ~� �a�ӭ�ʽ��P�2p�1�Nj �g-�*i*P�׿e���b��?��H��]y��[y��;y��[�]ɋ�r�g����b��=�>�@�����8cv@4Tӆ�P`iU�*�=�� @	�Tem�¢YV�j5te� �-U����	KV��pW�C  �$G�j��m0��Y��g�}{e�Ym�����sF�=�E�Aª��9P��ơ`<�iمj���X�rۅ�c�ۇ�U� 5�E�6"Z��@�f�Y+hp�AO�É,�s���XEΟ�Z� �*�1h}xV�j�G����V!�U��'��-u�����{,��������#7P)!�
��j-�x���G˳��g$��>��1A�k }�s� �J��+�	�:��	�J�l�m���-Ն�p h	�	���������\T�z��4!,�&4�>�,pK�O?��&���>{��e�@�������t��6��x���y���$��?Iwr��̂JϹ��,D���|�V*���'fA�YJ�ĥ;�`���*In��$0P����OU鐈h�ڃ���EX�1��m�]�U�9~ime෿���r&�k��,W�����S���T8bVQ�*d�H?���f�z�y �v���H3��$R�B� �
��s��Ԁiغ�c��G��R���=�[V��~I��2U[��G�W"$5i���V,�,�=�C��S�#}���]�ގ	*@���ƴx3 ��cQ`䁻g'I��/���o9v��(B͉��Ô��Ѽ܋Q���DHv`�ln�i��:���\ýܬ)�v�X��9N̺�7�fժ
�_���{�'�/�v1O�wl�Ji����fE��_�i^�E�W}�W�n�^� i
�q��}XH��}�����5��*��>;�?LH�(9����e1!t:ToϚ�-��E�Z�GmW`�Ii�z�c��rrP����%��Z�ThT�D��P�|���Y�����O���n�����{GTL�x�L"�]o�}~����q��gn��aLm�����J������}_  bsB��������|8�������&�_(4��K� ��r�p���5-ZH����v�P`A���MV�9���T�%�C!:��i�9�|~+_�<{�[{;�<_�n���_�ɋ��������*i_h�[\�[nNyt�O���r���t:p���rs�����G��.b�?��y��z�๎�CP}4Wk3���
7q}�b���-�|������#����+޷�e�̽��< a��õԏ�<' 9�/�z�o��ى��?�Gy��Ϟ<vs�[��9l#w�&T�����ܜ5��d[j�W�������s���t����\>��S9?}*�/_��م�ܼ}�X˾;ؠ��z%/_�\F����J+��~$��TF���y�X��#@�ֵ�u��:�k]�Z׺������J2hWhoܢg�<P������#9��P�D-�L�H����)���xB�$m�,u�H,$s�sU�*Y����X>���������j�d0�;;�rssK���+�|���Fn�z$�x(�ǲ�\�F/`Ѱ��RD 1#0�ŰV۩�5*�Y�� x����-v��o�F�{�m9}�X���s�������'nQwż���ͣ7ߤ�Çi%�0���xC��.���܀EX�-�4�``���`��cz��� `�����K�s�Y�����H+����BUkE늲���^�em#1<>�>��Te� �Qi�~C57����b�[��g�]$O��^����Ez�S �_#�~N�	� T�g�a�a�Ѱa�"p�i� ]�2U_sb�F~��]2DvF�6V�[7��2*=
� �r6M�-H?;JH�r7�Bj�ɝ�΀yL%��z�c��*�K��.���g����G�������+^+����j�Ъk��D��թdHbO��5�� ��s'�?��	T%9V*1A��H�lN/b�8C�A�#Ƞ���k��@э �g����8�j��C�I>��jr�?irj�/)Y���Ѱr3a貴�=dRX�G�Z�@�ڹ��_�VN��k[sy�oA�!Á��+`���m`�7�'�e��V�j@|�=�1��q��FP�̈��61�����y{[/�G!�ZOB��_�Aw�1���X��&����3SD�mV���� 5�Ix�k�E#r}5��${�|�3;ځ�UY�ش�ʍ�	��b,��gP������ϙ3@w-2[�Y1��@&�Zx�ჸqNro�%��2�~H�4@�k+eN�LF,�Uc�>�v�Fwn6������r�J�{��l�N�L\�M�m[�s��}���G�%bN�"�9�cGศ=b䭐���J[�_hNO��qҐ-9_J_���+%P���zxB�l!9(��V ���bS�X�3b1΍]H�R�}��&�eVb��F�՛1�ʘ�n+��<��x.Re�6�F��I���kV̈h^�g���nx���zQ�{$��U�ٓ��6�����\^�����=GR��ݓ�n>�m&	��y�dgύ��e��T���n^�T�_�r��� �C�����Z�=�G�	���@8D�H�
0ء�}%`�
��������g$r���gw�`���Pv��*#��3�
lWQ,3��q>	5�3���\]]�y�g��?r�"[��0�M@a	��r����}d��f��}Lb`����;�+>��x궥��v�����
'B+�XىƜgq{K%�v�G�Zr�6���p4���)����<xpO&����Ɉsy>�D-1NsΉ<7{1�#S7w��١���������[��o�Y���[�:��ۆ��{��$306������s��\5d�H����k<��e[�[�b ���<�<{.�?q�y#���-ܜ�������|������L>��w�?|*7ח2�-��ܬK9������;2��}�mI׺ֵ�u��:�k]�Z׺��6�� APa�"Lq_$�!ӽ�خ,�KV���{���S��_\������]�OB�����|2pۅ��n��-2Le��dG�U��o����A���.�a�u�꒞�����o�O�\�c����M��Q�~lHc��k[��E���� ���}��e�c������w����ѣG$:~����7�|)��L�#H�u�ux| ����/�z6g51����US
$�ڻ��̀`@�*h� �}�n|M����L��3[��������aBp���~i�4�a�~���� �{?�����S5��q|���=���@[�3l����� &v���%��g �&A�t�m0��s���;�A��S� wۀVV��eP$���Vrj({D�:U�I_��X����aր�J��e�GZ��~Ap���\7��E)y���T�Z!��jr��r���j��u,Ȩ q����+䱽��,IZ����v�j�z=�&ȸ�J���N'����f:$V�J^w ��_j m=A��`M>�Q�e ��r���+I�}��o̶�+���/�����40�����q}DqnU�v�-E��}���1.a�Ĭ��j+��
b�_�O�0��&'(H~�F�
���`&`���#�7h^O�q��8G��7 ��eD����o�&rૠV6��V5����^9����_��cƂFP��R2$z�f��$t���g��J�Y�uU���Q������EE����Ͻ�7��C��:;�2a��&�t?����U��wQEh9�*	Ay=׫���9�<�#��p�/V߳�[��h	���M���õ�x
��
��H��	=�,���E�92�i�	
�s�����o#g=����v��v�ٕ]�eC��W2@IP�k�2�2���-��Dj&�ْ�36A����►����,1�<k��+/�<-Lq!�5�n^�w�٘*�FaV�x���u�<���=IV���:���~`�7Kc��l�LY�� ��q���s�>l�<����5�b{V��ʨ~�zrԧ"�5#,��+�T���T����ٓ'��s;5s����+�a5Z"�-�s���ե|��o����?�v��;S%J`���=���x�0�׬����s��H\�L�2�
ދ��-������xy[F����v��<���وܹ��[`[ "#V��U%����8��y�z$���4u���s?ž�$&pPT2�]�q������6I���*r%��ĝ{�ϣ�s��7�RI
el�6J��=�?8�_��C7�ݓW8?'��p�"���D��;���Z����|	�@ ݘ��q��цk���=gh�e�6�"�|��ǲ��'���|��g������>'y1�EX�o'���]����c���;d�])�^A�`�����ۛ��_�Vj������Z������>������1�)_���{%`�𾽙s�,�K#4+�ᒄ�u�k]��O�uH׺ֵ�u�GmnqRUT�qP�eY c���r�Y���	>�P�n�6�bb8�ސ������{��S���\��<a5@\(9�Q������-zn����-�a��tꍅM����)_��p,~���
,Ƕ�{n!=�U�������ݢ�e(���U k,t�熃�a�P:��y�ǔ�u!�� f�&�+�������}���4q����>�M��3w�E��B׏�%[�n[�=!��l�� ��qqSAt�{أ����o,�	�`������X|NG
�d!�3�2qj���@��; ��Z��XШU#�&(54�թ�^mg��u`�=��ͭ���f0 ��-URآ���	�E��^���QBy-�4���e(�Eh ��U?o�타��.����f���Q���lk���������,�
�|`�q莧t��O"fg��wl�zc��ߐ�N��W�h���!�kbW���RI˞�W�r����<4=Ҽ�H��2�V,��g�*��G{1uH��Qz����薳�tW���1?�I%-V���0+*Ot��(����[W���ڴ���Z��m�|���k۫P�7J����>j�Cmգ�#4T,�m�zH�H%8��h�bʀpo���AN�W�p|�-���P4'"�E�z�{��hѾ,7
��a��j!�vT���0l��K�<�!2,��Z��-4�y$�WM��@��y���~)��X�Ýƪvw���y_���	��P�����Z����EM��FNR�ݘ��ekۨZ�c@�'G�
�l�jHU��f6�S^�Q�t�H�6M>ky8$���"�J*�{&�*@�� �9���}� �!	)8�}����:�KSX�u^sJ�5���` ��\�goUV���J��@����-��S�C͏��H
|.��>�fW��BmaF5Q�~�R�vk�"Hup�xrMϯ��kvd�OP�ԊE�N4���=�v$ � �R@H����)ļZ�D�uh��=�oDnc���X����d��}��)_�PS[!U:fي&Y���P4��Z�Xb�I���IG��jۭ$�}�J[w�)nh�yrr*���j���6�abyh	?[�s��땜>&_}��\���2a��|j��R��3rP�L�k � �����k�}!��Α���	�|�(nޥE+Y�fD�qgPH�7�rBfD���H�}A�G����&�KS'�_.�G`;�^O���P��sa|���x8%є�RLUn��A���t:���^/88<8��ji��+�mt���4E�E�vR|F��KE��>��C��_|,g�/�O>a�I/�����k�f�7�m�~��
�-ȫ�34�� �@0�L�Jv�ew{G�ޓ��GB9��鷪����;p��@޻'�W3y��\Yc�Y3@z$�����Y1n>��ͷ��[��[�9Y��O����ߗ�e���y��ޮ��/=�v7�N_�u�]����� �ֵ�u�k?�� ]�Z׺ֵ�Ű���4ǊȭDF�[E�T�b�j��h4v��������i����/��w��D����ރ{n�{��)e^qw��D~����
�Q�@ހd�nQv"�?&�E����L���м�x%׬��������=�Eh���)v]�A��媸R�0/�bY/���JddB�M���6^�>,��M������rx�|�������Y޲*���F�n���Ȥ'��y�����\˔����Bc8�R�5g�.�3����&� �� �6��������J�&P� �*��p)I�����o4�v��bN�������8�
ꄄ3J������իk���ގ[�n�6�v6��z�}�+�>X��w�J��3��,	8 Wd
��X�M}Å
�˛K�Z��}31r�go)<�{I�Lm�4�:���� [���=ZU��u_�ߓ��HA�k&K�7}?�_P1m}\������t��H.Ukl�@L��'H�7��!�$b�!��y�3��j�, 6@&��T�R��@��	[���i�����cZ�y�RJ$�J����R�༈����8 �m���>��SO��w�U]K��@����ݓp�ig����6�֟C
�T����TYղ�(M�T��=�+���P��B���l�X�����c%[��qOE`_����_V>��>��y2�۬�clL�]����
��s�ߕ*?JS>x��$Q2ԙ�ޔ�s�A�)g�پ��]���G�v��m�Բ,d��[C|x���x��(�T���Ͼ*k��C�7S�M��9��� 1%K��FH^�cI�Q+B�_^[Xxl�0d����$ɕ(P����xOb�:����8�=y
�ղk@-ǌ����c�+*|�k����֩���x� 䚒�[a�ǅ����)��4����u�m��tp��_L�H�ISl`��P��ܒ���)-|����hy��u[�[���\*�S���=St�����|���]�y��%��gF����Ḷa���$�~Nf�&�<�c~h
6<������su�B�2 ���Wn�`�Y�ƪ�r'=l�XF3���W�V�G r+P ��(
���O40��k�̃��������h�	EwH���|���:#A�^�8W�X.��� ��q}�Sv5��F�C]d=7��"��7E�����ý� ������B�*�S��/��;�ժ7!�X��1�B�P}F�Ԅ"�;��k*���"��3�q,Ws��cs O*ڥb�&������ Djǈ�������ww�n~��yd���Hf���8�=�}$���=���{(��*�s��ܕ�M�.�]`���a���!�W#w�������"�jm�Y [�#7�ߓ����Ik+,��xs�k��W�>r����},�}�--�@�?ps��}�G�6�t�}��w�pw�V�'''���� {n����ͥk]�Z׺�nҵ�u�k]�Q[�i�u����d	�J�u�Z-�b怋���=.����B'nA7��e<��n����g,q?�A�,'D=���|�ͷ�F�Ơ?�75*����嫯�b��[o�%GG�n�.��nB���H�v����	~��k���ʫ�z!s����V%Y���$dU+�K �醯_,W���}4@�z�3����ޒ��y_�?,��.�^]�HX=�
���ѡ��h:���}��TJ�=�8��W��II�z�(#�<,�  k�� ��� �r���?��p_��!���sV�M]_2�:����X� V+����E+l��N���	������@����HH�`�j��2cWv�^V�@
"�p�I#^C:Ԃ'R����0��a����������FV� 9�z��U�g4���������x�z������PB��!���Ǆ�9�jT��@������75	C��F��y�d���P+��"�a�6�!�?$�%��:��a��ǅU�G^55����P����61���l�|��	�7��*�C�;^Kp3T��6�w� ��\/�xe�'M4#��U�sVЕ�H�O�E��������vz�Z�6>�D��T`�>S�#�c��*)�g��y[%��`��Kސ3�n�T��FǊ���M�|ܟJ%Բ�	.�D��/k�s��`��'���VI�w�'�ZjOf�9VSc p�@)�p'�P6�_�9(8p��ʑ��"��R���O�IO8�u�������
�k��@;�FR��Rv^��;�JjoX�z�����H�-�XA_p�{�.�#O ��1�59)ؽЬ��5Q�u������l�e�'�!���ꏢQg���`��k�O@�s�a�_�3�@$�:1�5|v�t��G�u����T˞\sOl�V����W��ؠ*�
��z+���q7x=2�C�mO�j�F߀"���^�U�M<��¬�`�����r�[�*@���z~��5d>GUŕ��QcR�Q/Rr��{��>�/>@���}�e�y?w������f[��	܏AI/�v^]]�˗/��e�Z�U9G?T ����U��T(P��x���h���T/��X+D�S�o֒������Ȩ����m1ϩ�9l+�D)��8w�*]yƊ�JL����Qb��c��# _�2w�A���̱�k)�V��s����PW���gF�FJ�VlB��	�X� ��q_vw�H���ue�y/�W�_���z��򈶕O�p�B����q�' ?�wewg��ӆ����a�H�8*8�@�տ�̨r�v�8.�N���J�ϖ,����آ�sE*��f%Y$�T�
� ����/�>��7��쥼p��Mfk��;2�w��!A"a!΍���|��_�ߐ�֔j��c7~�ͅ�Sݽ� [;P~$�H7̣��x8�w,�:'���k�E{.�ri�vs�̮w���d ]�Z׺�Snҵ�u�k]�Q[�W��ʐ�|�N�Y%���*(������{/��/��-�)��"� ?�V�
��-�7��&��uc���x26M��GE0$�o����E�����z+�� �dl�{k2U���#�{�\�k�r����Zf�9��_0��<k�Ȳ�|~�"c-���W�9 ab�JAT��WC��E�s��1�{�-wv�ݢ�m�Pu�ݓL^]��H�������ށ[�Q����s�8?��1�b@ �Xlij*7@5������3�����Bf�[��A�GΒOޣ�Q+�S��¶�h�6�&c���<�����,�c�ۡUF�p߬��±��(��`K�L��b`�k�ٌU��O,��>���VZ���j��X�?��8"�CK�2��Cl�	�JA����J�RV��Z@���;(h�̶��!T3cVY4�r�J�h8���+�f���vd��p�JU� #*�+Z�%b�dE� 5��,g�'Z� 	��A�V)���O��kZ��;���럤?� $��Q4�,�M��h�*ZUiM����@}��B�r3�8	@@{͚�*�P��%��}�T�KsnD��q�E�p8 pIk,`Gf}T()�*j�Ju�=@��YD�o��I�Gj�i=׿����I�g /I����U]��ݑ�VG$=6F
����W���d�"����WA�}Ԑoo�����Ѡ�P-i�����m���(�Z�A0>h�[R��|@&��N��aAmq7��+j��Ѫ���v%�А��ﶕ�@�jB���gt`���(��L�{�x f@x�3���,�������4u���x=�h�^��weVEނ�W��=�K_qX�w����`����{1�L������ap�� �糶u��=���Ni�Ԋ��9q
2`1�O��hȆ��r�'U�&��^������洛��|?�:�ׇ)ju``�����r��<�^��W��D	��H	*�h9�J�:K����d6l��V]^��)�h�f�9^�R�@m�BZw�|fM�T���q��e�'(������6�����7��\��"9[����9�z�|�GZ'�+��m�0$'�� 0�D�%��E��[H���Z�+�ߖ��!���7
+B�g��j�������37gz�"
�y0�A�D¼�+�y�5��^b��n�T/`[����`�ؓ>�z�w��;���7G���C�m���:���R��S��{ yݵX�+#N#��Sw�!@gA�9�	�%�:�{U�r>��x��0�W�OC�lG�ҀsL(JaÖ�[�������"7�Eh:r�P{V��c>�}Ƴ|oo�jXf��C�v?c��7�Ts����D�N�Èy) �&c5�x���d5S�p�]�c.Q��f����y�ö�y�rZ�jU��TW�_$�����}EH�0�\�>��6�[�r��#y��-w,k���ݜ�]�E�q_����kNޞ�߫B��/�ٳ��>xt��5����_��ƣ7��oPъ�:�nkkǝ�9�w���p������d8���{]�Z׺ֵ�aZG�t�k]�Z�~������}�����*��_n�,����!m@>�^���������V0RC&gWs.���a�W�2��e�",�>|C>��C�O?&`���êET퟼8�W��d�u�������"�6E�|�8J� �Z��R��e��}lþ�f����9�AY����9,oԃ[��(�q���ɘ@�b���<Lb�@
_,��^��l�`*�@,�3;[[n�7������}���-��R�Q�b~s='���~��+�s����9:���\xAQr�=��"��n�����W��2�Y��uL�j����<L�],�w�	�J��;^�����4no��E�( �\ ����
��`�u�����o�nF�i�q�
 ��p4q���z�{/�&��
<�Q��<�g�qcT��d�L  Cr��ByF�*zw��J�B�`���q�`�B2b�X��$A��N/8���$�hM�<�	���,[[��U��wz���T�l	U���
�$X��%V��5Aq�/��� *�f���ޚ���J�j�B�`���MA�+�v��I��?֌�!$R;��}�$T�TU�o����eQ���J*6� |�]b�%�K������O��c!��'A����$�k�辀$��RD��*Zb�,�"RWҫT�f hM����h �iۑ)���n�>�6o��&I�/�����L����3�Ľ_3+�2O����x,$�2���/�у�a���. �q�|b�=����!�>�� {ـ�m*i��8g�:�l}Ώ�oȌ�aKdv2�Yr���<��c���e�1��q��OS�5��l�����+I�F�n`Ie��Z �ˑ��g��&�� �pM�#��<���p�7d�@��C�@Y��$��̠R�P��L�$t|F���<���6�F���d����a$�u<0������@XB)���e���YWj.Iny~\���&#�"�e@��;�m��*7"�Kz|-� �ܢT-�p� ��!��q��pm����'�\�������]mx�l��W�z2���Ѫ���aK����Vo���0s	�S5a_'�SS�T$P�L��*(p6���%�e�((<��h��k����ff�2�F��P"�O�!��`��W�	� �ۙ�U?�o�?���{�����)��U= �)�#�����VR�R��-���+7z%��)�I�}�-�-����|E�o�n��^wy-׷���s�}^��,���i%7'ٚN�����|K9y����W�~���Δ�?��|c�g4�w��C����qo�l��+�?I�dJܟ�y��b�\ռ �1�r#�k�5a�	T���2��9�{>s-<G��оwc��9���_��Bx�!������]��(Nd��W�bP� ����,��S�/�+U}��]�_������80w�<ou;��g���hv���
�B&����1rs���=�S��	��k�ȱA?�nr�G�;��gE$s@B�>v�Ow/}��]���XpL�^1����Ƙ>8�q���_�=;ucO����~../�����)��]����}�G@�L�w�ǽs`<�0��q��xɹ��{rx�sӬ\��_|�*��?��Z׺ֵ���[G�t�k]�Z�~���W�ʭ�I�#fu4�W��@h97̆&�m�x��@��-pQ��zc��Wn��0����HTb�����-�����-�bE���\]�mo�pQ;�%[n?�lsъE�XPa�������� ��~O��Qu����lX%Gl�dey��ѵ�͸�Y�@|e+�0���J�Y&Ȗ[؍i[{�?��-��d8�_|)��k����F�q_�ݢu�\��D���La�z�H�j�6�N}�@H���rss-g����} `�����"T ����$�hF�
�� ����XH�V���"�z��;�w���XK/�X��F�lQU��h���r{0&�Ì���U�aO�uj67Z-K��X؟h��J�F��z]��������w�̪�pr���XM�u�0�Lm�DA+��IR� ��~`[����2������g�+ͯ����=��>Q �@dh�- �TC���� !��%�I^K%r?��)����؉P��|U�U�����lz|X0��Q�y}SW�J�@M���<�H��h�ކK�\�v��A���ƪ�Ö
B���x�U��;@FO ��ZA�7!д
�:���k�VL�F�G�򧔲�9[!O� �(l������~#F��fEE+w���5�V����{0���^6J�o��EU@QX>T��\>������Y�+���R�D�'���$W���u>�Q����M$nHtu?��ϫ�S���]�P�a܃@�e�#��+,��B)S_���;D	_0K��@,�3{AB a����$�Z���+���-�;�k��d1�y��Ej�V���|������:�h2�{rlJ%�9������Kۮ�VQ���JZ�ɝ\��T-|��`8.L����bv�~�j(n'�5c&~z�M���II
���
 . ��J#����kP�xp׫=�{?X|����f��w��}�z�1 �gрP�]�ݳ�2bU��t��,�jEN�R�T�g#�����&���@Ͽ����)��QR�Qq������Bo�E8�z���,s����?���uX`�R^�}ݽ}U�h����q�7Γ֋5��n����*���Z+-���J�\Fn�HK$dX�2�������z%c�y{N�z��?��h��ޮ��2�nf��"�tï��g�tk�c�c"�xqw��ޠ6VJ�����g'�cA%�x5�;��L�zC��,Myey����C6JAŕ�1��ߢP�|�;�� "	�������DU"�^�������k�����w������4lsM>�4�Ǌ�b�(���B#@���î�o�s��p)���_H�f�41r��Q_�~$�6:p��y���y�V..�x١��O��{�9��|C����ɩ|��g��ba��.����X&��Y<
	*��3������3T#86�\^>��>��x��/�����G?��u�k]��O�uH׺ֵ�u�Go��b�Z�ic0�V�$����W��p� `����QH$]-%p�A4�h�Y�\�=~"_|����|��s%�~uu)��/�������+9y~�a�}.J+.�����SV,���?��U��$��%جYM
`e4��j�z�w�@�DI�-���\��,������R.i�ⶏ,,.!��(�"苷�z�-t	���rq~.g痲��K������yn<܂z*=�}�X�j�d�5T+��  e�[��
���+����b�6�m��E<�8�X��ſ��J{�.�쭬��dI���a����X4f��Pű�d"�'�x'��v^��f�sQ�3+�7�~��6v�ʗM���Tp�d���!���� ����8R��<�ic�r��J}(p���K/����'Ѱ!( OJ��0���	0���)'�׋�+�i���	bV*Apd2�;W����V" ת�Czw�w=��9��:�ih>P>�Ҥ�� �W/�Y� Ȥ�:�]�屠���DX#�^L	�@�~+���L˷�GQUЫ����[[_���')jpɈ��By�H���vZ60���E+�ak�Ps��+�z�L��%^р/�C���Y=oM��5�����:� ��[���A���?��s��2���R��Ϯ����UV�D�vM�5�y�C���i��w�Bie����� �Ĭ�X���'J�xw!�nW�S�"�,�o"��2r�,� ������]���6��ᐖF�B[*����g��"��=�/r*�Zy�
kb�Y+T���?ғ���jeY(a��'���:���(���H��uP�P��*���������D�yJ���
�b�f��6"^��m�<B�m�b=��}���=,P!ʹ8�۾y%�'@���6� �~�(��Q�1����K9�`ˢ
����T����$5c����p���Tvm��c��7�D͹�ك�F4���x�u��J3p,�E�����D�3J*��~a�E��H��Hӻ���7��5�
��ޞ0��啬��QDru}+�I��_�9k˹���4����\.�^�����M�y�����i����S���H��J��!�]�{]Q3߬$��佒�*n.��Qo�m���f���3�����<�e2��ӓ3�#�d
�8���o��:������x�*y/�z8gqS/�˄*���+�o���Tb>�� :g	`#�B	fhU�PY�y֚��7w�n����@&nn:�L�׏��pO���n(�~�X���Ivb�����i�5���]�0�<��~�Q�B��atM'[��3�u��%mC/ݼ�$��ﮡ*����0�|�$aPl�L�鄪� yd��wO��؇n�<�7�-_}��\^�S�w�~a�u~y�,8k~|޸��ꋯdk��"%�������wʬ6��+�8;w�4%QR ����������M�6�./97������[^���?�6>��s�Z׺ֵ��t[G�t�k]�Z��U���ZPU�U����-�b����-���ﲺ2F�|���[��Z��-r>��3�������O�����淬bC�$���mw#���'�n��$�'�U��n������������Kk��[@��k21� T��}�v�� -� �*,�եX��{*V��
抂��q1pj�� e=�ʻ��}<&�~��C���ɩ<}�T�݂�����m�����c�-҇��*
8�p`Uj��Y ΄��A��
*?�rpp�P�\ݿSV��q���`*�#�JX1����.zJ�	��죁8������|���x�*���z��W�1�GZa���A��bᬙ����<1{$�v>���<�1�'���3_�1z$%P��:vϣhaXj����`�Zt�f�%��gػ�'ț{�:W�o?�*�0�Gurl�JYWM���a� �@php��u��D�)���H
���苊��Zń���q�wD1wx�{� ��a�{���eOի�����9��<!{�L��|	o����Rhp�X���wmi�"{���a�^kżuȺ	T (��{�
�o!�B��`0��u�/O�4'Kj-r̂琙����q-�C�=��×���S����<���:{��@�v�E�m�|�U�f��l�xn�FuS��0�}�IN�����_�,�6�n����}вR��y©��J��� �W���R��uL@��s@�M�$쑠�n@�������O�%Zq��=a2��x�ՎDf��-�ڟO~x��>*�Hzgf-���TIc�ľ�u��!*̆-Р�ʀ�����_��V�-�z�?	-�8%?�o�`����z��k�}T�����<y5GԐmuP�zOB�I� ��y�_��a�ǝ����9�Mr������}��f��xU��6W�B�C��$Q[�(���O@�hu~�s�q�M^�Y`5��l��TԜ��Bɕ
�=���%�� ���%z�3�,��y��/u�q��O�ª�N��RJ�Uj�����;4=�`t���j�N�^�g(
Fn�%@�+�n.�MLu���O����5�e�C��F��nI0lOwx�!���O��������%^Ѷ�|<�l�k���~�7W��ø�B�ݝ-�#p�R<30gyy�{��4�y\�1�
4��͉x-�3�閔����5�&��K%Ӫ�dF�l��l� /Xb1��\��Y6��T}%e�Fc�{���kD�+��>�e9��d��p��`�kѠ�e9_���I���b�6�{�Է�&$x�>q�>ޟrSP�)U�����}9�UVO�_]r�uzzbV��X�s��/�����+O��8UU�����.���)� �� zW�A��t,o���̮^��ũ\޸��ót"��؝�1��:�(I����_}!��P�o����?8�Y�{��g'�ʽg���<\��/�X��1�n��/�<ꐓ���=���?�Ǚ���Z׺ֵ��4[G�t�k]�Z�~�6�L�2X��C����᡾�+������3�6���e{w_v��RT!�E�f��ٳ����oe�<`E�[t�oo���p�),.�^`{+�D#02�<,���Ar,�ф`���5�r� G����q�VZ�̆��m�����g�`U�TTT̜0O�� `��/��ʶ��C�jH0$�X���VJ���ş�����_���+��'��������S������>�$�Q�cG�j�L3*h�k,��\���	�������yyqAB J�B1z�T&O���6=�?�N�[H�r�$H@���L�rŌTn։[|�|��_h$�~�n!?R�r�@qS�,����j��z|�R���5��j?,�aD�Q��O%���Q���)AFB��k����)*ڟ��˪�TP�`f�����]���Xb[�AB����`H�JI4|gE�؝������X+��k������-��%4�o q�3\L��h!A��|��Zՠe��{����>��)]�xh�]5n
ouS��}�A{��f�U[O�/(���`��h�|uz�
��	�f%{˾�䋅���8L4 �gn���~�R+P�oVD$����N%<I_Yn��o�*Rp]�a��U� Eevm�m���Y	�b�>�m���"�>v}{�/���:S������/{o�$Iv^�}��ǖ{����0�ˀ�"j�$�Iz�ЏӃdz��ۘd&�I���P�XtמY�����9�w="��ol����232��������s�]�*���%�' ��MR�U�1�'�X_�8)�PB�옝/�m��k��wx6~Z#D�H�A�D�F�0H����J�}+*!��s�.����URE��A�>�c���Ѫ���{࿋���������a�r\����!f{ed2#uz���c�����V�=S#�c
&����Ϸ���n�u�c������[0�J��{�22���� �y�H���:Zw����PE�'E"�q�p����&�p�E���J`�L��,����"��Hn7VqF�~�*S`��Z���E�מ��I>o�u��`O�Ye�sIgy`f�eb�H���:�3������cj��q��B�MK�Ǟ<x(�`&��=�d�:�������xE�W����Zn�يF�G$!�.(�`��\<�����˗\o�>-h]0�W���|����M$�9�#�Q��%z���b�<��$��숹��ǣXf���\mT�'Ȃ�L��t�5r$�j�L��فb8�MHj��(��&�5i��>�@!L�$?���e��n��V���@v���F�
Ul����$���ё��vXT�B�)2W,��f��Y����C�y6v��Q"�g���OhQzws�b!�@h|������%�o�=
-Ɓm�"ds����8PP���ǹY��՚����L�,�P�5�P8�	��4�&d�IhV[MEܬ��*�Hg����[�^���XX,�e��;d�\>��+�μGъ�3�#�,޿����_S�S���}=�ڭ�P0eR��kz��)�?������f�e���w�ܹ�wX��ʟ��_�O~�G2��mhC�n�� �І6��}�ړ�Grs���i���xr:��������Ϯ�6f����t�ɣ�S�����ۛ�*ݦ�
�5��-%����_|A�#X/!$VJ�T/n\i� ���eA�����H���x�i�bo�M���#y��\<z�M��mP�eś7�	��ۂ@*|�d\�B��8�	����AU!!�M�&��h�6�g2
ݱ}?�������}%����o�o~�K�V�G>��]� M_�m+�~o�Q�"�V�T����F�1l���:�q�Z�I@2$����U�V���-~Ep��#MK"$O6��;l�̱�A��Zd3�a��Z���*��  ����D�����_ DP�[
����65)�f�P���	G�%�q�r� Vm���2U���U�$�y���*}�?�N:Jd<�H�ς�W���zʷ�����Q�{��~ł��1���߅�U�j��@�K�V-ϊmd����R�ޕ�ү<m�Z��/��jc��ДP�fu�Wɚ+��=<�	R�Uٱ��38�.U��j~�}�i�a`6D}f,=��A��C �@�@0];�?��<`��,�B��a�G�'8|�?���0�Z���������>�G+����(�-ǣ�w��o��Z�Nk >7��8c�����
��>$@��]���J��$>P�W���d_���&���{�Te_�M;��{T5$ ���?�A�<�%>��
����S�p�0���Q9թU�� q�Y�=m�b��x������Ty��	�� ƴ�|��o��ji%F��:���l:c��P�+Cݽ+D���<��*�0����<���e쯉�k�5�-�W�uJh�5j� n*#L���p}b�����������b�W�\�u?���Zp��l�]�����1ud`�3lQ:�fEh�'+joG牕��-��`P:�Fd�h�����/I!XNz�ו�p!��<��
���~f�R���M��ʅ��;"��ё���P����f���ݡ���U+�6z�y��*��dZ�>��G�ʏ�פJj���r������5��O$9�Mi�4��
�n���Z�8�׋[����
@��\RM�Ǌ5Pr�.��bê���J�f&(]"Y��r�w�Md�Q- E
��w�*h��\OF�~�V�C�=�^X쐡��Q���H���\F"J�N��
7&6��G�C ��2��G�e�Vgfq��qE�������L8�0Pݭ3*Q��0j(~���%G� ��Lp|�1�~<I�ɓf�A�L�m���8��7�ߐ��Z-IL���ѱ�@��{2�@x��1gf��d]���C��"(~�~q#~<���F���uF�u^�@��Ϟ�o~����X����9�­�OΎd����^A���S��<ws@%�߽��ݽ /��l<"QRVc�󱜟�ɧ�~�~����~��g�'2q����AY���O���JJw=��T�6��mh��6 C�І6�oE;�f��i��s�i�e�#�!D1��t���w�C��љ�?�DN�N%���4�V�c�@����}�F�۵�"�n3z�6���e�DC�AV�y�N��>�l�q�I�v�bǿ�3��m֡n����m� ��a�6\'���;���'g��xD��b�&��m݆���a�+��WqN� ���|6�����m�w�Ƶl����l	 P �����_�~~!S׏����?ȯ~�� \w͎�|��1���hi2&�@�J�����$ �x���w��q�VC���kF$2аQ.Y�W��<��*Q�]�Z��L&Zd�=�Ya���2E�Nt�"�Ւ#��}x{����UX��яlE�Y�� |U�,hVz�z���i,�Oؿ !�� fk��]��Sh�I�@�!�T|�ނj)��Y	��Y���^K�����4�V`{��P#�V���A̪j�q�?�|n{�4��B ~���t�Z��� C�W���S��
���K��>̾�}�����B)�L�&�Ֆ� �\k���?<��A�A[V��S��h^ʡ�O�u��B����UA��3��y� j�o�6S�L�8�k��4DǖD|�WH�����  �}�E�=�Y�Jh�@�iN�z����O�A`O�2>g��������S��C۫6Xv]{��f�wv��S䱪Y��a��]� ��֜�r|�J���������j((1j:A�O#���
�iƓi�sl,��?'���3�h�6Jٗ�2��{�V�Ȉ�O(_����U���>XPb�wl��9E�,����������อ�!�>;�",�-F=Y	PR�F0˵}��S�~\��&��wH�����}�k�$3L쾍"�U�-���P몰���$��-�׫�ZU�����PeN�?]g_��5�Z���Zr鿎lS�S}�����qc���/�h�c��Ic9=�?ք���)�
�3����v�;�C����"O,Z(AKC�Cܺ'ϛ=�`��C����Ŕ��! �AU>T�����$@��~���E�暤�C}FW�̂�Ӈ׺^@6�FG�<��֭wVɛ�'c�F�X?bg
Fz�.�D���:����c�=�����������H�n�A�K7��n݂+���k�����*���D�g�sM��ո�qϑ���1�l.�ǘ�'��z۫�@F:�s(P�*��. A���tF�	�)r8��*ܱ��<6��ٮ'��Ծj�~ggg2������s��L���DT�rr�
�wnm�� �>�\/{Gj�<���
��ij6��v�s�[\����T�\U-��~��J.'I�u:�8���*����"����l>��Z�/I��]��?��W��������@�}���\߸�s��J Uh�I�ַq���׭�]#�ĝ��Խ���>c�މ[�#�6iӒ�6��mh��6 C�І6�oE�5�T�k���Ǐ.$�r]1_B�j�p�N��|��ǟJ2�i�� B ����bG 0����j�$�����'gR�����_�95E}�l�2VZ�G�^e�߰���jh�5,�Pu���s��+t@�\/$A y6&�2�����G;����Օ��7_�z���;V�aS
b%�G�������%JV�E-��X�����?��ќy s`W�O�{�m���J�	��vJlT���8��	������➶ui��(�H8����R䬔�R�����b��m�3�Q-w����� xX����u6�a��T��\ߏ�k��@ �Z����h6f��zc�[�s�®�R:�h�� ��r�}��SZg���J����X�N�l�3�Y��UFׄT�D�W�,4|"4�l	�ȣgw���o,�HJ~�$#�
�e+ T�P���Ų=z�Ȫ�*A���Q(SrS�;
�>Q�� �8 e�|� Ta����� j��ת��: �b����TTU7fs��=��� S�z�ڿW+H�*Yo��JU�^9�<� �ЀO�C� ���hE� ��gY �^P^����1�i�c�N	��n��q�	��F�,�F����ܼ-X]�	�8�[�!@���%�_i��C ��)(z兟C��f��ɦ>C�Ȍ�W����V��S�@!���>4��ɏ���33���s���<i� h� k�?���U!A-�/HsT�G�ZP�q|U�����y�����Ǔ�c��DLr��PT�H�v�v#w����ȳN�@T���H&�dr�Fc�$��9��=D��"qY`�,T �z�[����{g�|FW?~l��oXj�c�!���Pmy���H��߃TH�q�@���EI�ГפK��"X��
�s�FeEؘV;�ƍ�ٓ`��e����Czߑ"�_�ĿӦ�����t��U��'��%f9��*M�� ��c%;�mc�"�F4pk
X����q.�� �uZGB��6�T��XFN�$�'?��Ь�ڇ����{7�j
72���m��[S��"� x���p�absj�P�^z�H�3���P���݇t����"$*�^����,��X�j��j�����?׹�q�w��"�������F{%�*U���t6X�Aa�5�����6eT���
(L7[��xFBm��0���5�f���x<�Z�C®h,GI��/(b��%K%Hkw�3D=�o:��u� �q��Pu�	��$�S伕eh���k[K~��+�*�3�>��1�9�����\���ɒTU�6_�՛���������<�5�[����d2�Q���)���Um�l�C�9'�q���Э)�d�:����]x=��|�e�&�`ն��ь�d�Ѯ�ސ �Zk�4Ve1��FY#/�������?��B����t���ƭ���>���!�@�����{�/8N����|	'S���t�֠SY,��W���	��&�&� L*dhC�о�m @�6��mhߊV��z r���S9��	R,��$������;�u����X.�/$p��z�An?���m���')�������m�&2�v��@�:T�n�vn�'q�*2l���{V�����"	��@�����}66����Y8��
�P���w[X,8	;�,���Ru���ѩ�,p���L��3��P�ܱ�ݮe���v$��{}\ў
�plP�RC�;V��T� �א�N�ƃH*���������tgu���^�bŝ��ս�U��]�ʘ�ɱ$�s���,�P~`�����p4�(��iP�l<���V�>ܸsY�.�
��L��;����r�h���]_ 6�cL�~̍,*I�*� ��h_���
�L��m�cݠ�"���/O�<�o�f&רh��u��X�6xS5��ݘ;;>%��*�RI0G�OӚ�L��%��䢤%K"	7���&�.%�	`<F��YO(HP��gn��\�]��ҁ�B"BY��4`�̎ I[���YZXw���>*;Q	�Y(j��<�OW����zG�L�u@�H`9.b�3ql�jPD�h����h�Ш�ۓ�]3�(	�q(ZU������W��]�a�<i-��	�=�Y��8g���[����T�*���B�늄I�/`�c6G D	d����V�֕�p\�͒���"	�'����'��C0zu*\Ӏ��XtH-5�ȧ�R�]��W�C��W�k <�Q�Y����ǁ�렫�~��]�pS��Es?��X-������o
!Uf�$��ZIV�f:Ulu�
�$�*+�:o��R/V��Y�Ŵ&ȃ*mz�&� ���l�R�- y�jFLo!�o�{@@Y�{ؑ@�ϟfSŹ�j���*{���;SbF�.B�F�xR�@7Ƃ�}� �R?csX�9�I{P2����滍Tf-�V30:�i� /ν7��J������{�pAOG���&ƿY�ߵ���0�"���3"fs�=I�`��KvI��Mg���j#���.wj�c@82�R��W��6�IdZFOCR*"(��ukǧ��ц�'𚄯������;֢ɬ����r=qc$_��JI]����JTI���=vP�Fȳ�8'X'���L+%7��X����������T|z��A���
���Q�E;x�*��d�П���ȫ��'�[���g`} �@�)[�7T�*A�������9�1v17�0�8���'?�>$�ir%-����f�����rվWO���/]�6<�h��z�އ��^���s?��j�0��_�]'�W2���u#���P	`���|�sz��ڭ�ܵ�$!g�S^�ի5�MP>���q>pqq)g�gr��1yQr���P@�XQ�<轍!��v�{_�����NR�-sc&q��4�3�=��̊�0�������Wn������-Ty�m��$��O���\���n���ٳT�`�bʹ�_� �~�M��+w������yGs�Op�!����ycL�H�+B��)A<`|�g�ED�B����ۻ�D��j)��ĭq'|�H�������d1���U��m��d���p��t2b�ϓ���G?�}y��s�����u�j>��O�qm��J���I��
Bt��s�]�<�H2�p��i�.tϓ(��H�6��mh��6 C�І6���P[��Q�6g��_��ڣ�n�y~�՛V!�Uy��7o�H���U"��կd�p��:��m��i������m�*��=a����盝� �`��6P ߿ˌ�9@��
���
D]�n�qÊ<��t�+�6I��~�
�@[o�
��&��vn#��H�~g쾇Ppl��YKݿ���ob��fÃ��vnc����Zbc{�����;ywu-����■cK��U� oj͍@��Ik9# �ǳ~S�tܵ��Lkb�J��U�ذ�f�2gAQ�{ww�*]V�͍�KG�{���FBS���PQB�'#������\�n�P����B���,�H.x	[V���i#Q�E�����%���l��վ���h�2��1��(�e�!+P�����7�'R�QP}�E5�# � ��ULS	�e>��U�HA�ZXM�vq����d�C�y��38���l�d'Y����h��Me�����m:��Bu��3�a�tZ٬v5-I�C�)��fg�Y(uh
Sx �yf@�߶}N�"��-0	�*f��B�A^�����{=��ث|����ay#���������
����U��T�6�V�4@_��P����z_�s�) �(F���b�9n|7EG���4��u1�8���y�}�U ����_�����k�Z�[���w���9����n�\Zr��v���gx�)e0vHSZ��W�f��z�"����z[/�X�l�1]����x`=ԅ{"٬�Б^!¾rc�� ���[�Q��W۪�1=�����r���)4��a۞��k�{�z�2��V�: f���ENj�GqCk���I£�I�6Vk��=A�=޶{k5���*�{"t��ڮu����%�E�;�֓a���g�fO ��E�=s�#O[�Fh��x��MyŘZ��J�:��x-Ǆ֋���њ��~Tk
_HPh���T���q�<5�@��O�����a��$�3s������\h�sۇ�+��Ͱd�u0:��G�W��4V�
Ȳ�u�0�y+	�
�&}�C�R*R�^	� �������Wc�$I��T�H�S���@vE��&�;��d#�?H��MU�;��{����Fυǩ?�:bl$u�vX��	�����#a����ױ�<9=�Z$�f��Ѳ+�2_�^�J�'�S�^��̓�(E��fb�f��K;ڊv�D}�豻�(@P+8^��Ԛ1ƳͭӺ&!9�Ȝ�V�}����׿V��㧺�L�y�� Y'X�BA̐od�m�T��|˷[��j��,��(<�B�ɂj���rz�d�z����*Y@�y{�"�y��h�3̫�f%!�h���p����,�ykL�]�*g%��n�v��a���:��m� ȭ�W9符zF9�D��#(�y�����9GׄUp��*X/Wq^��h<w��n/��І6��}��@�mhC����[uw�6���`�L���Gf�j��[�!'�К�����R~���ȟ������Z��{��z+�IB�c�~�$0�`N�
8 n�ٶr�6U	�����T�,�\�\\�A�
7��2*��|�Ъ/'�L&��H{�]��x��j��1+0;��û��UKp��ș�f���]�
V�}ll�)�N���Ű�@U�$�;���wT�l�+*�\��P 0��A ��QE�N�`1���|'K�1��3�|��]1�̇�zp�U׏#������� 7�*�m�q����;?;憛^� uFޱ/aU����j@'���Vm8~������]OXV���O><|4�����ص�y�o"���;7Qɼ����a ��Y��U� ��7�;����.���>� 
c��p|�Y���3��Bȑc@�$��K ZJ. �����דP����U�4�V�k{=P<�٦��E!voD�~�ѭ�oL�8d{C� �+���k�k8fH?ZM���;����#����UPr�О�@uTٲZV���J�*�f~�}�3�:2�%oM�ǥ�� �������hڄ���<��bŽ������&�дQ+.̀р� ���=�`�k'�����
4�[��Z�;��ZPj`�X���4�Ϋ�g�z�Z�(�k���孄<_ae�@c�I��JH���]�_#H�h��:���@g7P(����0�2�fj�	�s�p��'�č�H�l�7앪�|�,���¾>�9Ƚ�9v��D�^A���3�QfD|�:�C�v���?��h+�}Fb�`��|Or�
�{���P���Z�Q9a�`k�M��h�8~+���g|�^�=Y�ʊV��[eb�p����5,<Ž����'jy��H�p>Pp�����WdV��&��̾�j�]�s�2��Z�A�{��Qrѓ"PTU׏=�V��F�-�m�[�x�a�k[���j-�F���0��
�B�T�W}6�((ݙ����*0e��'8�V�2dV�Y����?�m��m�).�:�}!I���a�O
��?���G6FCuP�I����S��怂L���m�:�0��/�ݨ<<e���ٷ��o����_��n��ǋ_l�r�@����=�#��=;�<�ˋ�j_���@|ޠ ���+�<�ũ����%U��;.<�޿y��ܽv+�i��!#U���5���h��[]m9����lDX�Q�mi��U3�{t;�K7n8N%��TX}Lz��|:�h	喑nn��͛�\��z"��M��5����s<����W�;�Y��������
9�X�`M�j��	�Ȅ
��O�S�	;��Z����l��
�p��q>��E�Icπ����"�j��"�:1B͝��E?T�f��֍��
U������^�u��w�=9:⚃����`A��u��U�HrkY��������+���~�v��ݻ��v}<=���������/�ۗ2��mhC�ε� �І6��}+ڪ���̓LnKY�9-G�.���y�683�3m6����ȯ��\���U�����̌ ��f�6�+fC\�]�ncɠ�P��Y��cK�_I�M�M6�S��T�X�!N���A�� �{�0,�%ݽ6/"n�a��\������S�A����:d�A��N�ܑ���>8���Y��VYw{{kVGf��%��kQ%�Z|�4u�?�U$�͚�8��fK?o���(cu��Zk���o���Zx�Z�n@`���,��O��9>�m,^"V���q^P��s��5�ڨ:^�̫Ъȭy�+��ktC�
uЁ�6ʨ���J9;;e{�h�YU2rY�H����V%b��
���9�q�>���l�@�Cm�s�4� 8<��j����<��OT1�s��Z��7����~��µC���6f�"�8	c�W�N��+
�z`��W�f��}�GG=�A��z�߫@�����m�X��b���7Q��0f:�*�+�|�s�atp}���S
B�$1�����{��H�-�@�}�8 ޶��h�;��8���a���>0�,����.�>���P�3��������>�,�Z��8m�)�*��J�����Zb�����G����}fz�\X���o��| V��b� ��vp��hڢw=���g�P�т��+��$�������}�����|A�Ԧ�	M5���s��y8F���Q��-*�m|���P��_�ߓ(��䞄�J�Ⱦ�J)��~��8��gp�c�����q�m}X�^7���y��R��#��I���)<�����?v*g"� ��F��`��]I Tj^g~K@��3���X� �wǱss`�̆� ���72� �����J�^����i��yEB�Vf��xU r����Ʃo������YF%c��K'Q<�gJ�D�X����!>�\��>ol>S5˞�9���$��G1�p��ފ44�E�1(���
e+<���ϑ�u˿}�Xա�k� �֣��П��e�y�.{���F�����������	�=yb���#���L�uW2ٸ�����nM�����=��#��$:�WնP�P$���{����\+͎�ʢ�F��)���$`{����j�uF{"����&#+]G0�E|΃��&��$�:����lCq��I&�^�,4��׵\�_��,�e$�F�����v���*���#�:������$�,-���1�IT��"Pc<��	�77�r{+��,���,�$/x��L)�|
�~	P�ïbS{L�u����]Q"'��}��uX]�T|�Z��z����vӱ\Z����|����g�Iu0�;U�1 �d/_������_���Q�'g���߿\߯�G��\�6��mh��6 C�І6���~�&���P���D�e���0��mܗ�|�Ꝝ�]��蘞��L^|�ۘ����$t��H����*Z��~>�Y�~��bӗ4/˂���x;�5�W�Ry1r��� DwZe�`l��(��x�g=�3��	7�Q�J�5�N[m�<F`i�_��w��i8�۰S��|�嗀�1�BIY����X�X�J�q�h���U���L�N���b�����������ɉ{�1-�Vn�e1}�y�
n:�� W�R����X��Pmj`�E6�gf�g�Y�n�Jcxcc# �W�þ�Q2 ���� ��A����͠~�@(Yiiu���k�0>��
|T4�G�d���<�nsڝ�Vn�-=���岫�2�B�qN#*=��Ε6DZa���J+A@'f��h4�U���Z'����*F1.��m66h KhE���2��{�S�).����?����,��+����
�JeTH� �I�����Ҫd�_fY�m�<�Mp.�(������֣_�hn�71`R��"����a����8��
��ω��i�=BEC��#fy���#B����вX����+��@J+؂��"�3��H�{�`AY����IF)�	����L����W#��ԓ�X����1�
(�%�|ys@Ą��jUP0�=Ґgk��
�nm���G
�=`k
|zMݽr�����X�2D��Ҳ4����j�w�u��[}�t��B�}�*^R�Y1�5C0Ec�(9!>]�����GsT}lf�<$ؠ���,վ����l��Zj��Cv�+H,�@�P����c����G���0l9�RSS��(�UK;UR���B |H
��I�<������,�0g��HZ>ۚ	G����1���Vm�B�f�R�	��n�^���`^ɥ��'���x���,��|�H�dr`O�Y����Vo�$+�zb�7Ağ�$�EP�9��5BgD"��l�"����(�T��UL�%T������\{��{ �lN�*���~
���v����Z�y#�*����$��v@,��(�����1��fNZ<E�Y#?ǫ��?���$oĎWIUͥz/VKN��r�E�\�� \�[U��^Ȳ3�Fi̵�>�����O爒�e�,f���,B�WYV�F�}�΢	��ļ�\.�=P�uG��K���-dƜ��Ad@c�	��ݰ�;>���
j�_��/��ꎅ*P� �$���P���XX�ǅ%	�JP�`>�yEC��[a�s���L./��:[��q����9W�	�@q��w��b?nm�m��ƴӐ�V	�(�T��Հ��4,�[�FQ��G�����Z-$ߖrs�^���Wn�s}�/��\X��q�&��G���~���{�۳�n-D��[w�Ž�ş����~&�����tܝ�N���q<�?�~x�J�6��mh��6 C�І6�oe�F��}�9>?�/��R�=����e#�Oݦ5��z��m�	�M�޼�W/߸�*�*����;�,�h���.�H�6��?v��=7�Njk�j��EL�Qh�*6˭��b�wtt"���F�9�r���|��� l����nJ��o���^�j7�y#^�Og�'��춴j_� �ѰJ����l6�F�6��\��"�|[3����S���b���7$@&�2�
�A�0��[�U�j�bk`Bː�҂�A͏�@
����_3��*�`v��4G���	x�} 0��N���ss�$�$�b@�歔��z<��s+�r�X+��
�5���Szd�4��A�w?wc!�t�!��W9 �D,�82  k%W�jiX����<ڏo���i X���b�Fz��-�j/R���D��A���n�C�"n[�5���F*@�S�L�,�A����}���y$#9�����[g�������� %�?wA���{�+.�HS�� uAq�F]��R�kի�>��Vu�Aѫ>>j�@�kUs�
%�4�f��'xj(�0ođ���e��֒�>'>P8D̊�z�j
S���������y�ͬ�BCM����Qa��.��F�Ԧ��>�TǓYHu�o���3�"$��V"�]bO�v{ŉ�W�U�����U�{�`Sf���ȇ �ɬ�@Q@ �#6�y�D"qAt��� b�/�f����g�_���,�9N��k��~�/����{:N#�������0�ya�k�^�c�9l��0�y l���5��]t~���}�����J�q�i�8�DA� =�&2�@T)�|a�� 0R�S�w��^���k�g�Zky��~�c��<�i�Fmd�'EI��
��e}���8dLi����~׫����,诗'U"#Ga���c��$
q�m�۠�y1�*�@���!�k�~7[�o8נ��Z�D"U�����ʼP2��l��8LSb�|Y�ߧ�z�j���^.F����̛�:�.XT�(���^Y�m�o���<��Tz���.�y!��;���:��4�|��&��ɹ��b�Am6�l��G\W=~�X��|��K����<��y4ՒP�l-X8���.`��~�7�(��"4�0>J��F2v��5[�2tb{��n���b	�N��WGS7~_����r�~-�M.����P�|���`��٪�[�M�/	n�_��f~<��W�iv�$�2��ɓ'���S��NH b�{w{ǿW+���J1�P����4�O�m"#@p��~A��H�ѯ����T��g�ԭ��P-on�v�-��&ӹ,����Bp:�F�
�
���Ǆ�̫a�B�������?�o~�ܹk{vz��g�{���=o�ե[/����������І6��}��@�mhC�о5�1�5P��} 6�c�����ɏ~�#�����#V?v�9���a�jop��=*�Y��r%���o��7����[)�Q�Z��XGTn�s�{����dEg�����R����<����@vG�d�i�*�Y���n�4�cDદDTȪ�!H�	zY?6� ��ӌ��(*�v�{$6�#	���<���@5�����R}�T9I"����}�\� Y�V$64;�2� N$���h*�	6�װd��1"4��F}��N�i�-��&0�2"ؔ!~���O�? �
�U��?b�L�?���0��T	��@���5#%���)ʭV�G��9�g � m'f9Ԩ'�����ig�4jl	>�f��6��$1�?��]\נ2+���P�S�{���MCF��PP`���T�%ib�;F}�0wo�U�4T�>�1��ZXDO� �wτ{��΢�@��pˊ������T����,�:Vy{;$�e~�[�Uo����#���
��"4r@��> :z5���>x;�lMcV9��䍌l��A#���V������m�Bw@zxK����
^S��1� sT'�>���3�Y��40�_v	5�;�3B ��s P�*j,ס�g:�%�6W�����f����9�!V�¿%��_ PWп��{����}n��h٫�h�*<a����<y՘B�n�@������A�o�eR{��$�tb�~���ωN�׻#)�hӫ�� �N�����9��ɤ���N�	kѹ[��8���m�hM���^�������`�筦T�A�����	T�]�*-��_�q��~�+��]ꅧ�b�^��Z��JF��~�b�϶0ҍc��L�mݞ���Blįe�H�ߋ���Tv�q]oA�ǉ����F�x�%����oS�Q���Pzp^�sA�I�m����掾Ua�"=������^p����j�8���*!�W�6Z��35�n���@+�ܪ�,�֐�i��A?�m-:dK<�����·Ǧ�����C��1�$~9���#"���><ƨ���#��(z@��>G5��°ѧ�K����_RQQ�]O����H��R�>{"c�>�c[]RA�1S� P9�w��G�y�����A�-0M}T�=�|�N��~�4�gQ��Ͳ�ȫ��TK�m����ӓ3�z)n�����r�v�\p͘M'$j`Ǫ���nMI�ʭ�T�yrrD��Ǐ�z�����ˍܸ��d�IT��$>�����8�������X���H�5jIr&�j��B]���V�(B���&S�־sǬ�n��}��k�G�ۋ��������_��E�Y�����W)���L~�˟K�\?�H��'�g�{�#7^��8����Ї6���;�dhC�І�ް�b���7���ߗ��O�T���+�؈��mlQ�� �|�6N�2�&*�8�:���A	���+��|$�n���H���a�*m�vt$�*����q+i���� i<𯕐,6ce 6ϻ<�f�y #��d�q�
e|M�j	�h��>����e$�ŝ;����VA�݇MY���#m�5~O�d�X��t�J�$��@X=��� 7�mgUݚY+p	
�LPI7�^�D���>��m��(���\�W��U�f�t� ��)VL�j��M1��Q5��[Zfn��{��x� +��J���魢Я�J�"O%����nCO�t��s�I ,�q�TH��Ǐ����ȢV���P���&���`NH> �<�5F���c?@p�w��	J�$�@� �qc/,i��5 ߠ�E�U��'-UC��n��q}�fu�4�x���}�?�+d� ���{��������v��fɪ1�� Uཱྀ�S;��W�5-�M��o(��t
��^I�}D
��`���~j��"�mP��-r�<l|�����(��
%�'�м�	�ˏ�Gj;ը% �H��([!{���u�Tx2�zl���
 z a�VTu�=	��B��(d�����9�U���IU�y�$:Ԩ	s7T]�vk(�]M �>�+q����J�B���u��<U 5�?��D[5~��c`�J�4d_��1ΐń1����Lr�J�ؐ��#o�$.�+	L]��3Op�X�Zhv��s!l������[�j�f�hn���6>}���>��뉶��k0k p�a�I�W�k�S�_�(�1�CX�luS���4ڿ �I
�{F���݀\?���Q��0��d���C���|1��iL#&�ku�Dd�d�Y�͇cS�g���JS�����y<���ùh���=���T�R����N��/`� ��+U+���5�j�J��5c�V� �H��VmDA�{A-��W��Q����?_�������a�D'����s�Bǀ�-2%��O��ofs[���d6��"Kg�'fH�Տә�7k��vY�*R�1/,�n��~h��s?"KSo�!j�eq {V������T-�[?�7W�;�c�y�v��[K-h'��|����0|��gR�;*E8�;��T�!�V\�ic�B;e�c��OXK4�{�a��4OC�A��ۺ�!�\P�$��sk%Jniw� :#�p���,f��L��1;v?[Pq{zz��u}M��Y0�8+w5t~W�@��-��G��s�H@��=vk,�c >���Gf��Cu3�Y8%�����:<��"H�؞�F�`��}i����yf8�[�v���,7�GX��ǚ�����'��9���������S��{�c1�d<��e���o����o���o~����������\��L���M�|��.�.�>O� 0��mhC��ar�І6��}+c Z�2�̉��K���3��?��r�6d��0盜�ͮU�"L�%CkU��@-�����'���A��7���L��t��J�PI��4^{uu-��� KX�M��ٙV���X
����������ۜ�|��dU;<�Q]���p�6_www��]\\�(�d�˹��c���i Bp������!��AF`Cy�c6�!�P��nCxvr"#l���##X��>��/_�gؐ�w%���n\[�������Ν�Zn��e�^�X���>;u�+(��V��U��u}���� �V�*H�%!ȣ��;6�~�f��Q��'��n��8'�����/�ܨ+B0��	�*��#ɒ�V�VG}��\?��xH�U�{�����q��Է��_�r�r�&#/h�c�;���ٻ݆�{~�Hʢ�w��KՕ| �mS��R�,j�F+�������ɈU� "6���-����V��*��@vsO�H����:bP�T2��1�$��a���&)��K�F-]��(�U��$Z�,��U&1��qSE%	�	�VA$�P6)h��蛶݇�� =��h��`N�d4�k���:�Џ_�/�:��f� �7U�$��תn�}��Z3�]����(Љ�y	µW{��,��NX=	ك�8'X���F$��R̦�ד�B�}�@�V�Ǭ���X���66k3����{Y�}�JHr."p[�Y/�����o,��daf�/( �V���s�*���V�f�z-rw�;�^)��h]��g�� r[*$x$��C$��[��Z�u;�Oo�Q]�z.�	j $)܊�+w9X|*�1^TU��ܵ��k:����+P�@ӊ
�]�(�����,Hz�P�վ&����ɮ���
S�D4�Q�PPW���l,�|�5��20��<�9D8$�?�9d�N>�ۏG���{f!3���PbQ��z	��p�?c(%@D�9H˘N�]T�@RTJo��p�Wչ>ߠ&�4l5�YL]���.�J��m�m���*k�w��4����ۖ��e�8.�;��� �%]�c�	�Ø1F����~>��"!���'�����uk�X�A$�j�J����L ��g����#6��]�J�l4�X(˜�_\�q��ë1W�^�3�M;%�q�k*a�2�ܘ���V]j%�ǽ��ق|�+����s�`n܇���S�Iᙕ�y������7oq��� 00�c�=%<"���f�M��<s8���+wO�����h���=���f#�YQ�g�;Ǥ�|^�E���t�����'c�F�5��P�L���B^�_�������grq�����Ѓ����/>���ky���	o騑�n�X�u������u��I�$ٗG�`���֤���T	C�rvz&'����{]���FXG�\��QĹ���X��&���u~J��e�}�h��,�<!H`��]��h����ֻ�}��[۞�`Yix!�c�k-��s�mw�ށ)̴x��6�gF��AA�"�Z��Lb-n�g^/Z��{�.�|e㵓7o���~!����\m��k�B&�y��3�|�D�}�\~����<{�	����ݱ������������%�������/u~v�0�Me�ֽx>��3h���rK�$
�.���w}�6��mh��o2��mhC��4X`����<}�L��?ӣ�0�	��\��F�v6v��\T�4	�����k����X��K��_���^�H�[�Jӌ`,$a�0%V�ښ�R�M�T������`T���m�ohÅMh��/"�>�{�� ��T<[h������F�%Z�߃Z���x#�ߟ]��V���W�
�V��\��;��Ƽ�W�F^�z�՟�|JGnӾ��{m��L�6�$����I��U� u�����f��%t,עR�$_هV��q ���ñ�m-�d��X�T� ��T�()�k����:`�������'�j��۷o�☺�����;�G���a���`d���ѱ���±��q����|v$+Y���p���q�K)Y�Jv�˲�� ��R�d��u����;P�����7Z�J`�ɤ{@���*`4�hl��M}�M��o��nUa������֝VςAMk~$P$��-�-�-��5�X�ɱU	�\���C�s���U�>����0�/9�*��&�b6�&j5R1P)"�Ѱ��1˞ڀ7�k������qڨ�m�����DDF؀P��ʞ�d��ok��L#` P��f��݂��_�  ��IDATނ����/#�%�*�#�bH�M���L+���'�\�8�	ڷ�z�̊���Ğ��FX��5	c�-u�Rr$��҂���g�=���V��3k����D�I�������b����N��P�pX̖M�U������ �^cxM�����Q)��/io�_F�D��#U�J��PuX��9�sBw��A@���MOlF�/��q�n���� ��XMg�WWM��'��d�}n��wu��H�@h�q���4���ڠ���%������s�TB��z�^T����-q����঎�J4���z�na���TȞ��i���a�!�mD3l|���d�4��_�D� ���@��b✐��S��.��C^@����3��H��T@�G�P��*�q�8.� ���+�8�s!���'�,�g`@��6�cD����{ ��z�Fs����d��Jɀ?�l�ԟ�c�e�IM�'Z	ό�p���D+-��*U�u|=PKB��	f�VA$�Pu?����30�`.1GB�&�ͣ8�d�	�횿b�.KnL�G��BX7 ow�PÍ��6�zi���13���q��#�
he���h�u��rdzDn�c��Ɓ�x��f}� �^�ӑ�/�}�s�1����{�(�� ��a�y��b[�b���l,�=�Z�����<~D���F���@?bn�� "W�T�U�y��,ZI�x�ܘ-@~@c9P�}�O�����w�me�X03���c#���u��������
��1#�V�;r��|����%O�i]
%�J��N���'�G����Z��\wiO��͍3��9��1��Ę6+Q*Xb%�L�
Q(�,�֯Rkn�L���}	�(��]��-��0�k�^���G��������9��'����B��;��zA����S���~!o�]�d��(�B*����}��&O?��'h�� �І6��`��mhCڷ��69�)�p�;l�D����_��?����nӾ��O>�F<geǍ&6��3?����L����M�ۄ]����������{��fG�`͑{`/l� �P�h����7�
jb���8 G�(F�Ý۰޸M'l�E�/<��|�S�KJݒ�&����1�� Vw�jʰc�)l&��G����2��Dx�9#���Նm-S��G5T.�޽��r�p�6�|�p��B6��;ߤI���'��_s������_]���(���z}2nv�W7� ����r�2H��+���)8H_��2iM����d��B�d���w���3=v��Kn�Al��ά��* K��N���d�q��]�bg���ߧ�Q˯�N&S9��ן��~7ni1�XN�;2"B�6�{׊D�me�*���Yɉm��=��*�a��/�$��2A����߯	�ȇi��C=��%j4; T �2�ǮI�ڀ?��{�č���Z~fàt :�=	,  �-� �)Q�^iF��@�� b�<����[6���& ���ƈXE�W;w=1(`�՚�b���c�$�3YBpC%b�� G���N�޻_m9����͑	x��0���?F�t6~i�ZCÔ�.
-
4CD �V�����DT�'ZML�&��Q�W��`���JP�X:�fy_���e��O��O �8�:�p��SQ 6 �I͒IҘ�0��Od����J(H�ڮ�H�!W��Tmg�$�'�� j35��*�1{�Z���*�f.��4x�)��|�H
�y�k� V	>��e�4��8G\��m,?% ��3�������=�L'c�E �x�u�/�����z: g`'e^�ח�����x~��
�R��	D�� R���Ύ4��V%·*#fP52�O$���=�蜌��mf��xO H`dR����T�D�O}�����;E}��S�'�2� ��V�c>	0��M�dOеj=�V<(B��F��(H�~��TYl�0L6��S��Z��:o�@3���J�UY)�Q�sl�Ti)���RYs�,�J��f��(�R��T�� ��Pz?��Q�5�� ʡ���u�x��3����"V���c?+e�"�x�=̩2ث	0L�x��b�R���2dpwt
���:��:�Q8��$�\( rX��}�Y3�-l��P�Z�8��徇yru��K�'(1G<�V	~Z6�i�:>�B����Z�cXW����M�����>\_�:�,�h�I�l���{�,*��U+�ϲ�6�3 ��?�s�E��k����ql?u���ʖk1��:??ca�j����Ǎ[�B��ړ�>���SǊ�#R	���(��~��j
Ô�G|	�'�s�� �6V[�H�I����vXw�[�'��씄�]�s6Ni����<r�
�ll%�\���������������8ѾD�Jp=[��3h8ϴ��Yܣd���1ޔɁ���Z<�9�6}��`ŵ����g<�qFd��P�5��/����O�����'���'�NP�hFS�{3�j���9�9}���<ҹ[O���'�l�ݺs>�KӡmhC�w��І6���[Ѱ���t�O�>��Y�]��x{��7���� o^�f��WoB-�ŏC%@Ƴ1m�>�����_�t�I'2��(�ǟ���m~w��A: �����)�B��~:�lĨ�nÔ��&�F ��&��m�$�(�O�辯���݉t%��FeY�T7k�*B����	uEZ��Y���>7$�� I����H�7wr�Z��ݍV>�2���������Տ  r�*�W�GyLp@7��eH<�e��1����Z�inȡpA��)�Pl �2�}�"�p��`s���$�VT�n�jݴY�hw�jDV7�j	���؇�@�ou+��+R�v�R�O��2�HhP� "IuO� 	n\��2V��Z��aພW�!���Gஷ�i��A�)�4������xa{eB�-�V�����zt�n��Ma᫰�N��� (3!*C�eZX84�Y�+s$ D`+0 +[c���p��	�� ��Ejs��cR3�{����r-��y� -G ��	S�JG
~e�џ޾�y*�����V�˰Q�u�����IT��l|	g�xC=H��hi��ɠXQ�KI1�X�3vH��U�[V��Zɰ6�:(��ؽ.�#�R���$�^w�ѵ�?2*�2Xg�8�@��
��X��n�i[]}��;� O��
 �I��.�Q�Wh��[��"��~w�9l���P;<j���3"(���q��fH�>�sӖ��%`:��(�qs~�9UD�����1�j��*uU(p��D �G=�W[Ƌ��Y�Q�v��)�bu������5�4��ט����m���_���Q0x����J,�W}&���?���q����ڱ�HbC��W����D�2ϒ��H��e���q�����U�LmhJ��|���/���,@v��q?�B � n���2s�WJּ�C�����\q�-������t<3+/׏��T�g��V�S�R��ߍ��� �q @Ĉ0��2
�<���1�^�ΘC@�c����*<#XA�D̈́�&
,Ӻ-���sB%��?/�����e��� �I�����K������,� 0C���2w���Ƴ)���p�@؂N's��xR�@��Kw�6r���ˋ^�g ^����-��s�<�x����mYc6d$Ha���>ڀ����O���� y�j(o�`�	���g��4�(
�F[�u�w��$���ټ�Wo���e�4n��v�vDB���w�8w�T�P�,+��3y��	���q܂����)��8/dl ���(���
�7���X��Ҏ�nܥ,�`�Y6�\E+��	ԣ�=9:U%
`�hPh�[(�0Fpn	��r�]Q3�}p�� X�����% ���6g~�LC�+���ԭe��׼���	Y|\;�������gJq��3�5�7[jv��Pq�Vn�Z�����c���c�t�����?y!?��?�?��)�|�r/I	��3��8���+y��)U�w��8�<����|�\�o��>��mhC�w��І6����̩��Fr<
赾`u^aՙ-��߼~-/��Z6��|��s�ܦ���Z^�}M; ���S~��YM&r���q&����lt��!����d�B`�h�̸���7o���٧��c�r�h�j��FUZ�W;�YC%W���]]�|�on���&�h��Ȑ�����U�U�ؘ2жlܱNV͏�rvqF�"KG|��)5p��n&���6�Pz�����M!�"R+�8RR��܉Zu%"3#t@T�Mz�u��2[%����#C ͮ�����������M^�l�h�B�AH�}q�h*��pS�~��R���"��GDCU;�_��8����t��˲ۈ��݈*5�x0�zÚ����+d�z�Ï �龊��1�L���ɔ� JF r�x��	r�#�$���m!�]���O�y�E��!��] 3�00��[fsh�^�\��Ѽ�4�
���x䮗�>��D�(�H)IdX'`�|H���� \�"W���,��}�B��W�>��W�� ���&�Q�:�̐�ՠyU�%�l�ӊc���� moO��F��# E�������=� VT��������?��Ӭ
��>�;�o �j�UJR�
9���q\Z����@~k9(���h�2����J�o�Z?@" �-��@�5r:*2�^	���A��k���T�<����U{�M"p��y`��)��ƌ�eq4���D��������N�|�����T�BE��D�J����+g1������R�H���q>4�@e�� [5��5�z���ޖ�������*��'��D+��#���q�F��TV#%:;QkF��sS.����D���A�rz���㯪a[�����!� ������xS����B�u�8�<�g)�a�ggt�S������'HF:Vq��u���Z��zN�2��(<3<!Y�d.I�h��6��Ze��� 8�l���hμ/L�13�L1��=a�~#4ZSȠ�E`D�}]��?�n?H:���~�C�p��6�8W4�^�l2�Iv�9 &jUGz� H*�d�d♆�#h�����=���+j��y�@��Ԛˬ��Z�k~�b�@c>�s���	����͕<�Lg2q�a���c�\۹�
�&��)=&��[�vT�"��{��ݽu�_7���r��8'H��;17?�'j�5�=�	�;�Iڱ�_c�<Ba�����'U)�5�4�f,lHN�����%)�y\�5=���Og�.�<I���~q�^�7X/OH����"|<y2�ܔoK���u��ai�M�[>���[2��p��w�6kT��P���<��>�zw8���]�-�ܪ�S3w�vn�ʗ��>{	���w���ۗ�<fT#�tj�{�+�0ﯯx�XcBE�E���%�@k76����x2��H��t�9q��c�>s��jT-��C��,�DwZX�3�a��l�q�X�������ܭ�]wu�s��V��'�ȏ���<���cٸ��kLi��MO�b����3>�q����j�հ[�C	u����_�����6��mhC� �І6��}kڮܩʭ�r��&�ۀ�Z���=u��G�.��F�Xg�� ������?��Ǐ�	[��Zq�� *�QY�����Xq��j�F��������c�ʨ@a!�5��U�S��^�W�l��j;�����ӧ�ً�Trl ��6˹;��{ ؐ��b`S��r|t*��Q�V�:vOf3���M$��EB �{����������B�NO���V��nG3=���'��Nf�Q�@�Ȋa���]B/f(��V͆��n,�`F ��/��#B����Ȕ�`����n[�r��{@�j$�¤X�׾�6�Z p� rTC��D	��̽w%�M�6�;�0��o�
}��__�Z����GҤVҡ���� ~(���U��LS�Z3J��,b�e��2��2%�p� � h�35DVI���)�{hUʩ�  �3D��n�Wk{ #!h��X�?�CH$j�6�3�! U�*^<�pA�k7& Z�u���sf�	��V�2'AV'��c
{�ړh*��ϧ�yO�(��8�g�"� ��%�:�v|�W���L��"׊��W����3BT��тǃ��R���<�.�{X�--��s��*e���M;��oW�,��u�;?r��H�jI��$��\O>�	δ'�oTeY��)6�@>�y�W����[��m��a���I6%I��� �
����ew��ǀ�)[����[3&4l`���͕�z<�p|�Zڲ�T:�D�CPs.�
Z'E���)�:��׮����:��=އ�F�@Y�y�9 �cS�(�()#
���%�`n����re ���ש� r�CKyo���ߗ�'�/��p��p�s��; �c#�z�Y1�*�_�q�	<�G(u�σ�@�>����*:�z�����r��
���o�#�K˥�g ��J�U�'@���ͺki���BQm�Tէ�@�{���~G.-�x*q�Ė) /������J��ƿf��>P��^��ՔJ��X�B��I3��9D��@	̀*���U�s�,�`mǘw����XD�>I��AUO���(�מe�}��Zb :�~�����~�ɎԧSg�n5=�3\��[ޚ�����x�{Ý�h�n���R�OC]��� d����іV]Y� ��swIL�w��}���:�a�7�y����g�`�d3��^�1��	�;1�iwT����c��(��R�m-p��ؚ�9�g|����T����*��B�K�P��Z�Bp�����h�Tڼ� t��&q�נMT�s��-���PK�	X��c(���g<S�Cߡ��Ľ|� ��[7�33&U����3?�j�����V�5�5����ʰ!�1��<�[�+�����n2�����L�S�In�H�8_����;�𬗊�xF䘙F�v��j�xO�M]�����ڼp/ι>"��x�7i��5J-\�PI~؀alQ���o�lF��ڑ? �Ѯ��4�m��[j�vPȖV�1��g�}y�����*I����N�.M�CU�eVT��k�Ө�*Zʢ��ix6�����g���o}�[����m=ҷ���o}�V�x�I~���(�ws���;�g:�@[+Gk�l�,��_QˆDlĢA,Z�V���q���(�*~2A��A��j.�d����驜<9f�3�#b�PE�
Kl��!���T�B���<(K 2EaS�c���I�lZA'2�i1[%��� ǫ�HZ��~�V�ƱU�j���X}�`ˀ�\VB�L~���6}6xJ�e�]��ȶ,�a���r����D
ۖ|KK��M�n
�� 󍦂j��7�� �x,n�SU��D�Xڝ��紘ag�n�Q)�H�? 
�\�^�[A<@�1H�����Ȕ?;�Q���Z��|�m�c<q� `��2ۡ��*�x�U����x��;�� 1(@<�Ło7�4����A��J)��P�j���eϠ����Ȋ�6A~M�o<ۆ`�j3^��� 2�]�)�R�G�Y�d�q�`y��3��W�;�@��~ ��g��#x��0��f]Bk�h���'3�Tu���ܙLm��Ou�DM_w���G���
0FV�� �p���0����h1�"�j!ؓ�����}�Qś�
}����ǞGvιvP��n��d����8����J�8�*f��{�[���!��Y���������t�ch+tkK�ѹ�|�/�ۚ�q�j�f�`��b��Η����)����Lt].�5��5-�@����"C(\����fPD���#�`�Ae8��x��� ;,�bV|��)��k�
�����HHW��3�x����9���V�` ���p���Ö�ql ud$!@R�i�4�$⚼�]))��Z�՚G�x��X#�'Ū I4��I�9jɆ�
`^	������i�rD� �Z�\��:$���Yy��q���0\̵\��g��k�dB�kC�� uЖ�o�wMC%cq]p�U��h���-�Z2U״�`��vY���t�?J��脽����]R3w	��P��o��q�6j�v9O�OV2H��I+���a.N����+HHf�.YSf��a�82��l����6 �5
����\ ���X3f'���*���XH��a�n���w�9�a^c�T݀t���Qt�>_oe�ڄ1ZP����)Qq͘푯diP:��P��H	�"��1eUݐ~g�a~.�2�[��=27�J��m��e'����*�����^4%b�!T!�c1%~�3�Rɥ�*x� C�a�F��5>��[[�X�����P-�imkv��,T���U{��l1uLϦS���P{8D��W��e�N��>���
0�<��v�vIm����z%�|������9��ȑ�z�<4�'�l�u�θ������Ytp{����C+������A�>_.�~y/7�7r��㵚�!=
s:�k��(<�%�LS��L���9(ZBV���]x�
�q��Jn+U���	��p�JƄ�x��uX������]�7�6 ���R	�RC�V
��Ћ�K�1<��q�a<t�F���:��o}�[߾[�'@�ַ���o�ʦ�K57���EG��#�(@���D�mm��N����?�P���GO��p6"X��5�	D����#V���z)����Ud���/2��G)���x�?&8]�a#�ʙ2ٙIf�ۨ�c��W�F�����K�:�  ��5xY���V7#���O?ef��ݨj�fDJ�ٴ����4�a���S��f`1����rz��|��g!r�XG'�7��D���ǅ�'pZi>��Qu6� /��1��H����[V��V����*fh�T��*4���BT���xC �A�+{�:#��6�}x&�ji�����JCw�v���j����u��`�v��oF��Ԭ��֧�iiQo4�#�5+���@TY#ԖU��RP"�3ѲF��@"]�o��U��Wv)��{)#}���U ��r� 
 L��F�Y=�$L�VE�e�;��#X'¼'���DX��l��fn�15^�-�p�j����j�-=�	z�F���!�nwo��~��y@wS�^�ɵJ�U��@4�ؐ ��y�M%�Ȉ�}�0aU�J��$4P�K;���������1Zy���*o��F Y�x��ח��P��P�]l	J!H\=��.og'�-�0�V�l?��)��M,cůk��0�9��h�̉&gF�:�纵j�J�UX��\�=���@Z�^�j�2:�\e�.�J+���oa�(�2ju?o �n��"}��׌�$�u}����JB�V�;h�j�I%�]n7�DT^�F֥i<��}4�����k�-%�����Gnׄu`���αĶJ��X»?J4����=��YJ� >+�	��� �#	�@�1�����,�[�\��6�e	p�U��Wk�p��kS�����*1��DI'�<�8I��ܡ�������� lb�W�VQ����M)�Q�81[F��H*�n�A�S4�@��W�1"����im���aWMA%��!yTh uU��x%y�Z��ê/h8>|��k\��Z��yO�:�d �zi�����9���k���y^\.`U�l�������]�5�K9�����s�>�����Q����$j�{!x�|���� Kh 955�*��c�\+X�`��ظ��:n9��+����ɚ�\sV����\�v-��V�}�c�4�*��j��e�
}��%�
?ռ	������y�*���P�M���%���Q��X��g6��Y[�Kt��e�Ns,@�9S��ùU���~��G�����DS�1໖�Ղ$����a�WK�q�����Ï��N���3�㞀qt����S�NH��9�2<�n�^$���1�ϧ�)��dKb����Z�3��*1\_W/j���c��w�f�a��8��h^I��O��~X�}8<O#sl���g��!��/����������
����>��wss��X�2���N>������2�N�s��\���;�A^^��ãG��(��ַ���o߭� }�[��ַoM;<:��+��8:>�(�dÒ�T�l$�^�%?��!�_����k�
�!X���� )�F��n!�'�|����`�X�|�M�ZT������~��/�8}�Z�q��ll��.6��;�c���H�p�!����{b��(������fk%ח�ܬ��7�f�;��go=��T+���U�J���=6����h��j�W�\^��o������b�',�!��w�&[VKYm��
�'�A��8� ���J�h�w&SZ�
��4��Mre�A�D�К&b�l� 9l�+�mN�F�(���f��r���r��G�ᔻ��M��#5���=n�	v��5�B_ne2ۣ���	�mg2���
���L��o^���dz�*���J�(��bA2ضd#��x�QI�� \��P�n|�.=�G��,%��G	�Xm�d�V�@N;�-�,uTj6B���no�ɍ��u�x��G���l@&�	�"Z����j�����UKȼ٪}�X8(�᳔�����vuu#Ŷ�ю�=I���u�f] ,��y6I��$CI��鉡���  � &�by�� q�\ �[x�k�vAӸiT���x���A4�&��Yp�f$��,�F��*���9�K6M�/��m�uc� d��4�%� �)k�H\;��i��)�rڦ��*���k����>���%gc�
�4�[��oa��o���۔�� w�ר�5��p��a)�h�סO	��½��^�Y��� ��0bG	9]�ا��9�̷�Ɔc(��oX�`��Zv=xY l���A8�/ƼC�A8v����Z���`�b(��\���8���syPo�eցXN�t�����;$�ת�++�?��C#o���)����P�
7h�L�g��	�S�
喥�@y�A�N�0}d�(p_�7����¼�ߡ����h���mWl໰�:��ݴ^R�)�;�2�����Qd�  �<���^��tT"<��������k8VS��ü�DU6�p�����$�'��ʹx�T�9����M�9G����X����j)C.U�e�E�ZC��L��I%`R]w¸X���������U#0N�p>����u�a�F�B��kbj�ʻ�HL(�p�D�,�������n3&�Ɇk!�M
�����^�e��J��o֜x>�-{��kS�B�BT�>��
�'qc��^-��529��w���kU'��A~3j,���ɮLFc�ត�W`}X/�NTX�
�R%&�'m�L���c͜�Q�����bKu�ձ(	�y:̌�]��PS�E����:^�
M��2�U2�<� ȋf_�b�JTq���mms�&�� ��Pِ�}">��*6��Sh񔒈�\��g1�~1as��2����܆���՝<��Sy�Żᜆ�XE^��ƞM���f���Y�L�sP���$<��;��_�j6�0�<fȰ}2��ۛ[�x���{|p(;̊��b/iU�5�Zš6�P+�~����G�٧����M����1^^݆g�ޯ�ondx�Z..��~�K������Pmsxt�k�fG��qM�J�]�?�۷T���;��Y��:
��?����o}�[����o=ҷ���o}�woPG��<𻓣��� ��j睽}�����d�������F�a����S9:>�GǏ�у5�=a��������Dv��2����%�~�Hp�*n�\��Y��!l�/�n������'����t<Ӱ�2g��25	�A2h�w��\���&��W�d~wG;�*��?2P	 �U��^)�`�(�T�0�P�۰�?ؕ�ͥ��������?�H���	̍G{a�v,}4W"�*!l�A����v� � �6�?f'`9h�@{��T�J��+�%j,� p�Y%?�j@X�7U��z����R��o��$�l�\��k�
@. y $\���.U 8ދX;��h���ɑ�DɁ�b)Q6����Z��c����[z�C!3��� ��Y����K�����јǕ$��`��t�U��8\�G��,I�C+�5� ���Ui�zA�葇Fp�jy~�ٚ�V��c�!5O�j,fOVѾ˫��98�a��c˹烔��2Sk7 '��f�HX��^l&�����������[S�hpu��pZ��n��Nh���g~]P|k�*�ĸ���<�8� �jU����:huw[���Y>�+�,pҤ	�w�ǹ)V\��E #��{	jK[�9A�1@�ն�U16�1n��e/D� �|��Q:$a.�Ru�W��W ��U�Wa]p�\S�~A[+��
 '���� �격N�kQA���QW�2�R�5�l�
�����n��+���ƌ�sWa�f�;~�냟�оu����i��~��@$�cco��c�I�9<_΅Bj��<&V�M��r{#o کT {��*��&p.��=�s�G��@庄�X��ƪϻ�#�r�<��z��W WI����t�ŢV��9�W�cl!��T��\�TE��UXNk|�{Hc��@�hִ�$W���a�v�=�.��Q�����s@%c���Ȑ�B�K���(ձ���e�צҁR�2u���,T@��*�*�V+��9N��G���iɍ�\Y�E$�[�Zbj~FG���	���V�����y���y�D@��b�¸#��Frc�Kf指���t�(����d'$3�w���&�3���0l����=�f���ó�J�-$��ca��xd�A�2�W^\\P)���˛�lVJ�����5 $T{0�)�Fp�{��mAT�5P�b\���@��$������pF+%����Д$��z豺U�۴�œ��Z�Zk��y+�5�#j�h�ŚE��;��� ��ڎq�I��D5shJ��hÅ︼���K����/�3�����{��x�@A
f���"�)\����p���=	����J�yҨt� ����x�h�$�>K�����,3g;{f��#k�v)�g����_���u�� �qq��-�g�l�(�t~u)�p��4��0^�H��������4\�ax.��:r��N��8A�C�-��6��7�Ͼ�'��t��_��o}��w��H��ַ���[������0lJ#�����t*�G'���g2Lb�ݝ�����oÿc���wh��y�ŊJG�}�t��a�}������������W���� W� �|���?�R�<y,���܄�*_������pS ��qB�6j���h"ka25@�*l���9ؗ�����Y `|X~a�D���� �,`2�}*�^��F���S���~&������Fv&�p��j�;�M)=�5�{l���SP( .���0|'lb���^Ӱ�}�v%�I��k$T���P.�;�  �p鐤�{�3<|<b_ac[���GC�4*IK��Z���א���(w����с�x�97�����ݪ��@M��R��&�W�:Y�C=N������(P��V8^M�B.�u8���,j"��Q� 5,[
ENZ��3U�A¬�V�b���=��z�n�#JZ��� �� ,��F�X��. �؂�ҪyK%@�*�ޘB�!����W���" +�NI����W ?P}��\|�b�h wϚ�����������F�ƪ�i)T��2j�5 z3a/������$�{�Z���LN*x~���
�EfgFp5j���b���k��$h?��jøE���;禶uPx-	0c��(�h��9�s)j��!���`�t_;M������[��qf�1�b'��HI
::%C�\�n��'c� �IP���W 2M5؜N\En�c�f8�w���ʩ PB����N�x��L�0�|����x�^6a�6޺��]��/Jn+��=[���E�X�:1��z+��5$�� t�'B=�v�)WUc}�}�~O��@�<��Զcʒ��I�1V��(6��0�2��\H��j���? E�Ǝ'�|���2�-su��-��YY�J,Z?���� �s��z`#ǝ>7����`��m�&�|�q���a>��ќ��|��GPꤍ�!Q ��Jm�<}=�>�T��ٶ9N'�H� �9@�ދ�'q��[+��y��H\�qJ"[c<���,$7��ts��<(�I�餳��x�_p��*%'�����&<o+�`_!�,���-<��i8�ƊK�$(j���z]'�V�
�P��&|�KTܲH���W2��Q���1VD���D�v�j�	�9gh�P���6��Z��u��p�}}8�>��6Xe���\ʺ%�p϶w�1'}�l~��A�+��lݒ���k̓�b|g6%�P���%BG1UV��U��\���
EAȳ�9}-�{o!Ϟ>��#��i������r<�y�-V�"�.��)�W�����`�)f-��ĳ���1��ҁ���p̂T�����]���?�Id��@�X��O��:��H	���+���!����@�}�����ɣ�O���1�g*N��߽3ۣ��T�}ɋF�s{ң
��^���>��������b������o}��w��H��ַ���[�N����+����2A�|.7a����Qz�ð�{W^�x��"6ihGa#4��Zl�܂�Ad���?��?����W���\]�pG��1§a�	 ���ͥ|��W�a�'�oo�	}��-��c{�VW�hO��uP�S������U���kp��L��a]��aÈ?�Ǎ�*�TD���T>��3��_�(��Oa3yG��`z�}奍
l�Fc�^$V�Y��9*�7�   !4����=CH����h,���o�i<���3=���B�����E�T�G�� Y�Yx=��->�@�&*S�\�eF���}�M���k��/����V�Q���!*��9]_]���F3�)f8�8Q����dD���y�UTj�4��4��|�h�~jA���ϮA���,C/Ed�G
��앫���i�Y&���|- �X�e�߳��GI���P�t�g1p��:�#���w�V�Ce@�o44`'fe�+U��r�����^�N%N�,�T.�wՑ���Ǻ��C-����j��w̉��9FUws]��ݎO��c�I(�H�DIY=Tt	�HeQ<8�np�� tV5D�=�ns5Di�F����&5`�A\��Mk���$U�܉Wd�[������H��QX��H�8��ƾ�`Ѷh��[e$_�x��vGG��۴��UJc!F �`x҂�~=�h�O����������[�` 
�R��M�hYc�����9=ǔ�H���>P��׃��Y��{=�9K,�"z�W�܅Ts��K%|�����˚�mK칒�B��~��y�=�Q���z��a�U*i��Y�9igw?��K�5iϝGJbx���S f���ŨmUٹN:����bèUpl���x5u �:���=���m��<���x�����|=�u����^pe��w+h�k�*2�-�[���ؤ���� bcY~^nKUGu�;�N:�T�Tl+%��O��}�U]��W%��*a|\�����nc���e�6c�yw77���.��YB\���,���:V�]f��$�g�ฺ�����c/9?;��&��A�ۖd���?j�Ր F�`��$��њ�$��dU��-�,D��@Uh�|P���
����D)8���Kp���Rk�NCh��}-y��k}e �D�ϬU������5�ϧw�}?�g������*��T�x�g�oNKY�籝���|���Y	�`*k�"�� |��䖉�d���麪�K���g	�%����)�|<�.��d��_�֟,�~A��mxV;==��>�Lnn�H����֜5���P	��ϒ'���g����?���_������p6i�,�4���>�{CT�*7�{	�$�1"�G�Bvw��?�Q�ַ���o��� }�[��ַoU;
���'G2��b� ��cV�ku�����#���X��<�`�/=�kV�]\�p�s��+��~�3�կ~%�|���jcS�mlb(i��rU���@��o��>c�-�8v549l���D�F��N��
<B�sFk.m�ð9dr}w��A��h����}p���DW`&%�f��uu6k�_����������aә�@�
Չ3��%��e�i���5���@B���_@I��>9>���Vy^���1��ϡ<Ū��J�{����@^��+d@E��
�:����	���]�{�W����5�*���=��?����PX��r	��M��H�mɪed��p�����@�o6�X=
� 8��|�Wl�i˒d
��=�g(�t���M��?4U�"�`uO|�(����5���(�
^q ���_(�064!6_z�5�k�w���h��U� �R1<��ǻA��5��U���	�Tԁb(���)ׅ���:$�p�^�;{H
����X3n���:i���X�jVv�aqSU� �e{�����l2EpWE�:��w�V� ��\��N�� SU������>bl��m怨�X���:(�X��Ұt�-�jm��`�c97%E��)MA3�g G��qO�C�S����аo�q$<T�c�]���C�ӺU�Z?wWz��Aft	-�����}dV,z�Ґ`N����U*�qJ�4�/_�]9���fN9���-���&P��� q����[�%|Z֋xВ���v�n=�}N�]��+��c��D�ۑUe���1A��D�j�����9�ű��G5�(���&���Tj]��lZ�eP`�� �3��Z�9d�
U�0
�"�J\!�����
��4���z��g�9t�	J?ܓ\��������d��t>r�GTm�Fi8P��2@w����k�RDjg�N�BE�@L��k�+x����{��]��ec#N��:��1��{@r��Y��Z.h�j��PrE����=5%�������R�I{ʒ����
#�zT{�EcU�|"�]U>scD7�A�����l�30��ZW��s���MS�q�|�
��-3'$|΃�e�Fܮ�,�`FP�dW]�RS}�b���Iɨ���ZIݬ�=AҔc	D���B	t� �4ܟ�cYp]e�*\��e���aDA��ex/�(��|�K���>@�kdvW֟qgޚ�	�����E���'N�32"cr8���
�%y%����1.�z���un�E��P����������>���?�!3��ְF$��sh����V���g<7�+r������1�gV��u���_���>�܆c��g�ݽ��������~�O������ϭ�c�y~}ƣ*x���� ;��p�%���/�w��$�ΤNc['*�7[x&I�q!óiB�S�7����a��e:�̋p�un�q�շ���o��� }�[��ַoU;>y,����v>���򁜿|%O�>�=Vtm�����	�� �6����&X(�]����+�_�˯�[nz���\�2/�"�U���eI���/|H`��wߓW�^���$�;�1 l��n[Z5�VFz��i ���(��&c`��!K���'n5������$|�7������A��?����W���<}�£!7��� 8�d���-�#�*u�Y�2@�j�VS����F�Ox������F�¦�3�cu�(' 6Pю�;6ȩ����A�X�U ����T��R�v�6lJ'�A�j��e@0 �h <�����-����ZlǶ��ahI6�P䬌�� z��n`(6�{ӈJX�,�z�<�H+fq���1��f��ֺ �me��U��D�{��`���h�nHXUG
6��aި�4 <�ZEA�I!�ZE|��g�b��w�5�}2�� A�XO9�S�$�<_��l7M��W�w+�'fSA�S�ר����y ����ኬ��pл�V��� �4�U
U���������5�\�<�� p��
 ��v3@�àU;���J��y�	Vzk*���G��*ƭ�X�k@��|&.�U�;|�j��@�6ㇹ:1�Ӂ~V�w*����]{��.�r�pN�X+H� ����bw]m�)o�a��R'"i��sՌC�J�y���j���eV�F4��,-i��K����1(���S�]�����\�>��U���O4��s@h}~f��|�%u�2+2��ǀ�^+�3�J�C�����P��_��%`b�5�����>���]S#>p��U����>�d��҃YH�N���a6j�d������ۿ d�4�x�<�-������A��LK�w��EN^�G+�5� �by�X��\a`t��&'Av�p�
�
)
 �[U4b�����h¿g��ղ�� �Ff7Xk� *�i)��pS)`��Σ�)!<�%�i�~ds���G:�>���`Y�h/犺�
�����Lx�~�o�iU��C_�v%*~O�gGX�wN�u���9���K��}�y��^s�y�eN�O?��5�u�����tqv�ݴ�C:�����ds^A�MA"� a��<�O�����j�	N�m��|��ύ��b�(��2�,�b���C�*��4�"��w��M�9�g���0�q�u��5�g�s+����I<>����C���Z�i� ����ʐ�+ɲ���<���w���G���ub}�ڨ5(�����pMF��*������������Q�r浫#���������믿�Z~��_���[�4�cq�ܒ8��!
wð6��f�A�����x[���:<�ŵ�@��(y�B��,�r
��\����NK����O�'�6X��'?�	���Jj�\Vַ���o}�N�� �[��ַ����G����K���{�@4��Æ�4l�>�$�yr"��>�,��>l~ bs����Pll���ԗU`�{fy��g~����O�~�&H��$�/E��Y+`ӥ�j�����\���+�B�̡
���Ɇ`��>�Ga�ͤn	n���UǨ86��4��h���^G�¦l�w��6s ��zx��z�Z~�������O>�X�e6�S�bs^�j̚ŶK����X�����>Cuo6b�0j��`7�n�X��I��,l ��{�^ :0�z8�%�W���Z������9i��M��@J�po,T�	�@��!�X�mPt6T��������I�*��'�H��K��D�*���<~��1 ��0��,�-XD�UΑ~w�i�`1U���e8��"춨n��d@5� ȩU�u�y2ѿ�J�R���,�<�0����G٠��j�����
��̰u��v�wZŘj�? b���k�q�Pҁ۶Y%v����s#el�$QQ���U�^���V�� �o` 34[�!�~^ m@0�f�U𼓸��nH��U�;�׵�rR��-5�Udh�3�X%u�~S4�Dzu�땁y~�� U���r�.�}���mǷ���"���:��=�fxX_b�� y�H 	����jS>�j��+��j`�n�-`=����	���	�,QE��;3(:6Y
H��a���(���͉+k4m�*����M�* ��:'\
#h��כ�Y~�u��O?Om����Í��hM���#/��pب#��n�E%HV5���1��\6]i
 *�Z� ���0r�<����
`7\�a���\A)�V9ǉZCa�*q-R�����s=��!�H���zh_e$:���r[4��
�
�[Q��E�X��ye���YeސC�J�l�s0�Z�ǔf�h@��E~��D��)�[E�!M#�Z��갆��W��ޒ����wR�!��i#%I�����D����mo횶vW>nu�S��<'4����f@|�g���ץ�YL~����@�'a���ޭ�z�r��]�)���9����&_�+��
W=�K+�����	3��& y��q๡(����Kn�?b�~̀�pM��������@�6�p7���v�>#)���v�c�:�#�S������-���t4�Z�(a1�}�ZkYx̀��e��Ox���V�I������z�"���ۿeq��zZ3uHO��y�eAC%\;A0nC?��L����Pä\�i��1�����<�BNO_��p!;�<^�����OG|�F�a|-�\�"�!B�'$��(E��A6a�e5��T@?y�$<�����֌m�L���*N�uϨ���������(@��%�Q��5�%�XG��+(K�Fk�g2<�1�*�?�p�WW�?<�o��0��\�@�����,��jK�Kn�������(�½,Bz��҆AQ/Ø\Wqԧ���o}��w��H��ַ���[�N���<l��Zi� �(�� �w���bMPlTg�q���}9>8b5B���V�~^]�V���h�F���Wkn8g���=lS�ϯe4�J����$>��sy}~)o��N�y����:��֊��x�x�;ȃ;-lT ���r������t8�3�����N^�z)��/�����#|�g
����4q0�U���}��17��B�w���m�&���k�!C����������<�}����u�D�{/�p�0����,(:7%ű ��4�4�T�.�5��[�7l�h�a �j�q � H���q�y���Ak8P"bgw'\�!��/�ι	{r*B�>{��ۚ9�Z����aW3��p"[�!�FnB���5E�U�+�����3�_�<���[�p��*a3��b���
,o}��J%J"dfhFK��L���3[ \S*�b#V�9PB�8c��­~�RR�ͧ��ó
�'l���)z���wAz�7���Ƒ�5Q��WeG���j�mlp��C9��A4 # }�bʿVT����(H:���H8'��r�!N:�x���ʶ͊P���ͦs�&�ݱ�bI�p*/䙫�^�Z��--<ޕ'�sL����ec_W������Jl1Xv��w�k�Y� b�!�PD������,	�;Tajţ��J$'[�Ĕ�t6+���Z�4��$��c�T��R<��r��ͦl�LϦ�zm8j 󆨲�^�$�S�qC�Ѭ����zǝ���Q�8	�fPD�B�����4ׇJ0��/�x>�r�j~���ʁ��!�����=ۚ�<�1_�����>>�*��SN�躠��XS�����!��m�t�k?�Nk�T~=8�͚�֠��[���8i�Ƣ֞͏���۹Tp;�u�� ��6sC[l�)��v��)�Ԗ0�O�DܛD��q(%F��P���e�z9T�0�̏�U8���r�
��D��$ ��k|C��r$3��M�ҕ_����"�op�Q����*��qWmh�XU%��|�?���h�s�y���g9�L[�I�3�Ubc$jTM~�{��ǯJ�({f�q7��$���f���b��6��U�Sih7@���\��p��Y�YHU�3y//5�,&�Ya�v���Y+�{M7�()V��<�m'l�J�Z� 3��7�Dy�d�p���Qy��+uµ-tPRN�ԣ�n$Q���a4�3l�!�����l�=o� �ό ˨���䌍��zy{sõ��~�c�������r��U�N���UD��J�����S񬖜�?:ẏN�]��p�Ֆב�W8>d�_�g�_�������bg�#���f�eN��d�c]Η��,L�S���>���z�PN�N�O��|���r��zyO%ԥo�g�d��Yk�\ӆ+/k�X���#���3ړ�������<<�]Uet.�]Z�k�[��ַ�}�ZO���o}�[߾5�œ#��F
�t4T�g����&h�l������=��J��	<}'ðA�i{�@R R�
��2�mc6K��X�� f��-���T��;Yܭ�d� ���}�/������a�Ϟ�����rxxh�Q��q�hЬVu+贖���3�X���]����¿�&������?���������ʪ8����V�z�-y��1��|sJ���豂a�<�!��v��)��q6���	��i��>y�D��M#���۫��A�����Wr6��V����f�?�S�t����선J`��z��	����?8<��Ϟ e�bɼ��՛
��KT�.�׍�1�GQ��'O�b����&���l�?}��{ߓ*|��_})����� ��pݖ���εRr8�P+ ���\l�X��7��8*���T� }j���1���#^�����ZY���)��PE�icq���Os%�G2?��
�Ě�j��mK�3!�R-	�; Kp���Z���Q
��RX�@�xe�V�#�|i��� \n.����.̣0���+�e �H��� ��8|?*0q��1���_�{^�x��t��y��s�����*ˈn �0_y^^:�е0���n������й�;dQ��F�)[�S�w"�PN��[%IWQ��\���a��6�P֪v?W��j4��^��O��"�U= B՚j�*m(Cx�������Y#$�{���w����@k��YC`�h@}��� ��r��+��z��x����V|$�6�!pӨ��p�5�`s�)'���z
"I��W���E��xqН���\#=�����#8Y��c
|�t�A�߳"��L����,x���U:.�[�	�vTFo�:B%���3�"dKJ�\ev0��e���{�����yB�T����J����������-q��RU��|٬U��C8���
�U[��m�x��,ѵ6MeC�z�1	2����jύ!ɀu.�c�(��4�;��{~oX�ӎ� �e��������Yj��� ��*��C��5��ǳ�����R��gl�������r-/6 .�:���$H|�t?ퟲYW��<K�������<����{��Ę�u�_�
���]j�t�(D���{���J��2o��g&���7/Cy����'�ս\]��P�L� ��n>g��p���>t���XW2�����i�%�//���=	��"<�����˗rv�:<��c�ܱ\��s�.�ru��-(JI��wU�Ʈ)7ZbY��\W���dTUJ��:VUJê�(�Q���D#�=x���@2�w�ނ�'����A���Tt�9���*�CxΊn��t#�7��{gz��#MG��r�d�3�q5n�qgx��/��
��8̅=+ѵ�Tu���cM����"BqϔEI��ͯ�?�)�X��w8g|�r�g{-�,�{J���5ϙ�w��([-�A�۟��G���%���gidO,g�v9_��j�FK���pxt"o�������U���0E_�I�2��W����/�o}�[����k=ҷ���o}��4lx�V�+������� ?�"��eD��1}��Y���v4V��PX8�p���~��{z���5�b��d���" ��|�x-¿����rx��M�o~�K���c	�����˸�s;	�L�11`U	���# ���&�a�_�ɧ�}"?�������ǟ|DU��ѡ��vx��0쏡*X 8cc0 ���� X���`�}�����yK�?}N ���R�������<����7���a�>F�
��Э�
��2���&��^����j'U7�Ry�1��@��Q�ҡL?���r��5��`�rr�H�>ݧ�Ǽ�.��掀XFeπF�}�p�U���2��0H�-�1	�}�QB��
)�F@��+g8�z5'P s��f{����BƬ�r*`���!���Fm�;_[\�Xqk*�GU6y*>���A�̆�H�Vys ��ەYթW(;ACЪ�|��W����Y
��{UNq<���a4����������qyy~��I��\@�190G����ם��hvA<�X5��bVC�<��'Q�c2[����Q��U���� {�>��;�50�� ��w���pX�N��8���'~}�J�B,m���y�9��X�:xށ�E{��Z�����|��?HQ'0Հ�fgM�L;v \����!^��s���j+12k���+�5�J�d��Mm6;
ػ�z�+ ީ�~��9�c1�-�VEZ�Y"���Y�^͂i� �5�UDIks�q��%/H����Z��k��$�L��T<sa|nsYTƿ��]i�5ʷm�n�}�ԀT�W�l�v��g�@3^�ܰ��*��qU��%�R-��5'qP����]����g��c~�Ճ����nW��~Ql�֬�����DO�L����\ܦ�k�=>W���p ;�y5~\�҇�#-i �`%VQͨ��:e�Ɓ�5�Cɗ$f��7cNO��2|Wx.�9(���l��]�x�l��zεKҫ�!A�c��O�'wR����-)�q|��� �ݺ0,�𾔨Kv��9EQ�׫����	 ��p��߆u c����w�yJ{%�GS�GC=�$Y���d2c �M����;�3"i�;З>�I��c�������V��~��|�ɧTX��`8��,��l���
׍���Z���Qr���������������LM��3Qw�v��L����ܭ�X�g���^�[ژ¢u�`�*\���~���'��{$6����j�ϑ\�`;:���d½vT��ȶ�Jd�A��k�������F~��_����'W�TU�P��YH �.�>He�ÓD:p��l5�c����q��	�%���3Q�y[4*]�g��#��?X�fYZFQ�s�*����˨���o}�[����l=ҷ���o}�V��G��,o�g6��a�ae�R`^��уot�qYnh�����]I�*�,��XQ�I�%SY�&�xQ֬~ŦL�;�X%eF/u���-�iUmiр��(�y��X���߄M���S�U�w��{����aJ<�dg��!�'��?��0Ŧ�*�O�~)�/�������Qؤ��r~y�\���z$��7�M�vSr3����-*� ��H�#�h��<�����4c�?<���ɋoq�{zzJ�	|�|��BU�6���nE����˭-S���rc�20bHBi���B'*��2¬�h��x�dwg~v4P�5�$�|%��]y�ⱼ��[$� 8���qC�ao�0\ӡ�>���[h���	�8Zʀ��H�m�-����ᯍ\�/Я<���	\��y\�kSV0�y�� ڢܡ,CpM�$j�Q�h�+�:6e(��
e�c ?a�BE�Z4|A�ߢZ���Vx���Pa��y�
hJg��JpUc�psV�
ȓJ�`�|��j�@e�/�A��V��}����������@'=���X	fJ �ڳ��,@� �0�cT�
�`��9�CL��DC��j	���yQ��y8�H �*�� #��m�!ѿ[U�+`O�k��BeӦʝ�@V� 47�s.i@J�>'��Fb��n���j�$C�u���w�s�́�n.����Mux���yD������.�; �V����p�~Vi��-8��ֵ<s����Oi��N�T�C`ݫ��3$"ˎ(��hUk(�R�m�=U#a]�N��㑪ݶ���#���*��9~bm�;�8���c��L�1�	�0v���V���C��� gql��ol�J1w5u�j%�ʖ�������)N�Yo*����[m9�����n�o怈*G\Mñ?��r��`i�Gi����T������k�QT �����1SW�a��U7̍-��6Tn��X�!{k���5��8~'6��Qb�$�������Iu�B�R�V�qj�p���$�0)�����З�'8^�)������֊�QIfפ�9�"��Y���7^d���%����{'��X�b�툴`����@6�qܓ�.�Pe`;�5l��~")�yiJ1��������jvV'�Yyd ����qժVr�'kј�+�'j�z��u���B��=��4q�yp�2�faV���������灋�]��	�)qԜͳi5�¬��u/�iI�����q�g!��~���9��U����8ѥ�O:�H3�I"'Z0��(��gܘz����	����J�{XPf1�+6�����:\��0ѷ�pOvҌYz�X�;���5n0��w�x�	�����{,H���<�����G�?����w�"g��T����3!��!�o0'R>�C�;�F<O���j��1�~�y��ρ�\/G�=��z�SN���
[���w����~��1���f�p���]{y<;�z����[��ַ�}'[O���o}�[���� �!��p�6\;X���	6w���J\�������3n�`�[,u�Y��8>/�L����S��M���3�`�['/���ٝr�8&�V˹<}����+��H��z�Rf;{�HtE���'������@��A�eE?cl�@>����>�Hnno���B��tego*�����-,��7x D`W�����9�g�܄�a�K����e��Ž�<�'O�ʓǏ���bN����Wg��o¹*������a������hAhV��j� ��^�m���~yu�M5%����,�5���vu��8���h��jC��յ\���0l�ww�����p/_��Zt��ñ����r���`L[��645A <;au� J��hg��� �o�o	� ��yBc���qR�����I:�`;�^���8(�3ݓ��C��b�i�.:�9-!�E�g<�:!�j�u*B`,���M����g%�Ъ�ùT�	�&@%�Z��f~t
csB�'��vKh�Ru�^H�rF�q��� ׍��@kͺH ���n�����S��$x]�
ŉ���Qv���!��g��P�*H\]��=�ߕ �cn���U��֫S=0+;�eۼ��\
#C]��>���m%ru=��Gs�n�wc]#�R��v2�[i���8�����zkp��xx��[ù�Gn��!9���Uy��Ө	�7��DI:'���E�4�~+v�m��E��V@S�aU%��'oK7cĭ��+(�-�(%�� rS]�~VWEDB���[5�4c�Ǌ�٨��2�����%	��F#U.]��f����ؐ}�PQC��T>�}|7j�Z��#�6j>��Zr��hWa��!�y<"���d�]�5���7�K\��������D�7
�u޻-�旨�~���T����<��p?A��'Ƥ�:�V�V���(m�B��u�	#']�4㚇��c��FHn6��G��Vv�',���ƫ�~�~�k���c�t�OA������@$P�bfjK�f��>`�T�X!��0'ݢp�g�ȕzlyX��>�]��3��`_��O��#�a�4M�((¹�jUI�`U�@�l�d��x͚<��o���o�H��)��?����?��UH�µQ���u��<�U�B�L�cڇ���2�I�N�k
�ޓ9vq}�V��ص�#%p�kR%����T��ϓv]�b�J�G���5����mx�(�����h;���kޗV�%NM��\���[AMó�ѣ9
�^|���o%Y^s�˦C�S����y���՗�ȗ_~)���o嫯��O?�"��Udk �?��
�
;�	�i*�����+��Hؑz��q�Ts�rg0��d�G�����"�!���n��F~�眄�r߮������r}�������ӷ���o}�ε� �[��ַ�����䝭]�8��\^�r#v����W�7 8Eq���}��2S+~���{�ۻ�mB�v��y`;a��h��j�u��H�K�QB����9>����]]ʫ���ަ�Y�H��r#�a�VPڟ��l���tGv�3Zp�B����^�����P�~֯_����+�@�����V"�c�L/��V+7�_j���*�ɝA�`NǬ 1p}u�����>���}V�ߙ�ʻoO�,���5A�b�*��ހ����n����_�Ztο#��^��P�N8��S*�qč>|ŷ�F��D���ON�q؄�����N��x~ɍ���w�������������]t2���%- �T�b l��G�0��#y��w����T�� �9�A��� w�OÚ(\/j�����}�����D��W��c2��H��2:�:�{�r��~u� jh
X���m^��E���Y/՜@1�&�m��{M|�DE���1�Z�h��Y��k��vK�@UZa TI#�%��ps�GK��r���6v(QU[hvč�Y�U�vmj�8����lȱ�$j� dA 
�N�w�����6.^I�V2����	�B�$�q��ǫ��m8y�����'i��[����]��3%:�8�`��n�Ur�O�<�Z�Z�4;�7��1�W�*���"�7��5
c	vW
�k:�$K�X*�~�Ǯg��&�L��Rɛ�*�!�D�� ׁ͚<�yX�3���{|�W�����}UF�A�]Pޯ �VaS7���W-��!�&F`�±R5��u:�ݍ(Z�|�5��LZ�,gp��0!9����� >b�Q�B���{�w`�����Q��YS��$�M1�ǅ?q�#�BE����=~�Yz���ߖfYfA��|8[ 4�(�Dm��'� �u���(`���Bj�#�E���+*�y������ӡ���,��7���IlsjK���F����idCA9 s��qj��m��A�,µA�{�^5
^�S�����uKl��Dw�̗��r�k؛�W	���z�)��ɦ��i�����pO]�Z�))U������9��"%�3�k8_~&fn��}x&��U1����V��>*�M�q�َ��3�T-����,�2sǞ�"E[S����Q�!a�� x��O�>e�J�ż�x�B@��^�D�Z��!GcW�j#G�*b&��y)Y(Y�6�n�Se<�\���t� �dd���ڧ�s�}�j���}�f��V����)
;���dqB��'�~,�=�gO�Q��灯��F��/9n�?}�?�����ƴ��D9�<��f8��
���B���s�,��3>��3������o�V��,�靆�i��`�T�`#�-�uG����HO���&{��?���5����/��r~J�����x.7s��\�*$�#~Nx�"?w��[Eu�Qܽ}�[��ַ�X�	����o}�۷�a��;o��o8��T>�����ײ^mY����-�f��)H������Y�E��{��-y��;���J��˗��
���
�(0g.u�a�,�W���w�+����������Cl��q� �Q�_c����\�-�է��ƙda�_s������ )y�VG��	Ȝz8/�ֲ	眅��g?;b5΁
�p�̾ Lp6�f��V�E�%�����	gZ9�bN���� ZV��:y+�B1t҂�a��nC%���1�p��q� ,6�,���P[�	Pv����w�{�i�`�k+l�����06@����˯/~ ���,C�:(��y�6��u<�h����P��o���N*!��N|ƩNJ�����s���ԟ����ׯe�Z6����)5�����5U5 � �о&�$)S���x���wuh1[��}�����	�X
��`Gи�L�,��ک�	����ڞ@�����W�9��J�4&���V�oU�C�&�i�
�#*�Ǵ�����.@�բPc��Ŋ��g�8u2T�:��R������h|M� ��P��(�$���M yM;@{7� �{J�݇�Gh �#i��l�j�K�Yn�7Tc���@���Fm�ʂ�e��)B�D�>O+ң���A~�Hs����J�����/nB㳘�cn�S�m������[f�M��ϋn����!������Va]۞��$S�Z���Z49*�O��B�����ݿ!
����j
=���8��Y��:_��IWTv-p�?�����ʟ��Nr>ȹ1Bϳv����][�<rE__�=\�8w��[ns�Q`E-Ʌq���?c˘)TE�ℕ�h�|5��o"��J�,5�4�Я�P��QQ��s�ߞC�
���	����9 +��5��t�d� �"i���a�A��KB�,�\��Z����p�~�Y ��"�V��c��'b�U�;��w7W��:�$�*��N6RJ��I<3`��� �X2��.<�m+�"�"S���"�~J����pyp���T#��rς�i�4�08�	��r�@��<Q̂�a�O�������&b�l�*�R�������T��{[����%j}��|�{�+/5��!����T`q����}��8!yӴZ�b�9�+eD;��=��U�?��hF~��J׊Ҟ}��$�1�m�Z��������E3wr�}yKU2����ky}�J>���U�i� ���������d����3Z�.�\���\�҂�y���*l^�ж��˱P��cK�ل9;\K2U�<{���n�ח��������ԏ��"���}y������{|~ø�<����+қ����o}��w��H��ַ���[���{��@~��psv�L`;l�ӗړ���J y�4S���� �e�x*?�������e<���~�;�����~�����Z�'"�왔I��pI�U���H�˅���ȋ'�h�����:������'S��J���i��.����}��wd/����f��"¾�s�a�G��d6��7Kn�p<�m {���o
��ߡ��+������e �{e���눀�k%�����!�+ �"��s17��~)ޫ6�JU2T܀&�'7ȗ��)�q��Xv�VkBa�.׬HT�$.�)I���@v��	n�z����;�֜�5�\+E��ly��c�����k�l`נ�ȋ����W���ޓý}6ܨ�O5S��"m�u��j�������r{{o�4F� !ؖ�:��=��|}zJ�U� E� ��_T�?�6`e�<���6p���H��
<����3��NCᣈ*ȔFS��FVF��If1x��,�;�göj�\<����Z����Q�Q+d�@����@p�� �Ovf�����[M��я �q,��Uc� �l��U0Ջ���<4�s���u��jY�y`��!Ҵ��hhvt�׺������2�1�-m��=�@�&�$V{!�eHސ:8.��j�6Ue�!��0>�q�
���VBh��u�Nx�%f˦dpLP�	��샚s��H����6��m��DSK/*Vl�P���AZ�����<]�6�E	����^��6�4��v�8&ki>����Zd��C��|��$�tL��	�V@����J��6@]"V�l�����\ȕ8�R�)q�R?X�QI���'Zx�X�c����O��o�f��˒y'4�)�FA�/�{YJ��&�\�����
t�㺤i>�E$�j�V�[��&_`�k���xӰgS��<ڔ���vyUǊO�P*1��>��n�C��4�Ĉ�^��� ���Ǆ����#%�O�d�U��=!�f$P��9�����|����m�<�r�<6�)��!QA��,��l-���*�|}�f9�U�4*;#Z8v*�n��p����c@�� y̰�v\�:P�� ���H�}�]9D�G�GCY ��D
�/$T�L�;T�(�3�l��<�g��YW��R�TfJ�����n��e�جa:�ڗa�U$��� 2��~W��6�CٲoU��*���¹;�B�.�CB
��ԙ�����Y	���>/z��h�l�ZJٝ���Ue��9� <޽��Cw7w2H�T�]�\I����}-����6p����4�٘ϰ��#rq~-/_�R�L#�z���9
at��� i�����ޔ��P3�L�]qݩ8��WǚD�s?����B&�9����	������P�)�%��vM��x&988 ������3~fR妠�[��ַ�}�[O���o}�[߾u���k<{�<y�j�cS�P���C9��9������&c��E�t�<���Ǐ��_��'2L��T�˿(p�U� ��թ�� l�PٻzH�`2���F2<����RƳ)-..o�o�\�X=
�/�R����5�9
$�a��b�@���}9��'�s}C[���W;{����L5H�����3�:��� 5 ����x�M���6�ۊ�%ػ���*��)�:?���{��D?]�\��nNpi4�t��o8A8��da�����熍>�+�a�p�&6ۋ�Z/�H"�S6@7R˜W U����,\s\���K���/��˯	�	I �1{�;T,V���	��A6���;*N��-�0AӪ�L�CU�<}�Xv,���l<%�4`��VbV�����n(xx�藢���c9
}��H�cQ+"�ɾ�C�H�C�_���(\��X�;6��l�Ҭv��_�V��NV �a]�(�����E7��oB�����[0��k��������j5c���U��[��n2I��;�TAp9&@�
�ĀL ��������!��W�x&�^�6(;2?~WE�Nc.2���O�G���Y�(��Z�  �^��K�~6k*�.�� �W�w��k���*z�XD��Y��6��*��H��v���$�L��?״8RF��b��p�8(���*��p�Q�m��D-E=���w?��/����X\�7�]k�6{$#"`Nɛm�Jh�{"=ָӯ �Fn�ga��1�6�A�[�𲬚k�ר���-���NP���2)�|������Tjæd7�>u�Z+Qu �2g@ �
c���.W�6X���X��$�,���I�L׀-T�`n�D�2a��T��W�6�Ȃ�֊����}��خcI�=@ք�/86� ؒhO�_���Y�&�u,vr��ں�z�������$%�L2���]���hҕd qE���zz����sU��s"����Q���oɌ���p?�^�
�]�}��/Tj��D���*�s*�}�����{�尿G�@E���#��c�8H����糏����=	Ώȴӓ���1BDH��R���J�8�ڠ�dNK&�7�e�dFn���|M�l��A~`�u���gx>�N2t�vL�`�QU6TK�-��ܯ��cI�FͶA1���9���1��ۅ�s��H��&�>�5�MP=�y��z��`aS>����/���_���Ds�R�{��3�!�\yFU烎)˳
�ܴz�@̃��!�f��NU]*�0�̢���y*�*��u@o7[Y��ȉ�-%�xҎ�W|^���*�3<��h�%���w�>?8��1'j����WP�Ts%m�zA�8��BAa�����+I���0���bvyx��9�.u�,B���a�*߭o9��̻?l³��������%�7��\7\H�֘�nY���M���oΐr<BR<�༱ΐҀ-f�ǋ"�6��iSEx���ڱ!�����ϣ3�꫿�/>�y;�9�F�|2�{/����+e�����?|�u�ŗ_�*���mlc���� ���6���ٴ���˳�K9�xH���<l�ac��bu"��ʱ��ꋯ�6x��\NO�r6A ga��
ؤ�����.�z���[��d�����'8
@f>3��C�t��f������幼~�*l ;y��sn'�� X}}�&� ��w�~G�+ɴ�����0��i��*�`,�VL
���@�a�g��ذ1O¦�|��/~���+��|�a��%�c�Z���Sf�p���W?`p���s<���+y��5�Q{�-0�}k���rvqB��AX=a��C����b���bN S����X��r� \��G����N��kٯ������^����UV
�1Na{u~.��tr{��vgW��Q��(29{p!���T~��Y	���.�B��.@]Z���7 �H�<nId!_�{�d�W�:��
���r'��n���n��g k��1V�w�j ���O��9ǀ�?���@~X������K��?���{�R�*|�K��3��$�~�!�
P	D�ш�B?I
d.Q	ܵF��ء�DF��c�ﶚ��6]���T�DA��z��������r6;g�?�Ғ�܂j�̪��M�HX͋jL:ۄ*�9�ci��JWT���s�$]E�a:�GBā��＃�Si%��1H������� ȡ�zQ,c;��iAE�x�W��m��I_�VP2Ty��{��g�ּ���pbd�@��@�"VR�c� ���nv�anA�ѥϷp �]PZͲ9=�q�/�����7��z$���dO�WK�1��yCP�W;(螠���� 3*`�%�'����}��j#Y���e���a�H�+�(�R��O�Q��mۤ 	�#IAW�$�Y+��\"Hh��o�,,g�5������7�L�UNx?��CSE�̭�`��[�e�g��5��D�� 0��x�̜����V	�@�r����={"T�'e͜���� �g<?׼��r�r5�H� ��<ƺ�{U^$*{A惨��4�xD����qXok�8:���BAu6B/�7j����=?[m�Ժr�Mz�4�.n�VH���tF�f���R[nɎҬ�R<�|������5�S���F�}k�*�9�:^����B�V��A�Y��O���ލ�g�LDI�p��0�zq,��t�d1,z�L����~�x��(1�LXTQ�Ks�	�'�qD�܍[��`�	 ��+����oW��і�[��3��]__���ź�cX'aAy�-�u( �k�0dNuB���-x��y����܆��,6��O�?�/��%#8w��LDk�����O�ϩ�(���:�73*4[���a,� �q����t=hx}&Sl [�Ҧ ��wc��;�`ɕ�+�����*�Uq_[�g)�cZ�~l�a�ϔ��$F"f�*�u��2Um�9Y'��)�'�%UH̝	c/OT�������D�1�M&��#�	E`�"�d�uA	��KH�І�%��?|�ӌϦ���X+Ú������@5��
�%��:�1�B!��3%q�d�O��~�b	U�0��x>�-��s�>4�V�Y��\�~Ă䓅g��ݞ��E�?��Q~���O�}"/>��$\�a�݃G���5d�s�$�>ff1�� ��p}�}���m��Yj����1CGdlc��~�m$@�6���ml�����O�>�wqC 01pü��s�x�(l�3�'B��$% ��&+�:�U�gt����*��Ԍ��g�V�����i7N��aC��� $�6 d_Ѿ�l��v����G���+Y�ћyj�� :�n�t	瀣An	�� "��|O`�;Ȝ���ɉ|��grv����۰y�����LG����j��I�5'X��Շ+�iQ���� �M�CPް3�?~�{�hXǠFj���,lja��ٮiS~29��٨�f���U��SEB+�&�klI��:=9�:�����ͭ����sPIz��O_���3V?�F�����L�1�*�&uH�D���l������{
��,,0�Z _ل��fV�k��^�TqHj����M��4V��Vi��:2+�hA�a����@�B�Ҟ�}������	2/�LZ����c�,[aU�mӇ���g����@�?����$���lww��ji�jG�Am�:�j?ea̭�� �p���&V� ������9\�����Ƿ���/W:.���t��&�>9`W(�}W�r�	��;�yf���;9�O�R�4w���-x:u�%|X�MbH2���Vix<���c$�]e�kO':�����b��P~.+�#�R�o�O��yd>�~��3#��f�c(��ah�@��Ǭ���W \�4�A������nh�v1}?���Ok^n#��f�}n$7�20EM���8W���x���!��섨i��N��rD��X2~OI�U���	d@�_Wf�C� �&��?̯�ݚ��zW �8���ui��F���GὪ$H�<o� 4�<%	�
Y��}��`�?��_bp{�V�$A:% ��$�*- �� {q?ZN��u�m�����ﯨ��h^���]Y��	��3*!\)7��q�Z,���)	:�X�c���q���q� ��r��)� �9��r�#���h.�!�/�[����K5��3_:{A؋��j4�'�пF&�T����>��yD�<D-چ�f���n��c����n?�������nno�ނ�X�A��;�}��:`ǔk����hbͣJ�����`R�{%����j���ơh��9�t�s�?�1Q���V�*��n�s�5]��^�$1�S��Q���QZ��p �@Z��g��\>y�k�Y>������pT���ss.8�J;9ft���3���3U��r����`�^�D)�B�z����Ovw+�nֶN�:��}bZ�p��̺�Z����u��jCZrކ����$��z�2�%,f22��|:P�5�IX'�*t�ؠR.�1���ylZ��1�/�s���p�QjGݴ@��M4K�R�g|�����o巿�m��"�|ER��g�`}"N`�x8nw�{g�S>w�Y�o���:�aN�;.�V%p�6���ml?�6 c���6�?����[���_������R�+ְ���^d��Jݡ*o6�KVYna�C���Ü�_96֕˨�%(����bU���#\;��zCP��*�'.b�:�T�$�ʠ�i��V=@H@c 3Z�:q�G˦��Z�>z(��\�.��l%�.7���r*���x�#��S�>��m�Ç���[���5� �@i�*γ�s/��7���k��l���Hf��N��F:A���K�pG�%Ν�6��sn�aS���v���9*i2�J��=LB?���Y  L��;�����z^��e���G��O�ȗ����	��������B?�r� i{��ƀē�%-�p\��I���u�:miI����8g��@�k��`�-� �?HB�O'� �����	�E�#�Bo�HO�>�u
е�ڨJ%δ
��{���2�qTx�� +��\b��������4��	Z��׾�`[�k�sI^�>g��M�ّ���V_��-�6��jA��Á��ޏ�qT�
&�3j��F���nG�ƁT�A�˛!�����0�U�k��,���*N��d�e�~F�Z�;�>\7�KP�xE6�Ŧz|�&t͌�#v@&F:�XQ��p�{�%����㯦*��h8X�a��=(h�8�äy�7� �Їm����1Q[5�æ�i�VxhXKu/��6kvVP��&Q"[��	,��0&K!���(�����o����n�5��W�w=�>��)S����Z���@2*	�Yj�Yq��j��cM�^$Jڶ���6-$-�}L�*&��=�u����x�8�l�!/�pM#���ji�"Z�]��������-�-��_B�G5Ȕ�,
%�����DL]������50��I)��_�!��������0��R-z������8�L�RAc#�j�єA8sp0-���Z��,��?OMoK�$h��F�5�(�ҭ���P��k�/��U���*�Tcᵮj�T�WI�a��������"�c�,s#~��:�#\ ��=s����QI��Q�w�x����Y�XkU��ѱ����)M����'��%"i��YH�.��6��7XL��܆������l<��wK/��I57�:���x�³̱�:D�U����Df�A(�$��?{��z۸�g�;4T�q�_����`��g��޿9/�j2+>�$-s;��ϳ_p?�`AIo�<�ˌ�JJ�j^[���2�l��r�&z�_�o���C��Ya�8�|1S�q���2�Z`�{}j�E``q�IJb�I4Ik�zBI�}]q��h�WP��o��V�Te'���_ɓgϔ��b��]����J��nn>���~+�¾9{��s;�ɐ+����c�����g�|������7I���*_�6���ml?�6 c���6�?y{���w���b~Bp��ak��[��ׯ��`-f:�U��� i�,�}�xc���+n�?|$�~����~B����6RV�OӉٺ80`��a�M06��� �,
�1�Eh3�J�kY��V���a_�qs�?<  hUd��F�]M0'1�3�73@��O�M�c9?Y�l�w�b`��1�����ÀuL�6�Ծ~�A~������@����x!��q�\q�.l��>\�� N�,Pq�%��0�,��k��^���|���	��n#�ݖ�K��N�9V`P�'�Pp�`
�#��$ο�IA����sVo���'�88�9B䏙f���?{�D?z�0�7�~�5�y��}�b6'�p	� �h����� ��Q%�j|X5HG+�D� 
�O�����$#���4;=#"��,V�jX���/��
�8`���X���
 �b���ZΊE�/�j�����=�+��g޴_-H�ݫ�[�=Ԇ���m�O\[�(8���Y3�@��S��D�O���y�2��%�߫U���vB9�k�Q�2}�,��<��f�D�׈�U5�Wq�:�'I"Xש�F; a[ebU�p��Ic���6��wQaAۯ���V-'�XH�Sr"�yf��>;5,9Q�ۭ�P��a6J�յ5A�2V��(���<r)�*�Pp�e�*������,�AH�|0����yP;-}0�&�^�Bˮۄ9��`w��A�� bH~�y����X���}>���m�@t�H��4;n�eZ0�3nn?����k����!� |��'C �b�Eهx�����@��a��҃��T���S�.UN��� �Z�G���P+�4�%F�}vP�=��q�9��µ�
����\��:O:V�{���#~ܮ���S#����$ ��]N܆O �� �e�0����,󲢿��a���������^0��1����� ��(���J�'	�W0���#I�
!�ƨ+dN���}�'��>�hHb������r�l]_���(��wq�5¤�_��NFRR�c�T�?�@ �,U��>Ei��9'?#�]m�v} *��u�o�о��O���\k݇�w|���������w�oM�k}g6x5����^�2A�>/4|�"��S$z��� !�a*:�bYn������TsT����_5�>��,?$��\O�O(������	���k���2q{�����E
��_���P�uw5�V�5}�P;����9ù�9w�T��&�/�D�V�c}��$<�d��rҖ�)�FT-�0y#~l��|�=���$5��x��y�1��wߑ�FQ�_l�h�٘���r9�"d�}�����7T1��w��M���;,��矾X����ݭ�I�elc�����m#2���mlc��h,�J^��_��'$2R������o�Q��@"��Q9 �A�K �߿���f���C����ki���fu}�!l�wj���T�r��rU��d������ثc��p�б!y}�p���,��4ʥ�+ ��me����VTh A��i�Y�<���ĉn\�<zH�YP9����� "p^ �w;��h:�������-���)|��!�(Pn���@����)���:U� `��$���D-GP�@��,�����.���6��P��,�Ѡg慴tק��p�l�ި�w�X���=|� ���׷���e��8)`CvvN�ɓ�쎪>f\ЊcN��í�o��'�q}A�8X�
H\K�d���l��Uش���`C�
gs# [ѣ^��*)�p^����K��MA�.-Y��*Ţ��c���A���=�3<��	���� ���!h\�(Y�mć�P t��J��õ�N+^; +���ȱ$ ���;��03��u0o�@r��(^�*�%-scmvl�Y��{��uu�[�0�4U�.�\�5� ���������O:�,�� bf�{�z28?.ە�VH+��D`�}�5|]��K�(�P=۶�D�ڢ��Ĝ�����	��2���V��"f�4Z��@��P��s8�Z�H8Fr-�{�A�J�Lb�UupMp9�$��11�� Y'�����Ā����}�Re�J�̂���	H�J���$H��� k��B��rҩ�5Q�g���`�* ����4 4�9U=T9$ �J�Ԭ�8��jLap�h���  k'��Q��ú�I�Ҳ h�Īr��S�ᆅ״�k9^ʶ�N붪{�n��'1TM��1:�O~(�bV`�0�����?&L��j�����P�椂�?>�˘��������ݢ*�\r#+L���3#<���u+�bf�c���i��Ǧ���b����>c�Q������ �����<��xP"S������K�]Kx�c8	�#�̡���0dh��뤆��{R��I�/?�d�������]�t-(�4��qX�}�u"��^^����$<v�q�x{#A3UY�#C<�Bځ�Z$z��<�<�ic=�1�7��җ�X��z�[�s`٘:r��/���&s�h&��ܙ2k+ܻ�t��l-3��B�V�$Y4�<� �b��ޚ�B�4S�|�6t]����4���9��s�p��ZY�r����v<���>�V����6�<�pY�q����꘡�ψ�g����Ӊ�����ЋE�p� m[UR�5V��B<�ȄE:��t{M�J��aG�g�r?�qw�7��ɻ���͛7�����\<x��<�׷T8��Q�����L5<O�󠢂���}��x�����o6�w��_����'���6���l�H��mlc���������޽z-�6S���߇���U_���[٭�$�������?1�dT�as
K�W?~'w���ݵ,gs��XU6�i=��J����ˬ��v}'���ӳSV�tlT��xc��*lxa	4�̸�].�߮UA���ڂ���y?��v��S P�� �����҃(@u�fS� �͇[y��� @zlp��/�b�&�(޾}'w���V�P���) T����p��b�5@ ��f+�7w��z��	�ǆ�h��"�x�y��E�j��~�䗗yn p޼~-��a�ܔ[ ���G�0��|>�C��"�`T���39�6^�a�knpA y�vg 4�|��Ϸ�u+��Uݴ�p d�)�{ �������`^� Q %^�VEdS͒H�+|g�V��˓�,D*�
2PA+�k�k���=Ē�`�l5}v��yϺ�*�¬SҘ�Ąz��xM�06�����޲#&60�=j��UjG���w�OgyT�1�� � ��n����O"�O}T$XF��Q�R&��/��P��Pb�.%-~=Y}�J�(�N�~'�O�.yE9m9��Y��xϵ�z��h�!����O�����&F�����:\�ih	�ۍ���d���@��u˱��UWLD呁OCO�{-
���lbP��,�ڊ�lP���dV	�@�V3#��z��=1a�`����$���4;�>���8A�e�P5�1��/��I��P���]X�}�8@�i���E������R��
�����F��8���@�$��_u����3CZ�xn�҆ʛh6$,D�ʵ"�
������#��1�}���������� 9ؚ�s�b�"��t��Y���kݏ?_���:FkS����eN״ �N%T�E"H�������M��?�9�G��\
(4�Z�<_�8��T�� ���t�.&g���!<��o�:��5U����sZ���H�a�~�����2@������^Z���|��3��6U� ����j�}	��>�V�]��LTa�6\��I�����B�Ӛe
�&�kSnYNY��ˇ��J,�~Yj�
�FE�%�縜�	x��pqa�
�5�>��%d���6�C*�I���ú���%�\l�B��䇫B���b�NuHҏi_���`��k�߷�<�5G��P��|=FX��&����s�+I���+h�l���g 2������)�{�><WLgs%;���M��T-�~w;�jʟ�Ъ�S�E-��v�, 9P��g�ޭ��~��ρ(��g�����v^�V�g�0K�~whA�ͺ|2�#�?�?�)�������/��h5���ml?�6 c���6�?}ێ�qG��j��"�����_���[�8��n�fh}sM`&���=6�R�Jᦶ.�r����odss����ͭTa�<T�a�(�E}��.��Z\h�6���&{�hm�c��IC�Zc�_\��Վբ�Ŝ���>���S�ڣ�>ʨ*���a��[��S[-fji��1|����^^��������r������咊��O�Ծz��߁F�L��*Y��v�,�*_Z(����� �S(vaS�e��1�?�G�.I~ ��]��P�n`u�UO�����g��#�O����~̰����a��T.N���H�<~,�=�\��l�b�`�GYk�*��G��
���� ��	�
 @����`��z}9��0G.R#��W�/}`���=;��*�Պ��V?����?,4H~J��V-� ^ �Jn@]�E���xM�z�y�l��7�+ �*?C�<���� dh �*�uh(އ���@)@q��/C[1� ��1��B��_@Z�TK�*����N����0>��6⤃j𡍖 A��}'s�@~��W�z��jv{/C���+#Ok����S���-�Ї���%�x��z+����ژ$���ˬz��  ��I������o�>�F���:��M����}{%�j���`=���G�%R�[�����A���aU���̰���r�k��2l\���{�;�,m�1�@/@�tׇ���l��y:�y3"�/�]##Z#y��R�d�1�<id�$�Q���6}$
@�T�=�ͫ�1�}��dx0*λ��l�9��������a?�|�>\�!I��x�P�dI(U7�vu@�k�+9H��eT͸����m��������2�O�'���������o���؝(6Z=b͂J¾��Ɂ�e��"@xΚ��I�dn�^�}�`<�1�	���£���<Jc^Mj�="EFk�����9V0N��WE��%��K�VJ@��������>ue��'��@�r~}�X�>��I�����	�m״ͦ!a�� �'����x�.Πp#�*��S�����.�بT-<פY$śJ�f�^s�F� �!�R-fT܀��
�OP��%�|@E3�eTG�}��.����:�)��&�����eTj��U�(���Z�IOQI,݀�%=ޚ�^Ii�^U��k,�E��*����i%7��sn��y��f�-Λ
=\���SnY�y�����H��D:Tc$t���*=R���P�$�*D힎u�@\+P�P�N��<|�X.�8gɛ7��ݛ���íd��d�q"\��e��AU�c�߃>Ü��Wo��mx�jR����6���l�H��mlc���� }�������<m�ru{��rTkf3*&�y��Y�,�k�)�/3�) c,�%��/x���U�e�өվ�-ճM� �ہ�+��a��+*$�����>����U���UR���h�,��	����W��ކL�{6�[y��e8��	�#�5	 �y��5�|��>�!î�y��{��<�	��_����X�T�Nt0��A�U� ����A��#I� fg��#ɍ:|ǧ���S�>\���+Ay�F�/A���kQ9�Z.��Ç���*lb��B&�γD.�O���L��T��X����k� �~��9}�?��PA `��p�AG�%��ꅭ�Ձ�۰ނR����
%�H��-h	�Aͳw��@4���*���>d@%a`�E��'i�}Ő�Jں�}��Pؗ�i��J¬�C�V�pa �<<������mT�/��\G*�&�$Z�ٰj�A׶u�U����1��Mm@L��A\���b(�Ttl����c�<�,��9��1�P�LXb�ﾃ���ǘ�g�.LԷr��:	� �DO��s�O+����C�92�{��{8�O��;�q`���Y6�@c+����y��a?ϣ�#8������Y�*n� �*V����X0[k����H |m��م����N�C�� o֓$N*��O �2U`|M�R��!
�*������wJ=�����iX�>�V���k��{��$��>��!�w�q̠��D�{h���A��*�a�U�S�� �B
6:i���}�19�!ؘ�jWs��0�_�c��HB`�W�Uɀ$��s6���l����O�����FЪ��Z�V�B+�Sa�b]�ܘ�=��Z�c�׷v`u��"�'JUզSt�*�1S&vr�I��,�{a��i�ǩ��v,x���GdD`P ���o��H���#^��?/�Y�y����sb�5���g#�ˣ��J͢�����TnV�C�[,dB�5��"*�|��H���>��N������'F��<��
�V
{�;i�$i*- ��QA��:\[�<��9��d	<�e-���I��?�3fF�U|��9��Y�N��PdS-�@�G�EP� �����,����܆��T��sƜ�4��H��[�.Т��R��a�gg�.�T�x��]sY����IT���?��g�)�R#�r��hv
I� �s�E�b�U��{���E>'q}��:Z4�<�xM4k*��k�_�����c�g~&�C���U��M�g!�٩|��W����ryyIK����o�폲��H������� ��-�U>cT���5��t6�~z�}x|K5�glc�����n#2���mlc��jӉmz�o�[�;�/�/�W����p�b�K�t�d��D����Tum��2zl�
�FǦq>_<�������(h���,�ONV�ֽ~�N֛���F�Z�簭9��>|Ɠ������6�7>��wWa���Ńsn4Z�{�V޾y/�q/]ؼ�/�ev�T`&ܶ�
��aC�0�Y*��|��_�y�,|>�f �h�Œbl��=�wU�r, '9RLÿ�e�JU��M �*����I8�S��cs
���۷���X�i��m����Z������������W/��a:�$`�<9��G��g���g�iY���k���O���?��K�I������$���I$Q����>�qc|\�|�|2����sZ�Vrvz�M>@u�y��� 4����` ��oՠ������bn���
�Z��54/�̗g���j�2�g��MI�mf��玊b*E�x��&���Y�G�\����>���p��nȘ�烄��y�RE�6��T!�t�σjJ���;nN�x��U�k��?jS�+��ϟE�`>H|��Q��*�M���T���gG�u�5e�����Vi@�W�sy��p%���1j�v�y�� 2X��p�̏A%=�f]jD��v�TtMB%PU6\`]�v,w�7z��3��Vh��z 2�Vm���tA4�1x�S�fG�Ng����j�����Jtb�s�$��Y�89h���`õ��|�+����Z�(��Qu��`,�:xe��x���R%� 8�$T���8��We8�0���8KfH��I�#�^�B��*Z���B��:%'")��X"[%p�k�� y�a��>qLU�B� [�+��OG �9��v�������}���v$'�p�	N#d<+h����R+��2���#�����XU��չb��d�+�%��	��й�\,LQfya����5JZN"x���'S�s�@�bl�ߝh���R��Eu>[��r�Ľ 5?_3U��C�ZX9�i$*�e�̊4�ED�=��?��q�TH l��C$��30)�x?H�Op/��~%4��BQn��c{���]�;Z9	��`8��Ґr}�A����52K:�l1T�,�0�G�Re�Լw�:0��4�4��N����nsT	d�*�S���>\��p'E�  @
�'("�^iҁ��@������m۫��t�9�r,r9��AŋuT	�s�	sm����³Uy(�w��S��d��s�f�m��Qpqs-�p�rF�"�m����U:�Miק��1+��c���?g����9Cy�en��M��J4�T{�\�����HC�نgަk"���+�ߣj+�	��c%<|�������<I�AA��Ǆ�'�N�ڴ阍%�+%�m���ְ��R�8#D�4�M9���5K���tI�!�i�Ǚ�T�!�.<��?x ���Ky��Ixv�D��B��?���_������Qx^�~ yx�yEIx^}�kG����L)�p��z@�����~)c���6��w	���mlc۟��X�h�����ڴ@������ �a����� �1�H(/aC�R}T��,����Z}ܪ����ҕ�}�	B�Չ� -ZNh%ކ��<z�� P=������0ps��Hha��Y '9;��n�l:Yp��J�L��`㿹�������jC�V) �]^���` (��/}�Snd����ܵ������o�Z�U�`��p=N���'rqqN����F��?p	�7�+-�grq~.gg�vy������� |z���|�"lj�=�,l�˰�]onB�nH�����\�A	 ��  ��](����Y�H�l�US���:|gC ����7��WL�s��1�h��b���u�y t��'������
cІ^C�$SUHb^�����+��ڶ��VpE�`�-���X(h�� Y�s�KV���ډ��+�rI��bf��x:��4 G@T\���1�1:Gp�`>\��du��nO,g�+�Ӽ�l��w��݂dh�䀞��ǐm�HlDz�T�ώ�W��Ej`��!Y�7�?3 ���Xi���<Z1���q��lI��*�@s~_�@�
�k�c'g����E5���7jF\��m`���x6p�	�̑X���L�(���|���j)�}��F+������W[V�����ȋ���-��k���^���it ��n�$�q ��"ޛ�먽2if��Q;��c׉'����1����`)�?�ٓ"z�R��-oțr'*�J�F�ՊJ��T7;�x��������k�o�W��yx���G�h��J�,Ԯfx��F���2$��,��N")���>p��*~'/�t)��*��q�^����@^�RWQ��뗾.��ޏ�8UG�?p���hشY9�*���u���y�/dB��vv�j�x�3@I��R�m�=g�Y\���sR��rm�c�u1C�	
\���;	8g8����`l�>�Y%��[6 :jS�J���rzO�k�ݿ�Y�5��y��,r�4�
�2�
�D�X�{bKs;�@ú���@��ք�sLk��~��F���>����-B��+��Tʏ|��.|/���,iň���w�W�9疟�;f��zVyƏ忄5`�Oh�
	�Q�v��w%�u��8Ԟ�S���µ��F�Z��%��W�tRUH*����Cg�[X_2vՔu�X�k� G�h-�,�cDן�>�]9�~�Z���Ń6S̊��z%Z�s,C_�L��s�y�_�A�]J[�rZ�*�yT.�����p���_��$$̶@��o�=j6�|)�J�k����n+{7Xk&Pݯ�6�����m$@�6���ml��������n���D5ؾk�"灖=�V�b#�
������r{�M6N'���n �8���{\l��&~۰�"��d��{TAu!��a3Ҁ�H���v�ћ8+f��¾`�&*��$�f���,�MF;��WW�.+����S��\�F��(Q��F6�=-�޾şa#�������N
�8�p�����
�׊k���ѝЏ��ƪ�*,������Z:z���vB��y���<�|ȍgy}����K�y��l��O�+C�� ���N�u��`�G����;�m�����G��)O�<�Y���fC�
6����i��^����!�P�yT@1_������	 .�*K��H9&P��kP��AH���ܘ��pd������q� ��D��p�1��b��Z�yb��$Wbd��$c-�U�@d��������2�����[ɠ9�� g"F����\p�~ ��Q���#��������J�۝�l-" �d��p  ?����퀦+Dؿm�=T�H���k��� �x��G�'|��ѻ_$Z��`x��%*�S�
�ME���df$�XݚF�~臟��f݃�$�`�d�C�$��} 5���>��N9���I���9�����h�?��UE�*��D&�D,�0W�N"�[���f���n��	N2W?V���m����!9
uC7$�
%W����d�fw�09A�%�.���g���Qa��=�������^��6=~�����Ș�G�tH���1+(��BIG�X�y�����G�,�����uR��h���
J�pLj�x�㚤�q�< �#��� )3����O��J��}�cܕ��˕8�s�8?A�;����:�^~-꺹���yU}���m��-��䨇>;�9������ӵ&3��IP�3� =y��̓���_�*y�#�X���f����Q�`��R��2�HER�r|�| ]S�Xp?X��G��4�k��_���=S�vJ�K���b�Tҫ���us[�N"���w������[Q	r�,
�[&�'$�2�h#��ɬ�9a��ޮ�{H��M�;�kJ5�W��?�9�)�M*�����q���&�~�x�;���ժv� �:�fx��]�����u�l�k4lޚ����`����A�5-([f�	5�LUI1���6("4ˤU+,���:��Px��/A��_I��x��Tb�c=Ǣ���P)u��+����0���ǹEEX���h���[k��D�7�6;H�7�*)Il��2yj�J/q��d/� q=�j[dƽϜ�~��d��ř|������f#_���k���4|��-,W�p	r�P;���K�����{���6�����H��mlc�����ݨ�2��`�^��ۮR�= Pk5hZd�17BAmҰ��Փ��%��Tԥ[�*�}%J
Z�t���,cd��3�=��> �w�.��F�B>�FṕT�b�� 󻻍\ݮ���ۀϫ��p|��k��_Ȼp,���VU�@�af솘�6P}<y��ۄc A�}8>(# ������k%h�YF�@��ac��:|/6���Kd����Z��]��ys�9�U9��i����L�=*��+u���W句I>l��Ky�����S�|��$�zs+]� ��/rq�X^�y���Y��3� : ",B�!��;*T�s_�94P���UC�\�����?���ji�F��͕W��s6S`	@|Q�*C=�1���|�[�iP�`E׵1��Y�bZr�*M�=��8�	@X���6m�P��̻oTY�eK��q��|��������:̆p@�mXbظ!- �]���T�uwK?V�������s5����x�wys%��棇';qr��nf�
&7F�$Vuݓ>y|?_;P�h.���|�߽hqbp6�Jԝ��
�0��`���+����r^��J�Ac��<�?�s�\ �������
�k>��l���j�	�AV�"�xP$����6G�����= ������<U܁��!�<��ʧ���k��󒀵D�,�T#�@d*}��ޘ�sg��e����y��1�"z^=�����Z���U�B�s???���ʴ����*�1��d"�W��(�g�`�v%@Ӵq��y2�v��vB lq�J��b�;���zs�ua8?u��T#	  ���w����C�q����[�V���듫>�:�>$��:�"Y�s��A�TZ�gW���Z�\(㚑��������a�T{�r0��|��2����x���ʏ���w�g6��e�0u�CXF]IF�}��*�r]#�N���>�{�c$:M�̒dC$����&m�h5g�W��N<y�ɬ��v��nny_��
��`]�+ٮ��:�1����	E'�c�b�j��Y�CӫA4O��$�Y�eD`�8�ϙ#��:��A>���"�3i�iP�%��^�y���(���gE����)-ߎ�q���\h�|h��/��0�2yO����cۘ�c�R��g'��I�s�}�k�ۂ�\��ni����^���H�Ǯe8ᙺi͊Q�"����ɥήS�6�������F4�[trӤ��s��yɎ;+DOU3��i�g� ܽj��۷�/��/��(�V�E*��"<[�-���_� �p�$���
�A��v����h��`�tF��W��mlc��~~m$@�6���ml6����z:�Hr�x�= �\sp�@��-��hz[%��}���]g�������{�TC�m��:Z��X%�*���s�ַ�s �T�`�	?�.�]�Y`nm`�t:���IZ �@%\G��p�G�h=��<8;'x����V�^_�ʇ�[C��N���Y-O	6�[����cUj�q��� �a��~���n@'Y��am�5�	s�ʔ�K9Y��csy��p:_�+z�<�{4`٭_��@�/�B�<����Z�o��v��y%E6����|��_�_��i灰�J���BX���C�+-ʃL�7��
��Z�/OV���nx�x��]5n�!�L���A��zc�]��ʇU� �p�Ń�I5�z�$��E�`�N AX1���� >"%(Ԕ�T)��F���.J��6P8�h8e���fk�U�� �c8������-�{p.n)�>�'�����匫�X�:�����4^W���\�n��9(��w��U! =�`��p0�}T�2��p�M<~f�4=`��IO2�gE_~ m�j�X�j�����m�@]�[F{D��i�<���1=p���Zǉ�Cs���1R�>TK4��ju�P���Uǒ���1k��e��*.�a�C|�]�O��¸އ�GJ����@
�-\�0~�T�P- ޮ+�����/���1y��ڶ��� ��gR]T5��0�Ѡ|;��dr�ىK~�j��h�nx�t|�௓_� |*��`�8X�q��&��ݷ����)����v�9����v^a��C��r�P�jHc�j��9���"��������X�O�AJ��έm{�ox~�n�5$~} 	�xK�x�a��ݐ��x=�yH[{��ىfèa��xt�ϕj�3'�H������{���5�j�p�΋��zmD��%z|� 3���N�Ը��**�8��~�v�c�P �1���9R൭�ط�f����T<7���3#z�p�����WUx�B�ES�U�,ZVJ�m_N�:��}BU�կmGi�s�W�T�J*�t,�%s?L�ǀg$����E�y�$���[�i^
Ɂ��'�������P��B�	�ՂV��n9�lRP��9����}�Nj,/�m�d������zcvm����TJ2�'��Q�x��Ir�6��%����̉��2׈�$U�U'$U<�u�uJm��yX��8��_]�[zʹ�9Y����)��Z�j-����������6ĳG�l�TI#ѐ���k�kM�X�$�"V��trx]CU$׆ԕ�)��΋Ōq����R���w����*�_���x�����c��Sx^\�?��_�_�;y��'�7�Ֆ�f}ᙫ�T=H�)Q�FI��0���mlc�9�� ���6���Y����{*	҂p�ps7E�O�Q��M["���p��v4J dfo�a��N�n ���1l�*#�t(>��ؐ�v\�R7����$R2:ɥ�^�l8�hPAk^ŉ�wZ-�
T��&�cN��������Ѧ��n+�wkV�m��L@����%7~��x��xi6����*zъǆߟ��Uu���a3�R�Ѳ�߁�v��s�y��U���1�6�Q{Дʆp�.=`f���^�(�_�D@y��g����/�����?ȏ?� ��B�^>a�*v��d� 0�.�ͧ��g�,a����;y��U �)��a��v�� �L��<��#�H�mSR�S����o�  �Pr�8�V|� ��CH�oc��ف?u<�}W ��5CG&7�E��F YfFB��eU*��H�+*�� &M��>���c�>L���R�F��F3�X��a�K���6��E���JP5��Es9xN�� A��LL�0l�0����;����;��:4x�{�vfD�[�8��A��=k5z�l�$�@�����|d���9�"+��Dݎ��A��bN���2ԃ��4��~��C�_OP�n�\���W۱��p��w�����ޗ�Uxe�^#�n>�@Vᵮ���]��8�O�}c��!�U�8$�t��x� q�^��»b�:��dG�y��>���"�z�b�Iғ\�����@@���&*����}E3|2�3��*-0Ǉk���A� -C��9U����1��Sp�_l�R��rBj*)�<����T��c��2�V��,�$e����h�SUn�TF��?�#)�-}%�����)^�:����+|����94$N���)~����!	�v�ݕ��XF��T�@�`*0?'�H���XjV���<qbת'��~Tk��WCh~��	1��9��l�pR7��N���И�6�����{���$)��,<�L6�ܯ�6�Q�dN��c~T����}�g�D�ʬ���>�9���0ų��SZ��P��v���hvb�3�տA�LN�R���
c��
^a��oj��q<PGi�Z�0�JzeN�h�=ޏ��?z�q���AEˮ��S������O��P �+����]Y�s�Y���7��*r�#�����F�ڼ�����ڭ���CQ�6��a]��W���z�����y����ǝ�9��� %0�@d$�D5���H��'�
8�|���3I���6�4[
�Xi�eq�g�W�<
Ɠ���C\y�ו�W������Z��>j��n���_��?�O����م<~�,���ܠ�f��9��S�,Q�!$�'��Oc���6��c	���mlc۟M "��1��N�F.�9�!��̏Lr��j�n��?�(���'���Ԝ���V��~�6�Z�[�j
�	����6� �[j<�z;�}i��?����Vn#;D�BIK(X��ɄU���)P+������I]vS���-�y_lX���i	��f7����s�T�SU�i(�i;��g 9�VG=x�H�<y �Yo���U�8.5�7U���!l6g?�~��1A�wWo����Tx`S������˗_|!�g'}���T�F�gn�a��-��A����=�g����u��BN��r�:���-���CI��<�P���H�?� �U;��9#�&/�:ʝ��^����ՕPcj(�b��I��Ҝ�GV9<e]6ǃ[� �oP�	��~j0���ؔ�f�$V%K�Zh�q�P���AR����Y9��1^��w��U��pk��4U$=<Lى�<?F+&�Tz�@�F�[�I�Y��;��O�(z�]`���t_��"mH���=�^1ӫN�!�~����a���>8Ṕ���p��먼�n3TBo�[�f��윕��cm�h= ���]s�o��J�p$P�:��O��$�b �jp=kˎ���������fn�T����>r�p|9� ���z�[N�)#`��<��FÆ�V�E�I���(p+��L�m���� ��z��Gܮ��jr� �K�����y�3�\UY����[�!���%Q��j8/-�BL�z
t]��#�o���3�ʄ׏�R8����{֘����?����n�&J������a��A��N\�r�J�.��&�`mM�p�A��Y�ϊ���0TZ��焦[�8��a�����o��j�e�,�ǐj>Ǫ�`/Ǻb$�=�GCUh�?�q&������{5��Y���[#�~�wK�,����%�s����fY1]o�
�Ĉ���[�Wr�:ǝ��~����1T�it݇�c�ף�hdWAɆ�5c�L��(Н�����Ts�f���=�1b��\sr�Ǌ*�t�v-*�*;�z_�2K��mx�i���A2�EW�zo�pm����٧$�2l�4��R��y����㎄�6�)_�+Z����<���
�c W؞s���VM"�劶X Vn�ne����k�����U\qͧ$4JfK�$\a�%uξ�3X����b��U���yLM}��ǚ���I<�N��#Zdp�׾�k��� ��r|.����Z�uf��5=�D���k�����Ϝ,T�]��Gs�:Sݚ�����LǗ�� �����.��W�ý���ɉ�s��ry��jk�C���O�$�޽	υG�����	�W�����(�ilc����3n#2���mlc��7��.��r}��X�	P��P%̱���y�PP(��Ѩ
�Th�U���@`�C�\=�Q����<���-�R7���[��p#�z���,S����$���������� Z��~� ��2�/Y�E��?j�� L oI�Vl���Jvἶȩ8������CN��͚��P�欴��
B��m1Y�:6�׍U.�AUC_��/����驜��NC��k�@~�3K��|Fp�����<y�X<x���o�����ÿ�d�p�I�ә|��_�_��Wa�zI�V77�{rvvF`A� !���kv��i�6P�l�1�g����ў��˗���k^Tp�\S8P0�T�"���x���(S���\r>f4hh��U?_�`���3��7qb$U`����Z����I�d��uV>!8���3�@��F�UҎ����[���$S[�5
 M�Xv�`�C)���G�Jg��~ր�,��+$�J�{��a�bV<��o\�Ѵ����"�.�Jc��5�
�g���SQ��z�w�YM�c5��g> ��Ӄ`��|�rq�~�L���Y-_r|�&y�
��G��3�6k��*�pN�+nӄy�����$�{�4_'�|� h��C7�AJ j���3P����+�)�| s�D�7恲�$s@�f6�|,Tnj��^�Z8���x��a#H9=9���ұ�9r�03�5�_���u��~��[��8W�S� o�,�8i�@ά��� 0*���2��jQ��W��b�Δ>�v���}X�t^i_hH�m��]���f5�$���,`|��D^���=�d;umo�� ��A��if�fg*��#�`����!�q}�L{�ǜq?c&�����^s��#�����E�hp^�����Ҩv�s�c;���>���sE-�ڸFq�A�(���C�̕8�j�9,�^��3K�f'jg��/��}��{E�g�*��:���p����=�UR���{��D-��{Q�n��f8�|	3��_�>�b�@�����v�6KT��JFFrb�h�HyΉ�J�ӌ��P}���ekf]h$m��ς�\�>|[���l�k|���-m|]QT��ɐ��jJ�̀A(|y Q��u��>��G��9<��5-�T�h�d��U[13�QR��
p]����й�����I"w"�h��=S�bภ��s��3؎��˹��gX������Λ0��/�X��hj��f^����@�Jd�烖�\�G�#�穊��4����3~ϙ�3�I���	�W�,x��-�,�(�@q���(�t���#�$�[8&�4���2Ukg��a�	C� -�Ϣzw�VbF
ߟA�{)-�Ԗ
w+W��^��D��QH�\�d�.�Տ?���F>}��d�<<c�K������F�N����?��t�gO�{݁*�!���.:���mlc���� ���6����ۓ'ruu'��:??���A��\Ζ2͖ܘ�'S�8{ �|�M,�2Z���: &&�o�Gx`dm_�&
� :QŬvj����<WO�)�Vַw$���y΍֣Gh�Pͧ�`E��l	&�&+�>�~���N�7��P��E��P}Y1�75=�Æ�����^��y�`��9B��!��e�����L8Tu�� ���^���$��P?���u%��[���rPR����% ��p^��	l��N�4����r���<�|L ����}'o޽�*��N���_~J۫_}�K���뛯�!x���c�K�_��������*X�Tp@ ��f>d�����O�}UW��$2�AۋL����@n	m/Pmy�B�q}{E�f��﫻Z�N�2b�3��5%��0W�\SrD�q])�����̴Z~���|�7�J����>����O�Á�hk�MLɠ�ܴg�I�P!�Ѫ%��O�h�( Y�� ��y��ڬ�J�L�4���$�~>��kM۬#A����A�G��AmPm�$Yz��!°�K{��IͲ�Z�?�0�c��h� E JnE����Kb`p�s^�E8�41��趲��D��OP�)���o�a��3��pԫ]�����(AT���7�T��"���[�� ��:6WK3��tE%<��n�o�9 �?�\����]Y�
���^��"L����L����$�S��A3���~Ke�tV0/h2)�S;!���@�����<RA5��S��=����Ъb�P+@��	+��d�^$������$��b��$�X�<1(�P�@	��	�dΑ��S$��'>�2�S�쥰n/n�jc(a��S����G D�ng�n�3��J'��(A�L�xY����a)�1ECa�S"�0����SĞLf\���	v�\��+f��[-j2Y��b��T=5a�W��`u��g'a]+t�@E�!U7��/&z��-�T�X�2+���e�&��$'ʊ�WMLO�\@|��o��d��*Ϋ&��RQUB��>��o�C{�����y/�R%7�E~&2G巩Р�D1^������T��Y%����3��A���)u}?Y��� �џ�p?i�}+0>W�2̯DM�ky���a��l���C�:�-�~��`�9�߉Y��$Km�1�i�i-�h�m�߅�T{�֦<ƶ�, �3����2�4�e�0>�#b��v�[s'2k��=��V�ZM5D�{(H�=W�j)Q�5H��YB��ڃ�4��7-�j�t}n[S$�^��]
�4	}��M�@�X N�Ȅ��V]���}9��vw�5y�n<���q]>}ʹ�qy�}v'�T�צ\�cW�q[�z}T�I>ca�4��8���9m�J�=s����f_Up.�@|�n�4�󽼻��YNE��࿛$�3�p���$r��|�����s�h����jjQ���"<G����̞B��1fꧬ@��l�٬��
�ڱUK2�[��K������(�h�I��ތg#���*ԮƐA�Iv���)[2A-�I�>�_���y�vbX�:��_�������|��r�����N��8��|֌�\���ÛWrs����I��ȷ�d)<�{l����6����g�Fdlc����g�,~��� ������5�����P�X� �9	x�0�7���|��[A�B+�Z�&�Z��W��V��.{n�O�6���\�S��gK��4�駗��w/���U8��2t��^N�@%@�V�ǅJUVaKMpn6���RY������ `���T������<�k�Z��<�3��aM�V���G�Y���r~rJ ��斪t(쨎�J������@M���ߓ�3��|,�� b��X�~����p�Zʧ�=�O�=��咖b�߿e�T�zߤY+g'��]%j���հ��l>�����Z��n�Q�jsf�G���槍q��5�u����u"˰Y�E,�*���J�>�j�y�����A� ����J_�o��DB� $Rk*�A���clz��-�?G�����y�gR�7��UE�lw�f���!�%���vIoI3FFzHn�|��߱$�4�@�V�T9)�c�bQ	��Qy�r5�J�?�"�p�?�%�����b�����*s b{8��TbD��/�Y���P�P��ۺ�1 ��-�$�Q9�~� �`���JP�����Z���jƬ� �{P-�"Wz0�=V�K$�������*�]���`#�r�DrO�����S?x��� %$;<���[C4�B+�[S���3ڕpL����z2)b8s)���
�4P��HB���U݅�'{2�Pi%q ��(��x��fp0*�ak�k�'Rt����g�h���d�� �ʣ�u��kzL��w4*@tM5XJ�Y2hP����-,Z5��X/�F��Ӕ�r���Z�u6w��>�OL-���Pn�/f!��Re
4?WX�:��!������
���>na&�V7��� lõ����~�{�����h_"{D	3%�����J}8z?.b>���?w�����Db��U���3̙W�^�{{[��Y]Y&�)9@fLE�¯����<S�[ɜ�·T�%Z#&���:ڸ���R��Y~��+V�C� �L��)*�l�i�A����:g�������׋j$��sE
דĕ��ٗ�{�������x�ŋyT���ˌ#����V�s�q�T�@#���fC�%1��'�\"�����Vǡ����<ñe�_��~��H���on�d��s~K�#�m��U�����3|~՚�$>�����$x�56�ʈ2�Mq���Dpe����q�Юr��h��VĬ�@�g}��d���,$�}^Ĩ*&S-b W��ᑬ�gU�1c#���֯.1����s�~�pl�:��6%a�F�F�P�{1�G�J:7��yu0�x�M��\�&��g�֞Q2o���ɠK��HS?-��}��'锌B�q'�߽��IVs���|�K*���O�7,`�������]�#���"Ѻ{��!�U�s#c���6��o	���mlc۟�������r���L6�m��jขG�V�p�l�"���/26d-=l`c�Ѯb�j^���84}�k�d��*���X��`Rd�}KZ4�gs�x�@���V؆��_����d�jm�^��8����i�@m9��-C��*��i��� (����{f�X�X}��Z��53V���郞�Zv�1�BR�f~I�#�I�W�j���X�s;�`.� 	p1ߔ�Z�	�IKQ�|����۷/	8����+���s��_���	7�o޼���+V��*d�� i�-K��
���LC�u�FNV��ۛ;�p}-H}��UEULKk�f��e7�P�L'��w7������3��mu|8�����y�J�ă_(w���[K5*�-��`p�C_�U�B� �T=@F~��j`rB���hM�vGn���l�
�27"�(��	���9���0/}x �5�"P%Z�;����{_�
ڵ���d:'��.૳����򉝏�T���< U�B�b��?���qPM���sr��f
L�J?��{�+�yP�j�	6̻"�!�Y� �,�?��!�j���*Փ�$�c~��U�nM�9rD���"�?W�A'��9��a��"�?�o �2���c�M{%ɲ#��kx�oɵ*���z%�$Մ4��U�G���r$�"{#�ݵ�����w�s�Gd5G�؍��W��ދ��wq7;fv��Iu2B� ��4�
4"nÓP��Y�U*S��*7�?r�H�al�rp��hQ� _{T#�t)F��֪��K�
ʵO��}�zn ��`Su]m@[Bз�j�>��o��d$m�"#` �M�|�'�_@~��u�=H̫ҕ �I��5Tp#��N�� z'9�r��L����v�f��cn�l����1�Z 9c�## ߉{�3��.����Ȁ�ig�KN���p؛zʃ����Y[��UQR0g)�|����Z�v��N�x@�g�EIP�N�P�sQ��]�;r�<�?��=[����]�Ϝ�b'�: �q��ȱ9�F���I�z�ɮx�Z�t	�����H�K4*��`��s�k�s7 �m�&��f�tb�o{����Û��k_cBV�e������m#-�z�;$Ӱ��ڧ��,(A�^�'�!�:�R�u<� !)�A�acc�UkJ'(L��ӹMd򖌀5U��� !o�@�)}/�����M�A�!��7Yw����l�]٭7����`�����|����z���_�J޽{g�3F*��B8Z���(���$��ٜ�Kd�����ŽAkV����N\�R�B�T�G��/�)���V-F'����+=�+�� {�2����bͽ[0g��#X�Ѻ*�{6���Cx�_d�|��Wh�ٶa}�}�y��j����������ݓ#]����},��a#���ռ7����<���Y����-�d�K���ހ|8(�z��������!�e%?����a����oH�������0�W���6�����Fdlc����Go��؟L~���(�����=� ��_�#���#k�:��V� Ȍ�� f<#�����z/
�'�;�����X�� ,bP��V9{{0Z-�̢ H���r!��Ohw����v#W˫W��?�)�3~��&�@k�dJK�`�C�1 +@_k�%����������a�a�"�c�+�"d�熑����p�^�<������\�^��%ģ�r6��  X�K,g��@��,�\�^G(EG�%�$�.���J���O���?�Ϟ�: ?�x��*��/*o�X�Ss�����͖|�ǹb����	D��x"`�1 �fbD�
`8,��:��'׷���޲��@�g|�+��;ۈ4T�2���0A;7��'���`�K�ЃF����V��8��DN��#�q!��`Pr3�����|h�7�U�@c`ʎ!$�	�#�+��5�%|��k�,V�;��ɹ*����L��{��y����2��; �-��v����cMK8�)T��Y"� 	j��U��L�������G����z��e�TfY�O'�14�2Y.��5ȑ!;A����a�_�p���ZY~@K���?��v��#>T��?���@6�hP��,��'yzA(���Ⱦګ��q5~Mx�=����
�@��8��h�g�K ��&���wB�ƾ�����\iL��<7B&�(��~�r�'6�����U�nD+T�G	�2�o�`3bA����	#��
`6�A��U4f]�TF3�~dj8~�v1U���Z�ޚ�5��ޥ*m=���RDȤ�Hc������}@8����X�q�;O#�`��an�NL鹚�T�dIl!ɞ�A� ��[�$�����tP@`��sK-)>~�Ԡ��s���?��2�@*�����[3��,򺩑r�����{���yU��g����'i����l�:	��RlA�z08\�'`�;˰7�ܤ@���!=��|�<�$v���{	�����������C�P�H�Φ����Uk�c�Z�քa��ϨC&��R�R��,G�T�IN��V��ga�EvP�@چ�
f���u�>	��Y�g�ܦp�z�?�\���춏���?�/��i+��O$W��#�֩���?��~�{�����L]�w�sˊpǍq�ɢ���ƸP!�5G�T�z-�*�Ü,���.bm��p����:��OdR��nW��3'��P,����������Z�� w*w$�!7��M���GT4'f%
�l�������j���R�ݳ1����l�8M�%��꺚c�ͦصl98D�p?��V�4��Hd��>��?��~?��'����K�/R̯��y��9�Q�o���g�l�cMŸ��_���/����6��}w�H��mlc����m�� {\��_~̇`������a��f�f5{d��0G�l n����V�p�%��KSM��	@�A��F 3Qu�:,�S�2V���,�a���(#�^?�믿��[����>�����7�߲�t97&�5s�(E&m���e]��O&ST�M
�E���,T�A��zw�f����Q���}��%�	
Zh��%PEp(a��q�7�h�G.V~5N�4<��{�y� u��~�o�:�d�t.OV�R��z���� �h6�.��ˏ�?��*'Y,��>�n�$P��V�;�����SV� f��l��"�`]\�dB2c�?��>������ �O�r�%��>����x��b�{��a�|䠶�_���8s!�0���Ԇ�' @��?�20��@��Z�S>��G���B�;�Ce��C���1F��q"�n�F��Qמ-�
�+�Q��s=�X�w|�Z?va��X8L(bb���x��<�V�%����O-���@`{� 8��	v8�������2:�¶�5��h���!P�@hj�V�3$�����\�g�,��́Y���E]�' 2�>62�"�W��t�3lvb0�1��8! r������I瓍A돌AݙDG���B��� i�a�B� �C�&=�ү�4���֌�m��E�2�iFE����w�ʰy1�	����]Ȋ�-f3��έ�ҙ��n�d$�ێ��SKeFO��6f{�8a�ú�6]��q��B�U����x�מ�Br�s�j�>6'���é��HN���#���Z.��K�>Oݾ	䃫�B&�U/�F�w�" 	�i�S��k$o=������ʜ�K���w�!��'X��L ����T�#\��ԫ�i9ر:�a�D!��At`��ˆA�A�hFp�:\՞�67�	�K�5�|�(���j,{�]�����gԄ�Έ#Z�	�W�p���d0�yaFey�c`n�dK%��y&:~/	���o�`�,�>a��+�@��IX���]Hhf$"�P�r�ک�C�BX;`CI��$'l��؝7���$��lJ�+�,g�d �.��p<!��'�
	�o
��m��Q��}���6C��� �"���/��+z�W���$�eX:_��Lm�ba/u�����7���ww������MY��<�www���v�ݨ�����9矴T����]O�uv�F��AuY�5� }P/��8�����mxA��K�&��%W�p�Ֆ�dZ8fvY�G�)(��a}��}3���k��,B�Y4��^����%H��9H������퉝:V�a�/r_��$��g�$S�@�ǽ��⥮�Xk�`N��� %Y}?�+X�%��Ci�j��߫ W$c�����_���3�_�����/�TrIxO`B[ӕ��Ǎmlc�ؾsm$@�6���ml�6�r����)�g�,�CK*���n�SK��� �t'Vǅ���!�������Т�X��$���t��s/f]�n?�w h��J���'7��]�C�Q�I�������x����Q����O�3�� A����b���,<HV�>�����>�o~�gi`�M9���ށA ��{��� �f�W����lRP�������A��A�V  ��|���OX��q��>��N����V��A�w�n<Z��Y���r*�^>��/�ˢ���2�7EE�A � �L	������m��@��糕���&���a�m�1@��Y-�
�.#X�c@^ ȱ�u+I��s�dI���7�hQM遰�O�q@��P�o&X�5�UA቎��\bTx��Z
�5�踄�r���A� X��4dB���KU��t�<��sLYqUL8~�T�	b$�f9$��Cx_T�{֎��j�a������肪#�\.}���|�
�rp�> �1�����}� e�$��!�u�@�Y�$���E��~ G������I�yz��
}�� S����j*�5�P�+f=�ט�+��\�\Wg  ��IDAT���:
� ˪�B-u�3�ƃ���M�sn�x���H�9`���Z��9x�x<�Ho���"��v���ì�4�g��sU�+"c�*��õB5�bX��'ѹ��8�z^<w$ZUs=1���9�Қ�Uo��֏}늆+1Ǵ±E���f��[���9�b�:ױN&n] X�=᳛��~�?��w�c}B˾�\��'u+����e�@۠���	}	+�سUHl�հ?��&�06I����w��Lb9��"�&��"����xq���i{+��܄ڌ %��t�3�%�~�IA9��Z��z��}4q�%��a~��0x̴��bs=���u���15��㥪���/B�;��K���i�uqjU��+	����$|���BS�W�C�,�7�,� (����s����/Ɲ��w��������k�3ɒ�(��B�"������5���>�}��(We������uPӚ��dX㰨�����x��"����J����b����s/�2'�%�rj1�Q݅�]���O��{�5�e��yM��F{$��?�>s�"�>=+x�
P��"�랸{�r[���pU��{���1�����#~�J�Q�z���'#���q?�L��������0�ឹ�l��Z��~��X'S���Ŭ�@�L�.a�G'��'�ּg��F�A(yo�TP�@y�=#gH{Bk���Fܯ'T����/��{�%�}s9|����\eX��6X[A�2������Q~��_ʛ�����3���������o����?Vq�~��?���mlc�w�����6����O�� �7V�>[�����V�U�ŝ�̦>L�s�m��<T3�a��Pt���>����5r����= W��$���$ru��ϟ�˗����{V$Vǃ�ר����� P Zm�[�N���������uW�����*��io����Q��߰���U ��>�vP��[�4����D_܈s���i���7��ŀ����xr{ˊ`�~����_z������P��J��Z�Y.�>�#l��|�������{�g���V5�Ѭ|6��$���2 N-E3�N��b���zo��^[<оy�FvP�x�"� +bDRGV�m� ��6V���m�N�/�3Z�x� �ց(�ͽ{���9<`��>�v�a�m�g�*T{�� �z�d��D��T@#Ж�]�{p��{AF�i��
`h��a��k��~*���BO�SI`' <���Y���|���L�6�L^�~q �	�	`0��rk9$������ϩ�σm��t"'&u%T|� [u4�R=6��o�?�8iap�G��5r$��&g�5�ì��##,��f�!�Hc�Dvmp���q���0���ӷ�;��{��b6%<OX_Q���8>��	,� ��� >�Ŏ�+�u^Ot��i8��7���#�=�K�q���!�X-D��8.��32@�� /h��蚍���(��UK�Cu�,s�w��J{d�J�ĕ �j�B�2SX�P@%6��ǒy0i��)b��*��|�X���ʝ9�]WX�M�sv�U�'�?�F�8) }*}�2�$�,4����(C�}<C�@�\*#�� ��r;"�6�y��ֳv������'�v��ae&'�Y������ {�.\ԭ�ꧠB��@�� �fa�<��,�M�̺tX�WW��r˽�:��o�ͬ�b����ǖ�%g���s�*ܔ*!?@m���oև��X�׶em*#�V{���]wWӘ�����ܠ:��3y�3�OF��?��A�������ᜡ���u�`=7"'��u��G.F쪡�bq�'�Y�O����5Q�*�KK��T}��c���C��e��"���j9X^�r,�hgT)�Bj���«��î_��'p�`�(�~J۵�����\#�BՏى		'��C����ةmw.6�CX��U�p�e�V�8�SX�����g��޳e�ޮ��{S��(S�$��l;��µ��k?φyb��*���g�V5��'�x�{������N,,܈STTU�}��#9��y�c#�js���j�Q�Z��庀s�=Ad
`�y�>��������}�~:�#��� H�醽�둎���ǩ���p���b*�F�S�b=K�\OqLUb'�%�/�9��Z&]n9N��f�Y�ٺ�RA�q��I�󚃣��� ?�3�y��������V�WW��_�	���Q5�I���r�c�$�&C�6���ml��6 c���6�?��	Uv��{ E�(V%6���>c�28Z��)��ګy���<��F��T>��C�\���W@���U#ӂ���D^~�\�<����B���|0~~�R_#_���~���GZ�<>l�o� �G`�zn�4<| D ���ݪ�R�fh N�p����`]�|0���>�x��x��U<h��mNX�0�d�qC|��ɍ<}���^���tb��~�v���d�Nd25{�s.�[�8K"�����r"���T��c�������T]�;GX��J�h.�*��?�̨� ���fp
 nP���W_ɩj������n�;P�@��0�av	Z�Ÿ2���@�O�?�e��Q�sQ�������)����o�����?gH�w���u~�h�$qp���k>�ENg���1�ա;��!�ه
� �`>TO�@�.,C�o�w�ZC�E���'-
F���
i��h�S�9�Gچ�n׎��y{���l-ȴ�7|A��ۖ ^#�Po�2⠝�ZMB�K�߅�H����hu� _fdH���I@�W���1B�qok	���j9T�53������p<r�&W���h!������+��k�	�-�s ���*+�
�'m�+f� ؅�Z֔�0d�\T��5!���s-�����_7���>�`jH���O`��V�뭏kH`6X\�1>�2����l�V����x��� �ۿc)u͞�칰P
��cAb�s��������9 �����Ҹn ���٭!{�*�'㌜�c�YFL@�Ǳ��s<�vc���l�Ҩ�</��d[]��	��-� `#��*��\=]�|����4���c��5Y�c�����:�5�-�{�6K��t6'�p�c���
�I| ��!�$qb�w6�=b�D��噾f6��E�YS�I�HOSKD�M�~n{9W�7��u!S*X�e�x��Q�5I�H�v�������ܜ4HtZ0���>���麀<�<+��~��))L��p�`�GUA~Ά��v�?�����z�<�0��S���Uj(�0�p>��f����>	kŐ7�}�QI�6c�T�}�L�jD�Ƒ�'���C��b6�I�y��_����1�)�ik���h�s�L��, ��a��X���Ϟ=����<��#p��<�>^����H R�$5�X�)�k�{)��P�t93$�@��P�!�C�9f6U��"+����n����$,$�O2'�ޠN�}P�b����;#�#�]:H��ܩ��Z�D�[PR`_��kkSFz*{צ����*(*A��'����L>����Ȧø5����gX��@>��ƽ��ufO�L�4�"�4F��<�t�[��jB�E:w��PW�"W��8��޽}��u�z_^ظ�_(�qRnz.5e�����:������wlc����]k#2���mlc���ʫ���k89 ȶ�����V�n\����A��x�6Я|��`kK*Ф��X�+r\��kɋ�Q��PF��d:�H�췏R]-�f����R5�ɏ�\^|�}��/~�@����jT�A���I��t���V���# ���  ��O����U��=�P$��t< N�	M\��8B����>0�� �z ������B�8���fK2��Y ]�7r���w��HX�WzN��?'��z������˧���ŋ'z�*}N��z%����������$�i)ddH G}o�� ����o~����}_�|�����Ky�W#���VcO�<�C43\h�аږŽ�l�����p���U-��y��)4�޽����� 6K���
��fF^e9��mp:
��L����H����^�f��z�<�EX�:���W�@!�
2!7� �Mk�*ER�.�o[#}ɵ�'�5*��:��FC�v�#TP�љ���UQ�	[�o޼��lN��luZS�t�[$�X�����z�8'�VN$��{���S/PE���>�n	�6 �q� �� ��c2d"0`�x���x��I�}`�qP7 �@tҹ�{�J�~�%�΁�s�;~�Q�������'��1!�DN *B�<�,�'�r���T�<ؖJ[�`�����sN�]XNeB|[�yX�-�3�.��X nq>vL=ט^�b�3w5	�W�th��v� "����b�I�,' ���:�:'A�.`���q��|^�<.|j�d�X��r<a\�@`и��B�x��{����ͪ�8��a�������j�ytбP�s'�	���ĸ��p�;ji�y	q��c-=@�qA����s@�ɳcZ��BC�욨��~!����G�5 �����ܠ�N������^��
�)��v� ��%�W���C2�*��Y����:�����v�$��v �C#�o"7Om�Y�e9r�@\QU��z`2�r��؀N��L�*f���	O�Z�4뛫�Bg�qɵ�׋t��2g�o�k^G*�1����uNc|T��6k9�so�*�$2�g��׾SS��n����GTta}̨p�����H�nE�.�&i�c�@M�Zޟ�b 4\��xwo�ȏ0u
�\��hc�"��oQG����ׅ$�_; āh"a�DaM�4!����*R��}d�;P��#G�`m��rw�9�Ѡ�����#\+`��� #X��y��Q8�̜�ڈ�
��Q?�$Q���n�~e
\8�=��e�I�*i�p�뺁c�F;,�8��"�<Wۉ�#�GAqr�?��_�_��ϩ:��s��	U�����d�>�����P��f��{��_}�mP�Z�>�bR�>���X���{�c[�^p����*�#��Lx�J D�Ĉ�A�{S�}j�V~[�1+�d������LEǜ7�����	��5E,М�=��7k�q+j����u{�$a|�\�q�q7�NMZcne���1�4p=���{z���)� *��:fd%�F�z
���}-�t�+���g�(ֱ��2�@�^2%�������^Q��p/��a�A9�k�/2���Ls?X']��B�3�ՙD:<� ���6��x	���mlc��=�}�R��'gkZI%�h���Y�Kl��⡏�W��z�CR��<�c�"7}l�J߃��o�j[��瓘U�ϟ=��<�b9��~k�D� ��pU���z�@/��D�u�㣲���
�TjDV͇���}������)�}�
9T�ZU�I����XiBl��~���cX0�#ՇT���J`����aH8*���¬�F�Zғ��������O��f��KV�#�|:��T5�*�9*����-m�N�K ߰߁�f�� Ռ���d��p��^��s���8��>L� �h[�����R���X� �d+DC�a�`�={�[���zU�[G�n aA��n�y�{���V�BQ��W��`�}_�&7;����?R_��mr��u�q0X�uȢ5TsT$S��������c�OA�n�D�1=������)�-H'�Y�2�,��W��H�0�*8��*8T���G�x���߇*��E�>v:+XB�A����v���@���2} �P!����V�dX��M_����� ����� \w'�"ڑ�lY��x�G�?y��E�7u9Xk�Jv��!�ro�O����Z?���� �	P�ss�ټ�)aH�R4��˅�6i s1�*ˉ1\�6&1-�+CՑ��aV���N��}�9�!�&P�f;����Fb��J�����eV�e��ԍ�\H��T�Pűߑ���")�u8���é����V�=�A���u��֓bf`�۾�l=�X]ܵ�N�aL��@I+#l;��e5��kt�L۳����������7�\���Lmu"0K[&?�0�c��<5{���xk9 AUc���)��<�~K�q"���,@�Lm_b.���y:��сd��I7�� �c>a��Kb�Alv?�)��&�x�����K��uF��P�Ko*�$lu&f��\�Z�]�	ǩ^S�a�Fbe�X±P} BB��sS�@U�Qb�r,�
k;��p���F0V6�5��%|�d'�-��L\K� �{��N�Md�>�5
�=�^G���
���=���_
ֆ���yV��#�yU������W	�a�[@�r�����W��1���h�q|_1�A;#8�ij�oc�PzifgC�G��Qo6Nf��J��rb�?��������t1��
ރ|�������x_���u��=Y��� �B5f�a�e����ا�ֆ��@n�nyAp�
�����������hU�~���qW�~k\X�ϓ�Ԋd�Bv`�u�)�r�.ú6e 5|� ��|��}�s�4F�v_�v��C��q|q%�	j��� �1�ҫ��̉����'�P�wb&�1�=�#vK��ͭ�|����_���z��k��_�����Ɗ?�oHoG�/]s}Y�z��΅;��������/_s�Dz��%������l�����2���mlc� ���6�����$� 
{z������!�%��a�&J�)���fp  ��Umuo` .x����nϡ�q�����l ^�xF��_}�F6��FG�[�ʹx�s��#W�A��H�z�d5��a��9"��Jh�T���qR9�����lAz���vP�����:!����"�wB� ��|Y�f�|,O�<' �]o��qKp��{g�Qk��Ge� kՎ��<��f��|*��T��**w��<l��	���	����{�i�T
�z�^�'�0��q�z�C��������U,��\�YfN[�W�Mî��Lr�FU=�=1~<s�6M�g2�x9lx���'����O"��{���
���p;{�����f�mV�n WOps0�pB��lN�Dw�@��@EfY�$Vy�դ�[�� U�=��_�K`?T%�{�3����P(�XoK+������n����1d�4��>�Z� 0�`� T���x���>���`q^'�W�E�� _�=�470j�4#A�kU�'�����l@$�<������k9�(״:��D˝� �U7�]�1��Bݐ��>;�Z 61ߊ����B�H�$p8������~'��
!�6CIֲ�VIE�.�zz���)9G8�vU�`���������̏��� k*��C@2h�Ò�Ѽܑ��Y,sV[�rP4�}G*�0���%�Ծ�5@���(���#�2L���B�*8�� /�+9�5�����(i����!��I�y���ݼ k�?�)�k�-�l����Jz8�7� �\�J�-�GG��I�rΠ?0�J�nZk�Ɗ̇>���k	��ئ��6�n�C�
{ ��&�O�������������=��d(�9�`g��{�����#}�byƽ�����r�"��FKH.���e��E�B0E���r:(�� �a��q��-��c�� ?J(t�a60�u��AҦ���Ú*#Yl�n'AU�1� �7�j�� !��[����q@>J�!䵅���0G�:��SW]`1���]}��N�B	��t�}<����S�^ֺ�iȸh��Y����7�=�A��^��a�p�VY�u�s=\�����@\�����a���R�!��ly�h�f���,��~���'S�@�VL2�@�K/Fh�����B�RQ�x�ŠD�~g90��?�e#32�n����H��Bb��k:[�? �E�X�P���0�}��!�����wW�N��p� ���$3�\�b����-�&���	��$�GV���q���M?j���,ʍp�c��"���%gHO��p��~�6	,���/Hk���+�@}C;QHg�Sj�X(v�{�l���T��S�������sMb�̺��:�n/����o'���>'�Aӗ
[`����PbY	��)KJ1[��UEfki�\�Ǉ��۷o�E�ܯK_s]ϐ����\���+y��c�<{�N��z��y"sX�x�rdu�j�{R _���6`���Tz�ܐ����6��}��H��mlc���$�nic��``#�pLVaz�4��f��U�fn���K����}��b�ᝇ�⁊�����O1���j��"$V���C3���>��o����C5�,����\�+&xxȏ[}�3�� ��#y��d>3;T��	(�>l7�9`�}����P��`�����{�֪�{{ƙ���o������%�P�
.���'Onq��/��/������_k�6~.@@�R�|ƍ�9�a�vЇ���QVWSY,���wr�Ϡ]��.�{=�ww����c��9�J|5_�&��?m�\������%��~�� zV�_h����7"V*6������m��Ρ:迫���L>�����ܬ�8F:WKt@�c-��U�l#dK����]ܺ�=X�,���2�-3@����*Z]��=x��(�n�w��������1�� 7쌊IaU�!�W3�k�� ^1�acv<	�C�>�*��fC埅y�n�y,[l<[e5�&��r�3��Q��Њ�C޻�~ndΌU�&�����Enի�Z ���U�����ȶ,�C�)2
��#�Y�Z�U�`�1�m
-sb��Nh�r�A����W�Q�>���jT�vnk�x�J�E��v�a�F��k}��-�����x�]k�ŕg`��Ԕ0:�uI���f%��k��$�S ���Mt��%�N���Q����Za.]�pޭ7f�S�Į��]O�Z8.��`a���o$��@�/�Н�s��ʵ3�G r�<�Z~}s���L�n�u��C(? H���͆y�*���A0&A�N\!�Y��	�4\3��s����{�~��r2��{?�bo�Go1'6fy�xȷ0�J�dC@6�{u}�Vu8�5��~�^���s�ek�L'	�0�{���gOy�ȳ:��ZB]�1B�n-k��?�c�����q�¨�.GڶMrWGB!B�G� =����Ѣ,w��D\�R��G�v1��li��Ƹ�_-��2ѽ�z�*��Xq䚊\���e*?H~h�M��uL���p��-�����������>Ң�U�b<���Zf+��,o�H^�T�?�M=b ��w�0�D7����	�X���R�m^]vN��� @@(��<���gO�q�tl�\ T���l�5Z�U�>�)*�˦��
#0&z���K@����4�{�W�������lȋ���ז�,=��D�p��a�\TEյ�%þcDhL�7#@�E�{�C{M�j
�/1��B�8���K�˰��ɾ�����z,�4PP[��ׯk�׫#a�}֣�D���ߏ���1����z�|N�_!?Nu5���L�p�Ƿܭ>$D>��H�?T\6� ,1��'V���{�-ǅ�z��2er��B��(
�[�G�ͮq2!��6��˳�jg(B`�5[,~ ����ׅ_סB�=�G
�b[K��;p��k��g����	@X����<�(q�փ��k�~-ծI_p�{�����G�ˋ�/�ze����J��(��AF�B��Y�]mh/�>Գ/�>����A�/A����c���H��mlc�w�����6�����Y.�h�0e��s}P;���w�"z"qVx�n;<ܷ�@E +޻�]K�'q�>�<[F�>Xu ��L;��؃>\/g3Zk�v)K����Sy��>�r8��0��w�̩�[룚U�&)q.�RϚ�B�g9XQ�	 u�Z�{�4 v� ��O �$��f�5�O�������i�,u����V����3���k��~`��x���|Y����V�]��a+�w'o߾�����^ŰS����(i{!2�/�ȇXa�_����9P�v?�Dꥊ��yR,H]__K������T����ӔU��})�#�6���������K���)A�sOeT��apb0@� �����>�wT��+ �,fKV��_.������V�+k� �w�Vlb�j�W"�2�g��ܾm�l@"����s 40�慁�󴀙d���P�k	�)����	�ϊ�`�;
X��&����6 }����5?7X��J��hu�py#�0���HV �Y�����=+�cd4��*����3�"����8 N�2���w �{������u���ȌȂ�G��8y��рt��ɕ��	P�pOp;<u��qL�� ��M][>�.�*�C��^�c������|����!�h��1R��^�4H������M��w��|$��O��2�uȦ���j�	����v[�Ԩԩ�ʛU�ӂ�P��K����-mQp\u������o�2ofR��`��J�7 u��D@t|vS���Ү���8�JDE ��w{mD,��8[	�Z��_F�X�y��K�z��DVs���"����Ã�~�sEfӜ�~�����9���cl֥Y�� ��J��A{�z��f�Z��C�KFkd,��A�$P��N��?H�gϞ�|�"8h6F6�A�![	0\Tx� 檎����l6�yy�ύ�$rP��-��s;��
�k 	�Ff��r9�I��XƘ���l�_x��в�����mISZ��"��`ޯw�n�Z�J�s�o2���+��`�k��܄2�ýx�%�B��@��X�\	pcN����ܿO�G�R2�~Cc�kB@烩ŌĀ� ��~�cl��CV��A�r70Ċ���] Da	2�$H����:�҉P�::��uU��t �.�o����Щ�LT�n�e�?�2�� ���G�ydjU�ؕ���$H�Ќz��I2˰�h�Y��h��2�w �Ú6ا9�jy$�
����O�c���ޛ�$�i�vtH��2"����o��4��Z�3Ob �{W�vfmU��yo�}H����}�����lio�V��kQ�B�Sʂ�l {�{����}�t�"�=#2*�)s��Nm�ec���.�B�ϾE��ò�'TZ��W&��{M�VMuS�Z��N��殀\�̾�u�[�[r�>�wE!�8,�t����O~�#SXV5���W+��Q���l����@��x{��,�Mpd]����t��kM�JQ|��7��W_}�y�1��^����V�X/Q��$9���V�n�r
�XG�D%2�X�䮥mgJ=��l��$�,����n�����b��2���mlc�N�� ���6����4�k�9N�ԥ>���[�F �LB$���I�\,D��-+!d7�|����z^pkA}$,���A�.�fLV��}��~�T���K���V_sǜ��<ȹ�Oe���2>��hT�Y�.�Ԁ=-��xi�b�*��+�=�wznI
֌��~�CA�	^�qN����?�?����	\��$�b�d�r����\�\�9�h�C�7zNz؅�/�קŌ���{�Y�{psuM��Bۃ>}�i?C��Hf0WD���#۬w������=�� �C��샲�q�&��0��z ��xT��J1�a�DAk������Dw�_�~Q%�D�bx��7��{\Ӫ�����:�H.H	
���u �����P�@Hx�c, @J�@ɒ�&�64x�GkD��|�$�e�n _�| 'A���dCm��n#��sϺ�%��.�2@9 c�ΰ��� 9�~r3��I��80J%b��B^G��� Iv��<qK����H޿#����	N:����b*�dj _1!���Xo6N`l%H+�N��V�7� ��:�S ��
�T�cMA����$�6����9η�*�`-�k��f�s�} �%>��y �pܕTT,�=`�ĵ
�%�a$"o����@NqM��0RT��v#ͩ"��ά3� ����P0C�i=����=�tn�5�cA�:mPZ�L������ _�倄��r���ϨM����0��`U��auS2[��J}�,!d`��P�0��E�P�~ ��g�#?��&X]�G�~���w��H�ؗ����9wM�B���G�� ����Ph'4�YA2	����Cсu��P"���YLa<M����@\���=�k_���ʓK��qܖ/;����b��*��Kl�������$Fn�jA�l{�I��, ����k"|�ѯ7WK�� ��`�VY���*�Y8aԸ�?״8%Q�.a���߇;�~�gL��VV:����=�J��2̌�m�B�D�/����OÚ	˽��O:����WW�@*�.�Y$�<-�p"^S}�=Og�d�`�r�ձ�f�r3�,JLQ7f�;��}-�٩�r�`������<DP��x��b�n�R>(J���FF�[6����3"�=[�@X���O�4�y�0f�ec,�q�I3UAv��!צ��.J�+�C���n|������l��.�:Z)	�>wF�{�qw�‌D���5h��ռ~�����lO5S��ޓ1�1$��ȹ��>�>$?>�:�m����<�	�vA~�U�V���;�KB%��8�KJ�$a�Im����,�%��G	� ~�p���Z��^�o��ot����Rp�Ґ�j�`].n|���2�3#��0�!u]�.l_q?x@ADadH�_���^����	�]8>�b���|��7�����JE��z��#}����$�Ә�G��6��l5��y�'N�"�9��)���l�����6��}��H��mlc���$�Td0����W@.X����I ��Z<���9]��-�}��,��+?K�$<8�nSV�Y�BL���˗̯H<�ņ���s������{fs��>�zV�E��j�p��z 9�Z�Ws6��DY�^d@���k����N�~��kG��G=6 � :PUK�z�4(� >�Ńi./?z%?��������� V��@�<����rw�5���L �6_�
�i�Je=��x�>�"VZ0�@���=��x(	0 b���f����;~���L��v5������I\FE|���t���kz�{@h��/��%(,p��д��o���1�q�-l"r��ez��6�� �_}LE��8�Ή!lmO�n�S�7�>���p.�[%�
���JU� | &`.a|4%�s*� |��j_�"4^�*�Q��u�㏯�II(>P���C�i#9�y+�eBK���Ϗ�D�<��w6 /#ȪS��&���*�GT��(����*��$�k�Ya>&b6YT���b���a�0{5#�Y�����G:���A �t2�ۛ��#�@�y�}oa�B?�����T<�#�� �@(����a��^��� ��>:� 4�(쀒cdU�Pе5�guJb��yH�^��+���n{�����ha7u>����`�v9�S9P�?AE����Ah�= �� '9�Nˇ饯;�?}g���>�,W��� �`rK@� (Nuc��!� 6K[#X��� �����H�	A=X�����Z^3�;�l�\����md^�
S��妨!qN�"%�q���s�z�˝�a��x2�D�\�3}яIL�m�V*�	����?�}�{���,N+Hu쑪�\]-����*w�YLa�\�>&�nc��%X��i���x��>��R0� � �\=2+Ĕ���	�#�����H��Yf��o��r�=@\,��,h�q1�}��-h�!g�ֺp��b����?4��O�y�[���-.{G�c�a�I�9
R��3^;X#!K�cx�(�[E!��i��e�ǎ}��D)�Z��5W�8���k�_�*��d2(��/��\yU~�=\{�����'gҤ�߁R#��A�̬��(�'�.T��DGF�����-Uae�kN���'����ܷ�+C�� Db���%�y|�jD�a�Q��_�2����H�ׯ��S�Z�{�y��-#̔ Y��s����WT��F*��:�M�U��_�e[��8�o����'����$��МdA�K�-Wڴ�
���1�t���+�J5�;`?Gq��}&?��U���dVp,I��U:a_���E��H���=����s������t�c4��Ld,���96�ߟ�H"�[�{�0�$}����Ͽy��*�����?��|��������~�+y������_������˗��?��ܾ�8�Dz�ǩ�O�����H��mlc�w�����6����O��
�n��IvGmc�� � �[%iDp���{C��;�D[�V=��x؅R ��������:|��d�޳RY$u��Ō� NǊVXS�(a�C �!ѥ�����@	��*�`oA[
 q��XV�I�b�a�q��I�8��H�w}�^�IX�VS�����O>�2b��5�� )�V�={�_�����;T���Y� ����R�� ��ITÞ���*:����w��g��o~-_|�m7�oO�(�0���凒D���^�cT�ۻwz��@��5� ��x`�|�b6��_em5�*Gv@��V�ɉ,��F�� D�scIfıg*��@�G_���������> :���(&��!��_��8����H<�;�!H�iSC��uu��x±��@B��j:[��r�P��9���W1���LV&��6;#z@v0�sAhar*��P�x)�7?A ���&����~�Ti%�'��4�Y��@u�܀9�\:q����TA�`�d8�iNU���bꟵ�-&9*� �|�c]o�̱��	����FB%B��W�/��삟�D~+V'RL���|�0WI�ʿoIL�r߫��ics�����&��j{ڋ��!XA=�T�m��X���m'67�{T�Ê	$V >
��P5�����C�|���i{�G̥�[� @<u���~G���U
1��� �,�C�Vp�e" ���ځ���USuC�d,>�M#iOH�js�nG��|jsVS��]{t��0�3Z�a��+X�-X�W��$Uq��],V��|�b�2KW6��I�~C51����7:��;)�'V:'	�6M��k��������?���t4�0���.+S䰍 ���i��U AD��є���׀�~�5�<�5zS�@؋x�t@��u�s��n��^��k��kV�S��?�'�+�#���*��y�#��Օ�I��G� ��9I\��3!,\c}�9�c9G�>�'*2&��QaM�\�
��b�J��w��	���_��q�L�-A\�#������E�|Nhw[#F�X7�����Ș�.�=��P���Uu���n+�i������5in��i���#/�+냩J���Q�@[{z}]���=��T���y��<�D��k����T��"^���+Z�q<�,kk<
%�TUqd�-5��ف�:�u��8ɝ�Bc�$�g�)B'G��Y ��;(� Gl��
$Y<!�A{�8���nۅG����9�!�}�o��yOļGl/r���G��kk*]T��ɲ�γ%�7� |�<�J��~�Vb��(fH����9���������+������߻|S���e���*�u��9�s@?aN�iU��j�ӵ�CX�n�XB�o.��$��&��J'��n��^��P��^�V����~���#���s:؏�-�S挷v��� �T�FP�b�@��$�S���j���>�ߕ���&����7,6@��Y�u�g/^��{|�ŗ���/_�{���~+�ݞ�\��?��X�����S�PE�~�7���X��6���mlc�N�� ���6���ɴ�n+Wn�0_N��1%����8)d�\��j�L>h�����(�@��A��Wy��_s����,Θ[qԇ"y��`���(T�}����Se��]!��c)�É��o����r�\����G��4/$�,��C���#7��g|
������>�g��rܗ|�G�,���Z���e6{*�"ѯT~�����oh������J��Aۑ\Nn�cfPud���Z"�@��
�R}�|����^�A5�"U�V�凥�ó[y�͗�}x/��0T��
U�O���?���{���*y 6��F7oY=�E�,��y�P��ruZd��k�	�]]]��{w$I��gDE���� 0���s<����Q�:�.X�	�}<þ�c�FK˖����U)���X����K�����G�dIhd�� K(2[����:`�vP���,ZIX~�D����X/[|v9��t^0�D�q�~�	(��q{�0e�\|���PY��)�<�@@(6*-aD��O ��h���5��j�j'��Z��L:Q_�����i�3��l����YXN!f�e6��	*���]�)`Ϟ�����[Ζ��k���~�Ӣ�d�ߗ���3*�B�� z���;�GYZ����e�,�Ȯ�4�c��l���y2�H=�gU�d�^뵬e���D׏D�9K��z%�l{=ޔ0
����@�ꦭ�1�{�]�V��>���� ����B��^�u���x�{GE�rx�ܭt!��L�=�&�N�$h�� ���{��V�Ϧ�~>�P�1�m�.s�G}�k��1T,���z8�_Ο�MP�~�6*	߭t0un�V���U��tz�5��'���L9�;LX"�X�3��z�)��n<�\l-�P�������(�3��ӱwDv�ĭ��ɇ���V[�z�Ǭ�RsO5_5(h� 	���	�>�� u�n��k͖�I�I���+}?\ϊ_ui�qy��m$'@��k�U2Kfr�>8�=�*tEx5�@�����uw'5	���&��xҮ�^J�[(�N��vV3�'��*�i[6�zFB	qB�K��c�n ���c�|���@!�狶���:���k���~-t��HN����r�ɱ����ݛ�%��[��d�Za�R�R�-U)�A^���72��p���zԃ;���g:��oH<�D�c��=ɟ�*O^���o���_����_�={B��\Y���ͦ��ǜ v/�/�]Wy�y/�7���G�[���ff����wkf|�fN����^�|�\�t�c�<�cQQ���0�p����ŏ����+���u�X(q{�L�'���^�b��+�c��r��}N���������.�	�F	�j����:l7��H��	?\( �������6o,�uuTF���e�9�8�yf��~rm
=�E��]'�'�Au�=�e�Į�4%��`���L���s	2T*{�[� u�,B�ȭo+D�'l�3��w$U�x�󎢓�;�^Y��^��F�L_&z�RP�9�=K�wa?5�܋]a2�
B�s��zB�F�q�M��v��ʝ��e�۹���+t���f9! �-��^w�ǅ������A��x���U(b1G��a�;��P`���0u(�{]��������xǘ�}�^�o�-���K9阝4v_�i�Y���:ԁXc���c8.\|o�k%�k'�@´$Z����Y�AEJ �ZϤj-_kA��X|r7i���X�����:��r/�������I׈�Y`��Aq�������Ss�x5���g�#2���ml��6 c���6�?z��;�#��na�`$��F\ ��Ǉ�.�
�ci6$ w����Lf�����R��*S<��ܫO|T<��=���wk���~�����bVKį>���rg籸U�e �CUnP� �0e@DP��˙���T 9�IU�]�1x�]��� �L�?�0�,�M%o��|��;y�n,��s��|�s*iR>�'��]k`^c�c��y}�CV�h�hGU���6����Qǿ' +3�dEm[2� �f��ǟ��H�fѓ�w`����3I��i96��>�E��B�ik���`��|&���>��|ho[��۵���_cT�7e=����3�%�5���`Ɂ���MRԹ�Z�
1�.6��o�Y�:���H:�����J����<��6�Prn�B2(D&�-����e�V$ ����l�`��{���\G�Eߤt*e��wO��T2��w��Ε�DӘ o���(�r+�ÎU�umU���N_��<�6k;P /��ɜ48��t1�\@~��^Ǳ�:��D��|\�<�2	Ҩ��m]�� ��eӭ�;9��mNSy�c���s춼jP�eq��2 ԰��O[����99��:'�y����fY����I#�rح�y����B�*�(F6�|y�vPV=K�J=��o_���m� ����F��g���Rz���� � ���7�	��g��X��2t=���/ؼ��-��T��W{ \�V��е�>�@ ���X�n��q:�x�tl�����t���-�>H�
Ү���z�Nd�}��nK ����ۖKTX�f3��	a����φB�}[�tdz� w]�CV�T�Q��uj�T l^?>����� <!���s��5$KH2L|�!h�o�k�`L�BIr}Ϛ�µ*��k�uk����/�@�� .��DF��e\L�y Q��Pk(``o�o( 0��b��D�F'���@�Fmzm���;H��d�Z��v}'�^+�u�ԋ�[������ԏ����Bitزz����Wd��ǳ���p_�Om��4f�}	{�4��>�c?i�=��~O�#����a_cFT�ДB���!����Y���`���b��y�v(�Phݣתk�����c���끪�! ������yWG��4�{���B����=Ƀ��Yȱ�Mu��}�����^�WOt��9t�1W��~�ڹ);��Aʁ�kEV��(e�qqlu��~��٭�0~�)����� ,w]��v�]�9{(���r�.�ʺ�,���N2�B����ր�o\��	aئ����o���B��g����ǋ���e)�S*B.�Þ�ӿ��t���Y�@:����ek
�#��*��㵽
��
J�>a��d��i|m�Bp9_�9*<��g'���#�1��_RyX�y����	I���h����W`�|�*��9�ׁu�{Ԋ���^BA)=�m���w�?�X0J�����z�f�f�5��@��9�*d�J�GnWY,u�a�WZLV	��� ׬��;�UA�5I��u��&n�a��s6�/^���>zA���q�]h�����J2�*�P���Ԃc���6��:�H��mlc���$ _j�X��BQm{z���N���v �����|�G�@x4T�A�� &�g��(�����˘� �!|�3_m�j�7�|*�ar8�䡱0r�]3za�L�6�5���F6�V�W��7�EQ�~� �p�es�5
M�:{����~���,����OMn'm����Zṱ倈)`�E_p�NB�3�ӭZ�U���
 ��j�;�Zڞ�B���� :P��zp�yq���@.B*Qzs{KkX�=>�Yna�3��чn�����ׄĈ������I���$ �.�T�lr1�"V*�:���ݻw���'�Of�֭�����ő���b�H.I�{/!�?�~dU�>�!�6���P�;�G� � L�cHJ�9՚�{7 E���Ú����G�u LU�{v�y������! ��)T���A
�K�,����l9�d��A��T�0�ͣ��i!��4ov�S����� ���h�����8P�~����1��g�����`�q
P6J�a���&A%��?�q_$�y	�$K����C��<�WX9��	�㰼+k��61�iV�\�M�؍t�srV�nF%���>?�hz|��%�`1��$-�E�A�X.���.�ru5�J�x^�$U�
����㣱j`��3d���I�/Ʊt�KuZ�a���$e���9;I��Y(-`ކ� #w�G�u�t6NbcM�� �E`����[��i����o�55u� ��82���.�F����^���L
�T������߷�� ��ǜ�pT���#�s[Fg�Λ�xWR�T�{���OA��|1��.��ZtjMy�섈��Ap�8���,'s��2����Q�R��5���s.�#7+�-I6�<����r��:��U�n;�~�6O�8��Lb=�d�BR�CFJ�j��i��SL˵�*�뛥��+I
=�z�/�����8\��dT�{�z.�uhgQO���� 
[�A�����m��H�ێ��֤���_׋������#3� 1 ӒJ����h�J�c����<#HU���I�~� �@Z��'9��;]+0/�bJB	j�������$���\��u�X5�YFJ�� ay����B,���\Z�9�BH �:��%�@}"��T��6�z�t�K� ��dH��I���*2ҋ��b=u�Z�1�����)&�o@�A��Ա��x�+!9�u�o�ݦ<Ap��?�*}��p\���3�b���4T��W��M�zVH��	�7�T��F������B$
���2��R�=4(,;�W�ߋ�P��QemVXX��r ���w>?`�d��Kג��ovX�E��]�3�#��� ���'�=..Nr�أ�3AE��7�}����$����V>�IZcc�-�/@qٹ=)���㐱e�n���e���՗��U(L)S�Y�m����+=z�����1��V�ݗ�Z�{��+Tlf	�l�4�vS� 8~2��S��jT�T~����Z>��3�ɟ�T~���J�MB��̭��~��ҙ"��L��6�K�������6���ml��6 c���6�?���hGֆe$*��!���x�miՔ�8�X�J/����k��&���|�?��cy���U�$u��<̛�Ws�! S���`G%Ȑ�ø���q}s�ՓՐ'�PrV��L
����3K�^Y	E �8�U앧+���Ż�;�@�n��t�Q� � -5�F޼yC��� A� j� �|�2s�8�JЄ���ĐNZQ����FV)�=��,���c>B:�/�f*�!��Z�[��g!�͖Ձ�j���A��h�C��Ia�hcǋ���ET��:.N�x��4����n��(H"}?��ZFFo~� �(0����:�1��k��p��=W�v}��>g|D��).��*Y�؂\Ŭ�,�@$���̯��c����2���+q'缈�+�ݓ��"VmI��!�<���5���b��z` �Q��XE�5��BU����3���r}����k9�8}��a�|�� �ϳ�[#r`��=����R��(�S�bJ�m�P`H@�`n5UG�̧�
�2G�>��3��w��;��a�5Mr����EP�k
�����xz���P1��p��Oi�3;�z�͚�I�ɓ�:Gs�Z.d5�%���2P�a1��T y9�`��@���
(��w/�~�p�yKX �&(��	�QZ�YQрku�@�
��J���_�ޫM��J<.C��Y��B� BP��y��o�}���s��|��gz��M6!
��L:���s=2${g����~�ٕ�̈p�~���13:ǇG2�eg865B���A7�7���ׅ�x��_`Y��k��kfm&���YYB0:t�TT#��:�bg({�;�H�14�"ċ̶�8r>�󩞣ϵ>K]󙵴��s9�*e��|�޸�~m�_PͅS���`�E�ށ��1` hfy�j��cm�B�r���{\���q �ZZ�	�C��U�,�:���3,�;#����y�� �f Z�w�N�tL�;l[�
�1iE��|vF;��:��B��������`�3aMu��t#�¬�,��s��m1�����#��Ƙ�#[}���ʧ���1�@��
"���m�2�xި�}��ث����,[�P��N��r$0汎�S,�1H��u����/Vn*�
����ڬ�ᏹ���F]9��e(3���p��9�\YX��#�1rW�2����h��!^�U�{��ʣ��0Y扜�<!X�q2Dކ�����[ca��Z׶d�����؋�(��,�^W����ƾ�^�����9�l�x��4�{�0�5��=�7�J��+f�j_�8C\e;U~��+G^��gF�0� 4I���2�����p�TV�x W0�� �p�"�(`@$�\��z�qm��y�-c��_.��.�*/������WA�b��L7�s�P�����"����v?��V�M�.��$t�9���>:j:�
�ej)\gf��r����\�:�7T�Ebd�6����½Ω>jEH�E�da�\���{���E��
>\2�;�J]@ն?����WX�z���s*����s�)�\K�u�
���{'d�"�s]V�YZ1^֊t�c_���u��+������+����+�c���9P���9==���]��_(Y���Ν{�ʽ��M�u��{#o�l����5�iMkڷ�5HӚִ�5�Ϯ�R�I�ͦ�,| B� " _��Y,����1
�L�g���8d� 1������5B��L��)��S����U�������JW$3X�)��GTT���2"���!K�� ���] 7�����w�zO�'ܨ�!o� x8EPx�k6]��S�Q8
� mm]Q�N D HZ�Ү����B��b�����<��zf��Y�)�� R���PU�N�����>@g�(�mNdnE�--Qq�kad枠�3M��r�� �$I���#!fY1 G���>���=�=Ê�h �P��j� UÝ�9VQ�� �n߬C�!R: ܤr���^��K�M5@TW�^&7�	\ h� �������ߣ�xż��G�}��>�)��3� ^�UۀR�ލW���#�}��G]�rz>����#y�tB�C�ߗv'�ox&�s����-��C9����z�>���Ż��1�Q	�1��;�M��q��5�y�Xrx�ϱ������������� �V�j*+ ���9���ww啗o���#�u�H/G!>y�����t\��j�*����r���*7�^�+W����>��8��}������
��1�L%+�����W�<�c���c��~�����ek=N*8�6A$!�!�w�"W�����\=�B��/���}��de��2r�.�Υ���q����oK�kA�{�#�9��3����1���܎C�`�ԩK8����{<�{/ߓ��X�|����'�/��L?׌�<~.���|Fe�tׯ���gc�Z|��2����0��yϾ�� 50z�3�A�'�{�r����q�x��ǲ��!�� ��۝���aŹ��uߖ^�C�5�Gӓ3�꫇����d�%���(!�	$T�c�_�z ��@��d��'@����g$2�+�Y��X+�]����ܿ��ھ��?��_=z����j��vCK6���Z�N�`O,7�]��׮l�쩼�����MT��~��~��1��soO��y�;G$�&s=ߧ屾�t}jUֶ~b=��\Ec>\���[7���5@��|��{2;_��6�¡E�I䇀�)hIs����v�΢}��ײ�=�r- ��-���Ε�Wu���\�*{z�1�?���'��9��lx
ݣ��b|�q��￦�c(w�L���:�?��c���c�J̻п��X�*�"k��݁~��\9:����D���_?�9��D����<�B��s*|eow�sP׎���_���;��cFŦ�*�3��*�����ݾ���C��7�?|�P>�9|rz���9&���,t��5���c���{�g;��~�|��#�u��f��J�m�PChe�YYeYP`� ߢ�+�!� �Z.���]]�����I���Ǟ�r�f]�_�a�B���Dރ��
�PP�m��ʼ"�o�������I�-7$�V�~�����2YP�� ��,��ߣu��A	5Ԕh��Z,��~�3�÷/�G�Stm%!��atHM��J�x�� 1#�� ��I�1&۟�l��ɣNb�i�LϞ����u�����)�,6��WR�7� �~T�[�V�n�7�[����C�x�Q+G�V��R��c�I��{����y`��q�+]70�Ȋњ2�䥗n�[�}[��u]K�K�;��d�~�����?����g����Sw�ܓ�^{Mn�����%� �t�^V�_Ҵ�5�iM�V�� iZӚִ�����Α<;}���@)T��է,?���s�����-9���k�6��Y������|M;}������/���l"Ϟ=���3>0�a@�`7;��UL�@0�������#��Ҵ2�#g�`ȿs�N��:}8D0lY�� asXP�Z5������q��|���qげ�V�H��UA�*���9V~:lz��~�7�s=�
x|��Y�k�oSy���a����j�+GuwZl�`}��J�J�l:�8�'cߔ	 NNgrv~��t���z���ى�gsZ-�z�����GEܢ?�p` �M�w1�/���P�ª	�Zx�$�P�
�~/f,�; �j"��UK�=�}_��k�h�8��Y=�su����ZiU���囁��^�q�t�~Hc՘0P�{ڇ�m_�vg��2zoa�#�V+z�۱�#+�K����8oE��`БW�ޓ��{���&q7b����s��#�o��oe29ex}�ڕn�@��:�׮˽W���;�d$�Ύ��B���W���:�Ωb@�8rP}�\�	��:��_����r���q]�d59��|�����AٰY�x]����ޛo�[o�%ׯ^�[ׯhe���\���?�~����8 0�>E�x�����{��G?�	����g�'�����?�3�_@������	��y����ڕc�r��!�A���^�x��|��sIv��4�;�o_"�Hײ}]{�����H;h���k��l��_��LΟ���O�W�p�A��� H���=y���r��]�DG;�v����>��>|&	 ��2K��2?��c��՗o�+w��9�T�����x~�D�����<{�T��T��Q��\�5����Wnߑ�^zI���e���_��/+y���n���1յǋ�v�{:���t��]��rE��g�}J" �1�}���#�`�|>��W��0���cd#���~+�w�<�u}I;�	6��e&�����P��t�&����!ð���o�oY�t2�K�р답J�"��X�-/]I�F�����/ҽ�\��_�W���K���60�|,�Z�;]���x�c����r�|�/���s������	��ȏ�� A��;w�Ƞ?" ��d~"�������_��Ӊ�!�YB��ɶ�Ϝb/���u림�ƫ������7�~>���S�.�%i�ό`��p���	l��ߗ�_~YnܸF���7���$:?��w-���/C�f���d��z��-��[o�͛�eo�kȀT���wuJl/s& ����v����r��u�NW�z���=�����S�W �Q��u$���w����Kr��]2`윝���������_�ޢ��.�R�����ύ7�e��_���ӏ?���S�L�h��~�R���~��d��Ř�׫�� }pO�����_�B�����A@d�r�^k�;2��|��M�_�%GW������wߑ��!(]Z:�7 ���߄��#b��L\^�);|�O��C_��D{�ԙ{��sd�AQ��c<�Y��l�[��T�Z^-��Ap��l~�Aa�}�g5�Q~��~i��R.�G��}��`����E�b�eW��8q����s�|Z6�NE����^�k�|���5����+�����z��������GsAhm���h���W.aDꨏ���gɜm�����*����bч�H���A��'�FXo�:F!DqL]��홺�$XWq]�.b�~�{D+�Af$����(�Ao������aI����3w�����\I���P��}��.3�@�@����y�0{�7ߖ�x,O��I;ʃ�#��I���3��G��l�ꝕײ^mZӚִ�}�[C�4�iMkZ��,�K�'����������}��\�z%f� ���HZ�V�����V�@� O�,%�9?��!l�@Q}��AU� �P	�Jtب0�;���I���nǑ�����p@��ǉJ�e>߂
��C ievV�ְ�i�h���ԇ9d�����EmW�J6�P���+��޷�󪸰 b��~�UC�1�ķtHz���� �gMbVA%ú�0��V�yBpb I]M�l�� ��+����Z�<���:]�;�g3y�乾f�*OT���*���g��q?"�N�b���(q\Pw�	?�v�.+Ī	9�ief����jP���q�W�{���YɅ���2�g�R�򙊞�rʋpb��Re,-Ɯ���q��g��y�1_��͇�B�����
 �R8`��	�Ym���~\��Y�Dх�������:r����?����h�U���R>��C���GzmZeI�.���]y��Ƚ{w�+�����h,�O&�hxO��ӗ���Z�G~�����ӎ�����ߑ~���������	�
$��9��?����)���I"�If��wߑO>}h����8���lcU磑���w�s"{{��ztmz,����7���2Z/Ez<�)|��p����~�*�.�_Ǿ�ߣ+<O�BK���Ӧ�zN�7�<�"O�^�"7�ݠ"9>y��������#f)�ڬu=�BkF�ߕ������r썇6�u|��_��?�~]м�e�5��h�t��u���4�eR�������Ϙ��T�E8�=٠�<���۱�|���G?e�m��1	�_��K]G*�Кj��7�e�$���}���g?�7n�h8�9��5!���/��=�D_PY{��� �����^��w^�z�"X��l���Ox� pj�@��^%2�/��|	���:.�Io�%���8\M��z��&�j�h��^�2�*�d����2�H_���OK���ס��e�%�;q�ĸ��>��=�Λoȍ����������w��\~���P�ې��l.����;������5������,6y���A���r�i��F�Ck����P�����ӟ�L^�s[v9Nv�#�����s�ȸ.$�G�F�H�������G��<��.~��_ɗ�߫ٹ,f�2�9��\�>V&�΁��v�u���~B�G�2�vW���#���>0�w�"S k��W_}U~������>�gh F��,���H$v[Vh	@w�k���*7_�ɬO��ѕ+rz6�_��ot�M{�{��=���']K�]�)?���	�B��� �y�<����f����5�%�,k9_$���W�G?����~�}ր��=�7k�˿�ϲ�.is	�{L�I�i2�������o��=�~ �AZ~��'���s�73��`6����1�u�߰�C1��$�A�l�=�/Z�)��ó{��j��+r����I����8�$��#t�A]�N�w��F�N�Euih@5����$�kd{�8jlU��^��~�ŷu
Uq���J+��T`������%�D��{p�(r�:��0?XHS��&��y̬*\�GL�"E�H����9�eKZ���[����������PӮ��l��Ҥ&S����3K�*�{;�_B��B��Dbe�qT���+�0�c�vP=a��$���t*\�T[�-�:�*��j��V�Zd/�dUHdPX��, ��7�j%5�����%I�9�5��Px��üA�~:A�Y���f������Qݿ��w������4�iMkZӾ��!@�ִ�5�i�����Th�j�c;۟:��mY,����5`DA���*z�G�\.Xȏ6X&Yu]���C.l0�S���0K�+Ǉ���R��)UU����h ��CfA^���U@YlAmX��+�ߧIM~��� �ދA�fA���0�J ��LK� ��HIL0$;����>A�I�Hb�{��f����kA�l�!��^Hkd� �CP<}��|�a#�%����0|�-S��a�En�����^�̅��Ȅ�<ȶzڷ6yL��J6��Uf�#h4>D�௏p�UB@��=��ɦb�2z��!Xa� ��b�*�C�qB���x��5�p9�\�0����b�@@L�k���
�j�
u�>����L�0x Z _���%r����^ٸ~�n����X�{#t"�Pa\�+q��쾜�Ѕ�ת?�0���"_�,�z����Z��=J�t��Ձe���R��Y�m��	 ���޲�얺Þ���PY�@:H�kzٻ�f���RgoO��Zz-��Ȁ�������9?�  �p��ӎ�r�ˬ!�٘t$s0��vɓ2��kN���TIG���	d�٬�܇�#��Fx��Ң�r Ε�+|-�Q�f �Q��|�y$î�ۍiɕ2'�FJ �����a�Z[���re P1�<�$G0��xW�2�������A�����9��ʲl���̑#=v�� T�uI�ﷻ3���rAF�iiͥY !�������T��@���)�U���������lJZ�����\/�I���}�l����6�,}��b���=׻㑮�G<o,�^��@�WL[��������l�ф}H2� �Ah�(*�q\�.sy#�ə�_�׸&;:��� �{'�D}��Ν�q����B����� �4�j�5D�,�+΅��
�' ��uL^�c�a紘h_wH���a-Df���g�T;'�yz̰�;>���0еc�-;�=�}�;�w8g��$�u?���\�qt�]�zS�-^�3G���KZ���@Ǳ�`�t�2"�xO��-��A���{�u\b�e�~e������� ����C���t�Az[��ڎI��q�}P8�8����~O�RW?�@�T.T!�=���״�
�t�ٜ�~�|��m��8X����zrth(�*�٨�>2K���{�^���Lט��Q�n�u v �D���	�;��_�c v_ o�D� /F������1�n��G��v��>?�N\��
�w�^� �ai�kRF�(�gp�ҫ��� �XkPX ���އ�Yڷ�+eQ���z{ �W�rw�U{�<�{�(��q��o!�QU[��y�@�CyV�M� jUc]�A�$u֧f�
��� r,n��\��C��Б(峝�,�MY���86��B�7��JAm\E΢V����	�:�#����#58����z^�$~�W�\cdz�ƾ��^�bEE�K1��<�瀺E% J�^j���au�|m��l�-�����u,�rS�b�Z����ϧ"��j��	����qYz�ש�s�v/�}��u�b(Z��>	ܽn��vІ
P��<X�V��?�p��?����M"zӚִ�}�[C�4�iMkZ��Z��@_]Mpi:�1��a��=��x��^�X��b/���md�C:v���PE ,G �r!;����Ls�� ���w����`��t�*�0l�Z�&|��zz6wDC�jY|��m�BC��}f:��������Y%H��SX<�A%�^_ƻ���b��:-�C�!���x�$	S$F;�	t���B�������_��J���a@0 �VlV�_�!��ϕY����=��\�s�k���+샨@���$D�@�
��z��n�ԇ_ ����)
�B4�dŴJ�;��b.㝡�y��	����D����[ ���<!�;`��f��ãV*>�D��ZX� ���%�c�!/(5� T�ha�}`c���,��p* ���(��{�i+|K����*Un3Hp/�TH�"��?��
�8�l�-G�c@��Y�-�=�C�%dW \������,��9B�'�K"H,_�"�T�uYk������`��+A�rT�V��5���`�-	[X��sc�  >�{{[F�9��H�Y�86����6���"#� ���p�cY�u���q1��P��M�E ��� �l4�I=x�N`�c!�)�3�.E6���Ώ6E�)��gP� \��i�,\�:����t1Y�b$�Z�󩬗3Y�':�o�	���k���
���ꦐկ H"�w�6͓-�E e���*��p��j�1�=�}W�� �1nq����^�qMZfѣ}`+h�`y��k����(<f1a��KΗ�r}�XPy����q�10�	r��%f_�}Ϙ�����C^f��g��RV����_�����٬r����[��$�>??��c��@��o/tj*�m���be�ގ(be�dT	�{��$�5�GFz�����m=�]�v�]�6�K}�ܺqS����|�Fڟ:VF�1I$\��x���uW���`����$�T���q�dR���|�B9;�}}��)d���^���{G��U�Q��k;3EU�&`������m93�@��t�`1���ȔDC.s�3Z��g]�1�w!�ӂ��a������UIZY�6R��[ ?�X� ^$K(5#��f�A��$�+�f����1úa���NR�YV�Pa����c��qa�n}E <���I��`J�B�j�U����Z��`��`�C�3�i#��($S���uYO�'�k!`�����0���_ر�G#�!(�~�kAT+[���a�l6	��H�׀�Y��a�a��� ���ƽ�<v�1�8C���b(}V��t�[/�_A!�[�(���(6Մ�5�/s�
��U�Z�E�bAB݌��9v띺V��Z���Kd��\�y�� }�e�%�� ���,�^�[�!�	��j dn�B��f�L�m���jFD��P�o�:s�ş����Ҫ���{[Xo1�]��p��2�bG,��(�Ⱦڞ�?�/L�C��PE�&�h�>�ج�N�:}*OQ�C�іe��"u:��5q����U�An���n��"�z��Pc��j���vce�灹�>`ъ��!�(�'P�uJ������$QNNNx��$쫯ܣm�'H)�s!�$u<a�{�;��O��?����o��_w�����_��]�KӚִ�5�[��iMkZӚ�gѮݸᾳ� M�� ��R!��hx����x��W<������@�1Va���0<�����xx�R����B���K� �� K����c}�����ٙ>t=��{�):��������8����J��� ȼ�B���6)�J�A�+} ��1��grz:! �/��0�4# aA�jq�x��i9�H"�-�L�@%�8;�Akj���(,��w��w�00<u�"�����as1[�Co�k��\�� ���^�
���3p�(*�A�d��C���e��+*Y�o8�b|o}���F߿ݚ��I�e�*�pL+1�7�{Cg��>�H��'x���</�C�:��~�!z��)#@X5d�,��˼U�z�C8�(��\/��һ�a�X2��'�0`Amc�C?�/��8��U�6\4��� �XB����Z�X,�3X��	  *��xN�cvճu���+D~n�d�$`Ȯ��6�?tգ�CdNrg�r��咘}�gdBK����W�� � �ݘ�P���ۿl���d f%�[]Տc�����b1#�7>}������� c(�p\w��K�"�?��+�6t9�ag4�5�F�x�^[���\�jɬ�-V�b:K4�@ V�+}-B�=?d89	�ty�ch��ݷ�Cy֎H�Q��cE�:����2`Ѐ�j*1�K5F��|a-\!�G���\A�{�H�H�����r`/�V�or߮9r$`3B�0"a���F���%$HW�a�De6qP�`U�Z�		�~�GB��>�6xl�`�G�S2������
=*8�$Kh/�=�v�EA��֬�*~�	�,�ô���ٺd.� �����{!� �5�	��d 3pL��2�X����U��+�RD{�逊��{]��V #�;�[����$!�[ !�����Ǖ3(c"VvGΚ&�X���� �H$��F�9< 
1@��R!�����xܶ��>+\�C���IP��0e����/~:1&��0��$!��G:W���PDa�B�x���}��xWvvwt�]Қ��UN"
�����V.�\�#�8�j�1e׳��Ms���J,��`�<��wP��s���e�x@�Ab �����E  'gY�k>��IƙBfü܇�{�un�oYT1>s����r�Ǩ^3��Yj絝P��A����v�W 7��g�9�
�랿��d�P��#s��s��֋Ⱦ��~�#p�#췲���u�o�϶�����J�����}�F�98++˙@�ǆ�^���jT�����p��9�ڻc}�9_�f�R	�ײ&6�W\�.%���!PzԤ�:A��e����
�/������O&:>:T����S���0ܯ.�K�ق�� ����*�^���4��4�SR����s�9-�Wr+b�vO�u�r1���eЕnL{��ڎ��2�e(�Y��\�[�gq|N@�gO���tvfĬ^?(4y�՗R��Ʒ��s��o�o۩�P<s������������՛Q���W���kZӚִoqk��5�iMkڟ���Ϥ1�vh �U��2%%����I�aa �R�!�
T������X׶�<����҇�a�����J&��M����U�FV�O�'R��*���s�C�U��'Ǳ�퀀�F?}.��n����3y~z���ޞ��.#2+(�_����nӹ<y�L�����0�9⧪��+�hCfb �2��8�m�dE���.惽�j�ж��<���~�zf�;���lc������İ(��n�X؃;$�r�2�U�����EU�ؐ
�Z�2�! �C�l��)h���կ U(���X�w�������/ e��z�Vz�S�� `	�Y�
���%��#iB�1u���S9�-��Ew�Me^��F��A��^�AvB:N*�@w�X滽�۰�?0`��k����uߠ���� ��n�֕���<??�_6 Z4^O��ܗsD�G����Ep��@��O��䋧=�g�|�3V���4�}������:��O�*��j�X�A3$��ֻ���̼0��!r��F�v��"���AHP�}��K1v(�"Z�@a0��	V;]��h�r�� �^8�3��f�l��������|)k}�R׫Ǎ~�������9�k��5+��%E���x_-�:?VTX� ��!� �����[��qE0��R)B���>��1�;��t]�N�|ắW+���2?a4���,$���A0�ǁ��'x�#�v1���,#'#���Z�Qy�;ڥ��J�fP�f�Ae]�u�2 �P��M[(��oc@?���+�{�vR `*]<Tv�z�Z�!�P��*�����i���k����=���w��+7`YM�v�Ȃ��1�ZN��[��=0�: ��[%K�oX/���^����L�W�u�Z�i �s
�6��dg<������vd���h�e�_��:��S���T{��G���p+���Y" �X��P_��~W	?�fVnh��ګ+�����5An�B�}����
�c.e d��� ���T���2���u\-�_t����9{����e�tt�����k�]*��sa�	+>|a-"Ѡc\`�3"��HX��c`��SI�+���
�*�q�$ɴo��X7�\���a)�|�;])�k����-sh[G1O�;9�ޠT�l�Iv�NYRͯ	�J�3f��O��ͳ-���{ �AGv�.���:�+�����4m'�ZwQgJE�+�\.�s�>B�ߡP�5-b���JW3�	$TBN'�x� �Cͷ/
0�92]��l[om���[�,�ʡz��g�#�Hv�n	{�W�r$lQAR�9	,������+�F�� ����ˡ���ew��c�Z��9:�`�x��}y��套oq~��i���u�� ��V�}Ǻ�n��t���g��3Z>���|��=9;y��a�B�k$�u�,��WMı('��i���s�~�=~�}k0��l=��T~n$CfG�"��}��� ���zfָ�
��(p:;;��q�{����aP��4Y��������X��Xh"9t�4�tm���䗿|���;�"�����_��KEiZӚִ�}[[C�4�iMkZ���-���U�A�`�leY|�_sD�&�,x@[�Z�V���k�A��d:!��l����P��Y�9���6	 xQ�Ѿ�Z�(���2�<�� 9�
�- �X��<W8jI����=�LϏQ�-�����ُ}>,v�=N��s9�J�U�:�>}�����vS�jM�k]�Y:_�Z�@�H؋;��hk�T��`ٲ�6>ķ�L1��!��ުp�qK�#%`��w ��a�d��	B������b���2a�<����<�i�g|��o�.��B�S9�	�� �Q��K�{ɝ�*+V���0G�����7������kf}�pq�X:V0~�"L�{�n�'��ґTi������j��T|��K��)�� ���U/ Xe���P�CF-\4#�@�@��EW�"g�U�|��q�� ��/+7~��1��@��z㪶(!�>(�`^T�������J����c�ϼ0 V�^�2RU� �����:w��µ��>�6�8��z�$�r�SUϪ]�ְ��9"#� ��Ei�4%����s骋Kڰ@]֢M_��b�ڂ/�B O2%Y�Z�ږ�Uۇ5pGk�>�����K�u�H���rk@P����A�h�։�Б	I�2�Χ�m�Z-^Scb��P� �Exr�UQ�dT=9�׶V&L������UDo���td����y��' Zzz�*/t�kHQU���~�Z��k�c��v��¡@��k��JR׀3|�v9��`�i������YAe�P�C�D�B=���_X<�	���JG�y�*���Zs�b8��P��A gF�#�$b���Y`ǅ�J�kf�`�:����p ��^CX2/�$.^�[@�Z�?���7~��t#f� G�`^E�P�sL ��p��N�s��n����˫r�C����Hغ�f��e��|b8X7�ފ���2�5�-���$=iǰ �x�������܆�db��HK�՜�w[7PsPjꅏJS�x�U���	�^,�V�qW �<�$+ʔk�O��lc���� B���3���sv{%rGp/��ׂ�2�z�sXTa�`����^" �!��da�S�OCu�#Z������PDn@S��A��H>(j���Sp�R�yN��W��fB����&���=�cm/�R�΋J�\���Y�����'I�o׏r�&���:����L	�#���=@��
J�k���cK~\:�?�J��\���J=��˻����w�<�����(�bD�pM�}���:�îΡ>��<�l���_f/�?y��/�Tu���ֲ:�a�E�íI�w���h���/�����歗�2��9��<��+�Wq� 		D��|a��$H�����sy��9��I�fs��q=��}����A��O�Ea
�(�������ؘ�z��uPdc���j����˜���a���^��IE���X��7�;�^q/d19���L>:?�珞ȓGO��w�^n�-y�Z-��bJk�'_}-}�xg{%VEU4HӚִ�}�[C�4�iMkZ����^��+��o.��
^۴:j��Ab}pD�@��|FOX���@Ge���bF��,4���F����g|�`ؗ}(?�a#�J���V�
 $��!���ԁ>� <�<�;�"�W�d��BV��'X�A�)��<}�Tf�v����U~ƳG��O>��?��V9V}W:{���G�|�C�\��������r!jk��
�����]/�OP�%�֩H�$R$���Z.�`�%m
�{ʗ��u������Py��D���7�6�d�5@EV��?}}��>��������Fe�t2%���$�d�t�ɰwANE��v1��S �R��#*s`�@�^��-��e��d��r�z���/��Oˋ*]�k���j�5�	ȤI��g�n1�{� S��:����#�r$u`�eB�|g�DeE�g�\���Mh*p�Y�n*��b����&S*8wd<Ѧ =3 pV틤W@&���*g�y��o>� �� �5�������a�z��z���Ne�s;d6�YfY�|˔N�z��z��ba}�
 n��xi��_����ѣm�jOx��F���Qr�A� P���1�!<��ᒹ-��1��q��D<�� �sc� �	��zG툤�h8п��J
 :���� x�� B�Q���dcNKIu�8�)e��
��O�1ېb��g�rd_�	"���]+����)�iA���o���(rs�r�vm]�����^�"��|�E��|d��<�UE�,T��Ah����? �����PF�lӵ�YY�t��ə׃}%6%�?��&�Q�}��Z.�r>8\�	���#�n��&+�s�3Hi� ��Cp:�u�;�7��	̎0�P���ў���],�s�����]K�����[��:b�\����RB�B��xA�1�R;E�Q�"`)����c��@n����O2�9 �M>*�[������l� 0�mE�7K�P�����7K"\S ��)�t]�L��šO�1dz�v,!����AU��cc<�ģ�C�o���«��Ƙc�{�#Hm�*��*|-1������(���<~ڴ�K:�!�UZ�#?V��*����*�8�_���56=tp�:��ޙQ[���ޯj�faj�w�p�c�ϖTyQň
���5��p��\�*�9�](7A��'�0����[nUac���ɱ�T6�B��	���A0��"��ژz�rV�fs�\�I�����T$��/��!����.���s���@�8�$R؊�J��Yxy�q��s�9�<�.yX5��"�kg9�����֯���;Ŗtad;�hM��l�ݾI~��
?j��=88�7�~K~�����_��+W��m*��NKќ{�����+f��4�{��bLݼy�9R;���a?9���>������Ÿ���NE���6��5��?�Hfq�ӹ�qߨ���B��r�{g�	���3`��\��i����F��k済`M8�K7o���I���39}�LNN�X��&g���0GҒ�?�T�b�`q���~�y��?��5�iMkڷ�5HӚִ�5�Ϯ��ų\TX��`���P� k4��>z�܇�h��q��x�Y�W��G|�[�g�������'@��>"@s~~&�Œ��x_�U���Pf�	��Bk} ���JZ�]�&������-�� I�20�rU#B�rM&y��9�@���>7?��/����B>���5x���q�y�X���0-̃���~�YT2�ᒶT����������cşU��
	#?H,V�����%M>(��mw-\Y���l�|�����aq���#����9�����T�<~" ��>�H��ZA�tP�񧮲�|�ǣ!C�Qq�x�!�L�ڡȥ0`)t�!�ΰ"㵇m��O��`�"��^ĵFD�I��{��PZe3�e�

�����T1 ���]��׾Ced��׷bEgI�*;�	�8p�V�\�
ɝ��V��_S=9�diy#-�)hJ}�~pD�~G܄̄0�Yeb:���*�	��!�8�	����9c�%^x����Ri6�P5�:B>崱Y�Hk+,T�#����9x��ߐ���>��`)U��6E�QKh�#�~M��ό���L�/T{W�~pL�U`�T��$/�M&��s��p������`L�2& ~Aц�)�Z�S������Mr
߼��B r_׉uRl=����ˀ�qv$�>���8`Uq-��|Y�z֓�q�����{�ZNI ���a�o�G 9@���̕�Y��{����aeO~���	D�%/���bj=�!	�iT�8����jEm���w¸�z�j�\� �Ҏ����$�-3�	�e�e�]��H�y�Sqy"�� x
� �I�cf6@���@TLVB׼he$JX��V�*8.�? zu��pl8_Te�ߙ�cHuޣ��|bp7��LĚD�6Wum��1�d�]2�5m5�:���I���l=�ʧ,��|���]�@ǇGŋ�1�fh���N*V d뾇����/�Ն��&�V��dz06�Y�B�C�Y�  �E�\X��ȫ���7� s�s[*TO�s�0���4#�nJ �D�I���7)��a�4�q����j��`�@?��+-Ď� ��;{��?���}��ڮ{�Z��缚/]�H� w�� �A����~^�sC4�i�,7م��=�ˉ��߰w�����6�����x��觺�>s`|��T�#$���O���In�H� �Z�
$�ITP�y`8V����I��'��:ߓ
sґ���rA���)@�sᩨ(�
�~��@P(�G�&4!�S�g;�fʷ8W���:�J����X�NH��*��8��uj��S��K�e{�?��PVH [Ҥ&�䭷ޒ������c½���������d"ִ�b�{=��T�]q�����k��s��S�vdwoW:(B��_f�?�Lp��Mgrzr«�S�H�)��(�*�*a��:}������?�-q�.�����&Ś�Ys�nw�Fz����{�}��Z���h)�mi����ͧ���x_�H�|�!gL��T\z޴�5�iM��Ok��5�iMkڟE�ϗ�b@�{��J��U�[�@
"ǇG|ȝ����,�lT���mY�%�
t��X��EPd������e�Zh�>���u@�Q��U2(�e�Jh��i����e�����|��7���+D�5F��`����>x��,�W|��Hn<��+y��K}�;��xF�8�ͺªL}���a�  KoÐ_<PB!�m�4������s=_ `A�}2�Md5�%ɚ6#5��F��3��X�� ���Kn��\��rM?{���\�Q$ϟ?�Ͽ|�l�^o G�We4�x�����?'Љp�/>�T�����k2|&���G��G`�<Kx�pQ��$
�P9	���@^�n	�_7�
A	<�H��]T��)�o�^���jT^��& @�����/�3�w�""/����9Fh�VW��uj��@t�����Aoz�l�[��-��i�ԉ�V����-}Y�״��v̷`$���Tf�����i��b� a��B���a��	T��.�{`#���-^C � VCڂ!W:��dKb&�ji��K1�N	�Ԥ�zF{}��YI%�Q�M*�Ӣ�Kb�T�[mI"�vE���j�� h]�6��rd��@v;8�Q̓��U����)l�R(�r���J��#"f}$�x¿X�ƃ�~�ĲB�@�r'"X���1��Y,�t; �$p��e�1{(�q����2V@$���@�� #��$, P9�+�a�ħ�҈�sS��h��<'�Ǜ"�AϽ����9-�)s�����:�`+�hTf���\?x�s��R�.��r�V��cv@��U�q�v�����Y��s�e�͑WP�VW�~��~)����5�n���a$��	D��7�Ǭ�t�W���z�8��-����/���Z�+�K��M�n]��D?�?�o�n	O-r�X���Z�s�os��u��'��̖ҽ?G�=�?���H.���ѡ����O%�*�8+��+ ق� ���@"�d�LD{�
-��A���Q�t��t��ڰ/�{{����q�F�@���.]�*ļ����x(2�"+@b�я9�nBB��@ �;c��sY)��^��|���.tۯ86���Dሦ�^���_E�j��ϰN@IbI�����	(�+Ia> $z���#j����O�<7�Y����{��fEC�^*A�DaF��s�[UF�Uv���?w��5)��'�'DR�;��*A�t���Y���B���D|#c�ڲ���]�H���e[�:���a��#�R��o�+�V�s7�=m<��g*��?uv��rAp��(.��m�����[���1U���uk�/��r5'���D�S��(s�ߺ^�ִN,*[G���0�p�L��B�Cт2�G��"� #�?�l�?'''\<B�O�ꞽZ���׳�)�R�`�eV^$���Q�bI�>��-	���41�
[�7UFJ�}��>�-�t���O�ʸ��ڂB���r�Z�ÊD�z�υ�ͅ1�}\)��8��������t>�����_���o��4�iMkZӾ��!@�ִ�5�ivU�^U�Xhf�*�5�x���=��� -g���px'���a���g2=���|۬��p���C-`�Ao���٩F}�rx���|1�j��V�wa-���||������gʭ�wego_}`[%*1(�g��U�X�X���H�B��A���!��أ�'8��vj�>�ˀx]�:0���[2����30�U�x��/�M{��O沜έR°Et�L��=ڪ�j��	I\�f�ۗ�7oI�;�0�����'x����c����f�%��8wv�2���@5V�<z,�"�{w��ªU#�Zbz�0����(]&l���I�`�1�ǁL�!y2��A�>�I�${�:
Jgd��ы j2����,� �������GG�L���CNŇ������f>9F�E���� � r����JF L։Y_ы�,Y����Y%�3�1 vl
�M���#$��"T}l�����8X�̀�5�V6�S'���o?��c5Py%SĞ
X�?����c�P����+�(͓>�۞U�R���3�U'$Ċ4wY��v��~/������'g�SZ��S?O�	 O,zΎP.�Tl���ճ{�oղ ��Y�V��u	�ǘܠG0$B�o�Ck���Ā+�9�R� �r����Jߍ���8T	�e�9`�>�@%��
�2)|��\\P����d�.��NQP�	+s�D%��[S�R� �@��_�9��V:t��hq���q�	~?�X���Uo��5��5�g���� T��
�P޶���$�q^p�߲\���Ic����`��5%���S9�0S �e���p�K �cg�kK 9ݰڞ��Pl@�H5EıE�z��o��=�kW�I�i[�9�q��Ζ
#�*�3g���X��=��3�ȭ�3���,p�c�yĥ�YN���`i��c뀸�m�)����0\� ɡfsD�8K9�Y?��*�WԏH"a?���`f�IO�Q����O�=*w����m��c{*2T,;F�!��������{Nyfs���3P?OR�J�k�}k*�=��OaO��$ ��V;2[G���F����A`���PQR���=��ps�*2)]фɪ�6��H$�u�8CÑ�{)�8efVR��s�^�ш6�^X2O&IfqY�#s}Z��.pO���>uX����H�>&t�+�& |g�I@�9"9����s�C��zFT����;�@u�F���`M�>XZ�l�0\�9�9�3��Taɱ��LU��]�m�S��ᶔK����W�|�I>��R����Թh8����Q�U�a5�nm���J�Zqo �Wn�*E�TOs���}P�}�HpԤǿp�d�#>��-�����/��j�u.�^�9��"�~|�� ��?�,tH:�Eג�J�����FL�̼�8b~�b�T��g�6T/ ��Ҍ_f�Hu�-y�R�xk�Ġ)�E붌�zQh,�-'$��<�ƐZYi�R�$����gSKkA�?Y.g�>�3@'�{�͌�g�#S'"�j�y������}�^��B?��/)MkZӚִook��5�iMkڟ���^��w_��`$�ѐlx��Qm]z�Xz 
r���'|�:{�����-]�f�U�#�q����>���

��A)-�!xT$��#q�+�~��Ge2 ��.�P����	����p]�V:}V�o��F����Ǵ�X�o�y��f`D$��J�UJ�B_	���ڮ�"@<�= [T��/� @y�@�?]�a��X �ux.�w�ܪ��y-4�OY��}������"ɒ�0�vL z5O����1,~0�݃��8~dfTf���N@�|��W�!�����n�J�u�����A{��sĂ��ã]}��]��P�ݻ'?�B�O&�FVQG1=�'S��?>�e2B��q��:��Q�$��������V �*=�\���%�;�sTLS���t�������"��3�Ѩ�� EV⇲Ym�ҾG���������w ���K� ,
�1�����
@���.����!�1�O��M$� !��39=yN���|�J�Aְ���2��m�X�҈�+��������p�+ � 6"h��Fm��)Ӓ�� �����B��m5@j��%A�V?&m�*Y�ZJ&QO���iBX)3l�gZPZ�4kE�H,�����!�oʤ�������d��]h8�_�~�ǻ��1���#Q���B~EW�&��k=���ܙA��"൰��h���c��xGv��i��f( n���7>Ǡ���6k���^�˷n����W���ծU���+��\��v���`-�sM�����~D��j2�D�H����L��6� ��WPX�O:��f��u�o�E��Kw8��#�h���%�Kt�C�.��銕޽�B�4"��{�ot�[��>y5����5�I�sj����=�~CV���xꬉ�` ���bm���u4����w��
��'q�5 &0SQ��uW�׽�`w�yDXK�c�єJ�m`�MSX�_-oCd��I���1O1rW�@; yZ�����¢�9�K�7��1��ֹ��3�� ��u����Uؗ��A�r/�^0����
*��xc��pG2���lb�>Ò��5���Fǈ�B�7-���c��M�Y�3dr!�ABJϪ��Mu��ܣZBׂ"/:��£�rjN�*����ՠ�J�%1� 8B��#?"�+\�T� ug�����͖ǁ9���{��Ҿ.q�PY�	�W���Y�l�tO�=$)ֺMe���W�>{���:��f�����7�1+�>�g�3B�K�_�NSQgk����.oZT�N���y>(2 ��A� ��ve:?3kr�tD�0�a�%�9�>U ��/dv~.ɷ�vq X�L��^����'Ʉ�$�����	�^o�}��x�j�� p¨M˲,�H�m���+�_A���(��C`y1�GH|8�Hߩ��\* ��P��Op�5�w�Plձ�#��V�,k2V�|�KS^ �$p6oP	�S�c �.�~I#���=�h�c��r6g�L��{]�a$C�*u�\�Z�1��$?��#�Y���F��׊�T �����.��B������:(dO�g�?b|Т��SȮ[�� ��͊]6$�0WV��֯9�[�����ÏXt�{1.�iaFZ�5�*$��5��0�u���˖, ���F�Ԗ+(,a}��7+Qh��]r�0v�߀�-˶eʹ�3�_�w���x��$bWxo��M�yf
��&�t\,�:�+���>\ǥ�S�{B��U�b���u(b�|�o��J����]�o�Ҵ�5�iM���� iZӚִ��Y6Z(��}�X�mdYx0�}���h^�QĊ�R���Uzw�i �?������T�� �Z-I"�J�����A�;���������{��յ'6 l�	�D�����K�P]�;��QM��f?R�A\�WW�{=v<�&Vy`����0�.����.�_=7|6 �����,,C�:lX���!z�X�$�%��K���m��CfٴU��A����₲�x{}8���m�&�q�ȑ{�g�8r�eb!��.&t90�HnG��K-t�g�06��l��oAZu; ֬�����P28^�u�7�Lp� ��6r��kq��[ХV=\.M��?�sq�ER���\���
�Z<?=����@�Td���5{�}H���2/v��A�/��r6%	� U�PF%ȴ���prX�68.���tf�� MB;]Z���G�*p�ĬX/�ځ�#f��[FE�p0���=���ql`���ϙ͓ \�Px 5��@����J���h�ԓ�p ,�t��Z<  KT��ic�9��3��mI��"� `�/_ϵU��|���j�,�+�78N�|��薋J��6��W�K���.���j�>���r����P��Rf�(���S��fGĹ����w�k #�[�O'��H�7�	Q�nlT$h�8���0�H��w%�U�8˕:ȼC�
Dl���(�<f!�a��N�씴���T� <KV�S���")�%ASS��P��NV�2��	������2P�(�5�x,;�n����~��c���y�8��B�`���s�~ y�d	�j����"��H$0##q�m#�,�,X���tjE W 2r�\�o
"s��W��C#m���3�h�`l�׶T纎�)߁�[b!æ�'�@m�7�d�� �cl��M9Y1����#^"��b�'P̾��E�D�cg�j1O$nH��r;"O�:�4Cx9-�p��rd����F�8�2�)��b{���k���;��Jaй�jy������e7i��MW#��/y-7���b�_���W����������f����O���BUh�R�
��"M�ʓ:��r���1����2���{
���@$��P�I�TN%�������E�������	��dĊ9� �"���ދ�����Z�������^�\���̲(���s'9mA��R��"�}>u���ӷ!ߥ)�F�(m���Xq�>}���YFv�"������Fm_Uu���q����ا}gn�?���y�,�r�������S-K�޾)�B��b^�j�$��ր��"���5�����ZEc?���#Bb{I���#u��S��� �o�JE�d���\@h�, �LI�lIa3��ɗ_~-�Ŋ�<�q����9�,����r��S��X.��7z����9J՟����>l�\���݋b�A�b �?��r�!Uۧ���ync��|���z2gvY!�]��?���u %Q$��6Xʥ�Z�5����X+�X�WUX~Tx��ִ�5�i��� MkZӚִ?y;GP��*�ΟM� H���ҬPM��x4�j5�r�6�0Q�π�����2t���c6H���ٌ�ǽ�=9::��`$=�H��OI^���P��*=�uVH�9�V߇�\dL�B?p���������|ΰ_{x���A�?��-�K�ZW������yz~��&�7<���w�"'ⲏ2��$rg���\��8��O�+�?� T"���k�Z�(@i �s�NQ��ҷ �_���Q�G{}���C�7Z��β��q�v.��6#���� h�j��Y�l#�� ����pO6)�. ��� ��!��;<�����B�����=g�au�6�R�j{��P��+VdzT��`+ ��W�ɳSy��S=ޜ`�G�LX�$���2>ԃ����}V�����M&�g�{ � �:7z�����E��ѣ�)�sM�
�<�M�K�P}�3 V�G����qn$�2�����Z��z��MT�K�@i��v�#,tdd�צl?�2gI��@@�
�;>�L� �*yΛ$�L���1r���T P6��@��r���|µc��޲�l��a�.H�vl�2_�Z�Ǟ��#㵲�0P��oiH�lA@� �Ś@�� �P٫���$�����$��'6o�9e|!l:�X�<�/T�י'D� ���B���q��Ti���p0�p���w*c��5��q��7�j�x�XV�L��	��S!��) >A~FJ�u1[J��-\���\��Ҕ,^�Oac���P��rBp�@��zm*����Bz{��,��,�*S����C[�<���ZT�e�������-*�P��� {����A�59{&3�������@#Hp�x�pe(;m�č���3�B/�B������<�:�S����ia��&S�-��/a���h`�M����^���%65
��za�պ�����=�=G_���j=����stl=Kt�t�LO�4$1�E_��;��x�H��Y����%@�j"���~��O9����6�C�"��ֶ���%Tg��'�^���
�+W��6	��g��^��O��yF"PWD�I����Y�+�?�� !+��n��^��Jh�3�Ϟ�Nu���#׫������7�s���� 1@Fz �����ܿ`}�� T�$ޅ�{z�\�>{$��8�N���ýTpQ�6L-Ǜ�%MTF�-uܞ��ڭ��L���}�kr'�j{��q-�|�_��^?<�W_�o=�{���c p�\��'+��/+H���\�{(���Z��\(�.���P+�rt���@�SN�:��s��D�m��?�^2���5��5�u5Ym� �]��֚��a�M�$��$��[�ke֪	-4 @@Cw��~˼�o~���5��HH*Ւ{f���1;�FD�JH�FM�IVfFx�_�~ݯ�13�A܋@@E��Qbgӄ���q�����=�£�t^�7%���/�<�����w�����LQ�PaQP�i��O�w�,;#n����O?�gϟR�rlX ���^>Ϩ�}��<����ς�'��l�Ҟ��}�c8X��`>���*d�:��n�0�yx��=[��C^�ҟ��T��c�3Ա�b
�SHHSm��36�@��y1XI���dm	F����߇V����=���� ���M<���0��T���33��l���[1y��kZӚִ��u�� iZӚִ�}+Zg�/�k���O�2�  F b[q*;�����raOi,|��@���K�>����ە{G{��J�p�ŭ� ��ٳ����s\�ա�K��:V��~`{� �v`����CEITD��P�W�Y�l���TV�ٚ �A����D��΅Y�@�@k�������壏>�}|�R��.n-_��N����	T�ב������a1:��P��h��������`h��+y���5 � ��d�1˵+�{^�B� ���*�Ͳ� t�Q����h�]J	�!$]��Cf	+P��?���t���,��� oPYL���d�~��H�Z3wN�m���X,	t�A&�O�<��(�h���W��P�I_iP����o�t�nx���{Ƴ�,��L	>��������n)��U�%��?5���� o%�{��<yL���q`���R��Z��e �t���^5��:�Y�9���D)����D�
{�j1�˫s��<g�6l��H]ѶV �P�
p����� '�1�sg9%�3]Q!��g̓�k��*�#�AP7���㋳S���zy�〕���%V��uY-t;%����б/q��@`;c���$3���m9jz�����D:��w�$�:_,�{��f>��`qy ��b��&S�ֳ��9?V�O��K���W�5Uyڇ �X2�'5�7T-8�4��|.P;�P(Ib\�_ȧO� �^� ��9-��7T�b%2+7��
��H^<{*�/_2�������3T�`.��yJ��|��W ]>��vo�g/�d����D�y!G��:�f$��9�8:�F`]_����c b��)A�v/f�A�l2i�/�8������s���Od4�&��k�����t15k6[i���F4���{�۸�����D�z�T�!`�<�G(b�E��:�1u�_zfdr�#����5���F��E���{�e-I+&p~qy*/O�r�n빢?�έC�6 �������N;#pX������s�#�{{]�ǖ:�[��{;zޮ	�#S�	I�:l�}zs`�����ޗ@�,���<0p�
2#�Jz:�R��ryq*ϟ}B��Ū��NǏ�%�>�+���4Z�5{�_�$�/
Y�ܱX�e��A��dH�e�F���Wo�:��� ɴҹ{�s�b1���py #ϥY��>-TP�$up�{���K*a���{d���Y,`��z��(�#��<��/>�����s�-漠�y-���kI:�����_ȳ矓�ju;�����=c8�-��`6����bs=��\��|���B�	@�r^p��z�$c~Y����F�i�����]��|�r��\3��5�=��o�}(���Hk��q\�J�9��2]�bq3A��r�0 ����������*��nDH�p�^�Sx{(L1u,��%g�ff�=?ڮ�'i
e��父cA��^t��*���ͩ�%��
��DH @l�-*��� ~��s1�+�t��s��r���V�� *R�������������~�[γ�'�ZD�I�bAr�B��t
��J�G�I=��A&G��$R1ޠ$��|���T�2�ޗ�_]v���<��6���?�dx,������
��M�@�B��m��ŵ���1w�oj�*V@!�%�����,��^��L,_�t%��m�bXv�����U'x��bo�Ҋ��k�4�iMkZ����� iZӚִ�}+��� �n7��.䗕W�f�����u���t�JѼ\�Z.�r��G���p;�`ظ\�>�����
<�A����Ө�$�X|m�i�m�ju|��� �����.� 8 �X�!�@ٙ�oR�"�j<be�U.[šy��\�>�L~��ȧO�����}4�!��pjTy2t�6� ,���`]��΁ꢠM��3J���H��9-	�-��ӏ���q`�����T,rQ����Ҭ����$�0԰�G�ތ\8�:����Ǭ�ZŃ�HK;6�,`W������+�Z��>prie���y��AWX�  "�� X��u?���������5�f@&���v�P���#W��ĩ)R�ت��z�e�`��XQ�@�	o(
���$�QjV��ģ(r���o�^�8U1� �$η�1tvr�hwؓ�G���-�:8/8���X�mX�X�����G8�0J`dE��v2�ٞOo��SI�=�.}-y� ܃Xb���{Q�;�N��L���՗S�/�ٳ�	�����K�'��D��k�0���!Ɗ���9|��39}�LzM������;�;<��H����T"3��^>�\�~��)gȹ^��� )ՐP�����L�:�m2]���?g.P��c�.�nJ�����	�a��%µ�B?�����E_���k�?�!�2���8`�~!��B���F7���'�p|u;)�]�}d]P�?��"��2�!�j)�P&<��Si�ؠ��.8~R��w�zru}�j��vh�
<�W�����~��m�P�Y��u�עr ��.7BX?j���
�������~CЩs��	*�����ɍ^� b�0��؀z���������oC⨫��%J
����[W�+$sj���|a�>;}!�|�����J�>Z2��IgУ�y)��H??6d�s��xzMRk3�<���9#y�㺠�GG$T�@�P�c*�^F��OX��k����C��BR�7:W�G�rs�R�/^��yZ�<ć���MÒ���d���`��驜���6.��r$�x|l�^ajFS5��]��O����TǱ���>ڱ^cu���	�S��"�Z蹎-�ʄg��A~��_܅*���tDP���� �#��9G�\_���iS1�Sق��r<Ҭ%7�$�)�' �S��^ʵα�@.���$"��7��H���b5�}ji?�̋ ���^���^+��_�nG%��v
7[�����:�O>�-�R�ڧ�|E�xY::�2����b\@_��ù��k�QG�5��u�cnXs���{������V��J�m���"�f:w�@Y��TY.�@�s�z��$�⏴%C��z݄'��b!�P��Oj:���z͕�Px���������d��F}�����=Wbv���s��<��1G�Й��x�q#�@V�^��T�X�=�(�y�����#�ƽ����7�6��q������ 9��z���wѿd��ʭ]K���[ N��1���sB	K'�������5"��G����6�u��$ @��zreys��l���5o��<z��ۢ��4�V�z��ܧs���ɏ��{��2�NMi��$�p��1����W��usyE�&�A�;M�[˰�CEkY�f[Y�{+i�yʑ5��՝p�ó|����*�����4�G}�eQ50�u��C����5��޴�5�iM���iMkZӚ�oӫ�{�CMQ[XuU���@ ��NW^�.��,P�G�0���Z�ee4�m!p!� �R.�$h�"��P���fF��r	��`�q h5�AQ�H��{em�=��Y����gӢH���ͯ%���,*S6d����1�X���l>���[��Zn�2{���O�!x�����'����zPK'*��<_Y�
*u����D�vPP� ���'2�&�>��.��y,��"��������g��Efm�G��c��
��m��َ����� ��Ap0=�3�0��;m��ܸ�4Z��G�v�̐H_�r������I?��Qy����u��{X� 	��~��{8�5���A ��T��YF�	?gwO�	,�:�j6����;�����qF���U� &� |�x����>�����XA�;�q%���usmӿ�lGbͱTV$.Jz�z>�f熜
�o#��Vk+3 ��_��vK?d0���Ūrk���m!;NͬZϤ-�_�fl��+$�z|�� /�,����uL��
�G�*��`���,[��vg�����Ƭ:P��~Kiz2_��Yx�L��A5q+���kepc'�;.�=�)��H���QI��͢�Z�P,�X���I3�F��T���s�*��`�@m�*�v�.��a]pU�T"T����@��EL�s�H�
�$67��s� ����*�Wy��A�% �2��t�k,!�	�%�u�=�0�,��PͩĠEȭ��l0?�����oPK$i���l���a��S�ݺ�*ڦ,�>��� ��Q@eQ���q����y@ <��b�q�-+��#4W ޠJ[)-� ��	ܛ�0����W��킬\W <z.���j+���3s΍x/H 仗b�\��>=?���'����DB�웈��x9���vf���h���
�	-�0�1��^9^���1���T�Mi�})I����9�q����y �;m�s�C�!�dc�X+@`�H��3�T�� a�D�^V��w�9�c��@��y���y�@P��H�ܩ�95y��Vy������H�r0�y�P�@��t�]�-���_P�0�;���ְ222
��k>#��~�u��֊�so��k�>����t<�f�D+;��3��}��1RJ+�ۼ�Pj}�h'��
�4f�ۃ��*T�B�b:Fփp�\�˟+��]����~�s�ɨ�p=�:�g:�e�iA
�K��*��:��X<'��s�)����ݐ��p�m�E�Gm�>��-%˭[d�)'����k��|����w�`�-G�vH�YÝ��c�Ϛ:5����Ȍ Bejm�(�@�|J��Z=?����)"��
4��*�W�Apۼf�fT��s2��ǞQD�I��AA��ϴ������K����{YXP�k��#k;��V	l�V���;���kPDb̂����d}���7O�<�7�x��W�/��� �W<~�Y!������)��|+wwy֐�g�N�C��4P.���O<����gtmF�֊*Xf�Y�BR�L�9.�]���j)ސ%d��}#ױ�ǎ>!���Q�4�iMk�_sk��5�iMkڷ�y�8��]V�V����z��F��ё{&�2Oe��` ��ɜ8,���vh�D�6:�0�M����� ��GT
H��*X=J@$7�a pW�$["V�-ԏ�/��AT���o��ܜ]ʛo�!G���*%E�.�O�>�'��.�jet}����Uյ�z� 0����t��"����aM;�����  T���b/�R��L�n�rzzJ�
�r��u��Aׂ�	�Wp*h��
X2a|z>�m~$O�����]lw>W$nr�X0����r8��CS.n���mY�?�s�M���d�[_��A��������2`��H �Z�*m�Vs��R�L���W��i��
������C�ł���~�J彽ZU D�"���w�����<����+3ac�l��4{0f��"'�B `"��rS!��}b��_�����M����X�˪�X���ߕ��#V��A����������~^�ա�����|:��sE�>�Mݲd�z*�y�M����<���z��p/8�uA��ɫ�Daֳ
g������޻����>����8�Dv���h�#P����1�~���;��~3�FX�
���܊���r��t�� ��,��	��z�!���'/x���k#���~�#y��������,�?���	�~�͈�w������|��?����K�N@�����*�:�\Vz��0z+c���y��ߣ�_��$2wK����=3}�~N�����ѣG��?��?8�u;.����y�}����B�Q	k ̏����&w��1�$S54_�:�ã{$J�*W$�PՋ���.���@�voo��1rz�]=��۰)b�yMW�wgO~�}u��g�h'�9�6��K���u>]"�*"�;"��㜾�����y���t7�	���[������L��+q��-#ណ����Z-�`أ��g���X����Z�����\�$=y�cR���}G+^�/ ���d�+�
'ڎ����>����x�t�%�ʋ������ǭ*]+�po�yz���������3��װӍ<|��ټG�^�� ���7?���?�E#�W�G��\?o(��=^������-��ػz�b��8=��f��f?���7u<�Б��s�V:n��)���~��u�ۅEf��%���ww����qf�+h�����ν�c���I����>	e���}����QE_C g�;>s�~�C>�굇����l�^{����Wȧ��# ���#����#��0��k����<���Kɂ�
��ͷަ�OW^�[F��o(Y{z��=����X|�j�O�a�j����B�y���E�ׇ� ��������Y��Q�ZA
��(6s���sPMU�'D�'��§1Gu=�	@x��k�ȱ�E��#(-_����R�ۜZ��۸_�1T(,��h;��E��l���ߛǦ�ڈnH�=<{��O=��96��;V~���B*��܉�d�yC6�^���d@RǊx�  �!���eT���g���
�a�}	=P�eI�߹I�Z���D~�cF <������+}F��q�~��vG�f鼶p�T�~��ʌ��l�^�8�u��^���I�,�=�Av�ca�����tPO� ��>xNʍ�&qUnm�8m}����3Jų���qqK�/���~�~u���}���X�Ki(��5�iM����iMkZӚ��h+�D�30���͒��pd%1�-S�1�\������J��	�M�3�����D��yww�u�3���+@�$�����R�E	~��B����UTHf�x��[����WVՉ0P���-X�"���܁�
2v"��im^���ta���: �UNՊ�����󬨮�z��뛱�i ���s���Y�{px$��4?99�m����frq~E0d0�!���
Xm�jHT`ÃJ�Vfv[�0Ǿ �/�����r$/_����+}_[���.r;R�9���K;{������wޑ��{O�����Ī�3G(��j�41K2��N�H�v�k
'C��haA�j��Q����ʒ�9 k�ڲe̿|�h�Q��}���ˀ���!*�O>��<�]T�&1��I !PWVa��mU���X�����QQKT4#�`gwHR�� � x�b���ܽ�#�S�ד��~[�����ʛo���7�(�B���Ъ��F���z�p�Ú�A�-��ˏ?�P���	tƑbVH�KƓ���Xv���<�ֺz]����˃���C��A�Q�*ו�G��"��F:V�8#�V �F���?�����{t�j,*��!���Y��*�V���[�!��Ʈ��� Sj 9l�t?v���� �S��h�W�ß��C��~DOy3�e(4�����[I����l{��c�����J �5��ƻ���J�AMf[����w�}�����pnAjN�s�N���O�������������^�����H��`8\�7�� �w�	�O�������{�}�|Lb�s��\����=ٽw�U�PI���ܨ�������y���ia���#%-�f���~��k�N�J�sӀ�/³���wޖ��]���W��AF�`�@���]�:7B	���C��/�^V?^��L���N��̷�h��C�B�H�*ǋ��
�� j�[�x:8:���6@�v@X�����G��޻ҁ*J�&�M5�k��+��qR�� �{��=��'$QA�#�h�;��"y�����1[�<��g-[������I��{+'z�Œ!��<&��9��*1���辎��[o}�s�% �=c��c�c51���s����?g�<6�u�����rO������+)Y���������?�I%8���S�7j?#�
D>�� �e:��~��5���O�����4�1�F��Sw	`3W
�d�Cq?�����P�>�wmުc�2Gz��B$8�\K��;<����/�z���^: x��-AПG���&���j�s���~"O�zIb��)m�`���������s��D̃��c�?������$q�2kȈ�OG���_�������X�2����yH%^��!�k�2*~��dl�$���|��hU`ˬ��̂��2`֖����7X�eh��e+5�>,���=N\-�&�}1�2���s BB&�ݓM�cY[v(NE+�2�a�9�E�սm*_p��Y�=Ϟ���(-�#�
�}���(������x甇'�l1 _��H��-7���%s�h}�9yJ�62'<���'�ڼ�y'�%��:�S�<�º�ǚCp���M=2��Y���ez^A�������&EĳHb^#}惕)��Q�����BX���T�]ݴ�����n��O�}�ɂ��rQR��9
���b�	9(w�?-t����J���~JҼ�sH�˘�%)��B&�ku�,%�k�MkZӚִ��!@�ִ�5�iߚ�-bPj)�~_Ee�i[5{�� ��7�#�7r~>�)��J.ϯ��٩LiC!�I;2*F� v�gg/���<y��� �F��fms3��
vgg�� � <bq8�XE~U�E��U��Ѐw���+�� t(�=% �kwH p���"kQ�w����?<��?,;`U��j��k� N�օ[Q�P�wvvn�ȨT�"�܌�O.����/ߗ���߲����J��__� ��c줙�|�
J� J�:7�r���wrE�x�<��5A��b�t�jSe��樨N�8?�6� 0� D�������GX;�� �4dg�t:��VJr#�,�����֨�gT(��
�,^ ��;PM �"jC�P@�E�f�K`)P���sI �a@D�i�bݿ�x D��,u�Gӑe� �]?�B�y<�ѧU����#���^��=p���+�# o�:#=ϓ�1�Pώ�bF���Zv�F�`��{҉:$��H�¨��������ȇ�RG�����jM�TLE�\�uT��	<�/S(t�?x�X�V�
�"7���c�>�\:(u~~E�	��^;����|}MՍ�x�ڧ"i��@�xa�A� &Q�� ����C��ݳ��G�����@���2/x�XQ���؃�a�Gb1'�Zxn�ˡ��sZ� �������Cx,@%*(m�7:r  �쾅� \m)�նm��Tu-��5�Cm��l����yQK�D��P)!ק�̙E�O �\��-s*��\?0P6����jjTb�B��=��TBl�Z��;ߗ�==T+�����+����df�G�\��?�Gq[4��C��G_�TL�m���;_q��{}y���IY�67��[�$A��;_�Xh0��,uw�{�ӿ�;���~���$&(eT��똻H�i��{�������c@��R�Y ]NFf�G�R�}b�1(��ҁ
�;o�%���n
����f�"@{	^�EK.����P��������LX8M���MAE�a�Ȏ�o}�]y뭷�:��3��^1�q@����ȓ�l�2m��}>���������@�Ȭ	r\T��S��a�Js(Gސ�t\��=��>���,����4��g�U�9�� �~��{���@V�ӾǸ.9�����f22�慜����K���58��Z,	�[1�Ah�e֚z�W5��'o���I2�V�n+����|5�~��c��(X�����1�s��!1U<�1��)�������}��w���חET��&UJB	�&�EPG��i�c�G?�Urq�mq��=�[�#XM���^G�|���|��'�ˀr�OG��@�Ph����DLmj �$��<���6��NU�%�Ls��h �3���h�a=�ǲ�{���ܲ�*�*
!��zM|�k�+��!D�-l��郑^ӕٷ�e��@ܙ"��(�w����Ѡ?��E����1䜘��cNR��g�jn�9b�?����W_���y�G����-ޏ��ϛW��$kƳ�ݟ��3XVA�a�X�>kt�9�X:����Ծq'��굨
�.�����-�n�7���_=���9�<�`�SO2�~�E)�g�/ .poE�D[����}��x����:�*ԏ��o�k�>�vO�-��Bvє�/��*�~w�����Lϑ��n�����B���q�������y����-�`w;3�\>�z�V�]#�9b	���s`EkUUӚִ�5�5HӚִ�5�[�9�aM�/VJ���ԁ.��j��q[�ʽ�C99�
Y b�~�c�M�)�@[���@̪L.�Sz��D�z��⒋KTB�8T;�t=�{ą��p����2a��1JM��ﰁh1�ؔ��3�z�x\.o����	*�
���Z HTء���W� `x��Jƺ e��d�*_�IP�}b%��B��T�b�D�v̂
����OY��	�XŰف�բ=]d�="�b����I�0�H;f!<�a� 0~���B^�X���.G\0���ʁ����>�_���� ,h=9I��dTz
l����s
��0-�P�
�* 4w"V�� �e�V�w�Yq+�`=�e�≍HR�[X!Ybh:��Ea���~o���:��y�0��_�sߨ0�c�nd6��xP������:���i�"�yg(����ת�	��e�s\�5{:&�H��9�z�=���|��z*����Ψ�쎈�u�B�QV�����������j�`�d���-Y9��� b�|�J����Q����e�N�a��vA`���Z�Y0���? �elբP@��HV�@�Z.�K�k}2��Ŋ�II�����BV��Q
���^�k,����V�&��E�������; �8Te���1�@�������} �u3n�p �)�x#;�אقް�,�����{6��^@�b�sZ�^mD�[��~�qm�k�_dV�֮�'49�'�<�ڒ`���ul8/9�Z�Mݒ����yd^��W~���{)ò���`�k_��
Er����"�y��'"�=#I���Ǣ4�F�B�g 7w���s:����	�:�"Q�]��t��L]�k�Jy-b���UQ龖��v�Ok������EI�L�Ņk���`e�E�j���!��:f+��%�2O:b�W�gH��<>�k�H`�#<ͬ@O=�Z�)��1WP�e�^wڪ���Nx�P�VK� �, S�� y?���d����uL��V��ny:�ǯ�P�/FV�fqE2˳pM�}���w�W�lc�%C?1�ɪ��	xn�u�	��f�Wm�x�a>U>nՄ��g�{�W%�(*{��=-���?@v���s=�I�$�h�5�$y=�?u����[]�`�m%�\�7������s���i�f-^�(���"��\a�A��u����ڿ��Z����-�^)�3��{X֡����0anw�-���~�n�O��aŉ�0ִ���9Yhf�d�9X7��9�UY>cF~mTn)�+����d2�sK��2���D �q�q����|V:	�߬��S�ۃB*�۳�>�ύi��{,�pLؿ��|*/^�����܁���`W_�e?tVs�{��=�YA��C�>KÆd�1��+r{ҁ��u��3�t2��g�$����۾�L��L�ܿ�
h���?ˋ���I��H(��9�#-���hL����K~&�9�w2�>�f��$��kYE/Oϩ�>�Y>���p���ܻ�;ؑ�3 �����?��>}��|1������x�&��ִ�5�iݭ!@�ִ�5�i�f��� ��X���[�8@+]e"�x��ɪ0$��IYuP�ƣǏ���ZN�$Ϲp�"V����t���i���\`�2��� �P1x31��>ɍ���m���I�s.�#V\��С��bfA� U�|m�RzH9�i�g^兑%�z�E�5���!�G&S�� e 5�@e�U��4�\�^�P��������J�Q�A�.@`tx���� /ԝ����tI[T���0�Հ-�[e��Y�ɪ�Ewu="ؕ�v�'Ū�)��Y2YR��Ћ �\ж�m ��q��h�(Yh���H���N+��5�*_�! �s� �����P]�\����C���5�϶X�`�܄��-�n�V|�w �^����D?�,�ɒvC9�uk��F�f��蘝��ł�` 1 �\_!G��]�%Ѿ��E�<�R{���a�� �(\��~� �����)L�
��+E���]Y�0@�� >��G����0�4h��1��P^S`X����B {U��Сj>r���,X]���� C�% .3�v���y'�/�YB�$F>����>l�bW�`\�@�A�0��y1�c�Dm��a쎻%�� ,Sڪı�񚽍!����=Q��D��E]�A�І)6�<6�t+��w�˨��j �^ա�NlA��WO Pc��q�����č�ɚ@����ŕ'��ϱ���	�f�P_��! ;i���u	0��el`�qZ��a��6��4�|�##��
��
��DEL�#� ���
��pH2��q�O ��d̕Ҡ��S���l��9U?UbD]�jt��*��1˂���s���5�]d���"+�l<R����I7��_P�!���9���miIؖ�p��]�����ˏ$Ub����]�����ʕkȈ��\�>���<�;�iv_f�<@��fB�;k��w��@=b>���M��GJ���y�]��|+�����fP
A���%
yT
sw��02��v��L�>�*hyT���ʑ׈a��bvEŌ  �K��(r+��U4��E]�Nr�0x/LL�ql�*��ח�(�ad�C[b���$���-���9(K��T9~��~����C^WF�@��m�u$�@�?W�Z	a�h�+laց�b;�Hڏ//�s1��_�A��3�G���� ����c&T�,hof�	����'$���ACi���b�$�۫ж�d�/8,�]�I @*>�6�.�
���l>����z}fəc� Cd�x#Ŋc����O[T�sKb�B���d�X�0}M����}Џ���_�Z��|&�N��<�{]�?��3�P���]��a�H���^��q���F?M��A��9��`8���Ք�kxZ۳ɰ-����q�A�g��������y��2I�氤E+ȋ�̈́�5�4ۭ��h�g1ؘ�X�쉂'XP�u����͔�����9�Z<8�e���I�}��lX�ȇ*���u[V�2[��'h^iZӚִ��5�� iZӚִ�}k���F�p@���ť.��Y-���Ӌ�29z�-�BJ�X5�2�o�����g����R�1���$8�1�|�L� �N��E��]�]^^H^��;�(x�\M������\ZP-lPИa0�ݢ�~Ks��b���V$�� V�V)�����bVLs]^�n���j��\�X2��X�k�r��س�Z�n���,��E�|���]X�������pO>��m�گ�ON����ݧ��lk�KX)LT�\]��Nr�۴�PXz�(��ęΙ� K��h���]8(��};P��w8��t��B��z�"�&,���Ɛ�܃����m�`�e�n������TP�l�F�Z���_ c��X�
0ف�N��\��rq&�����2�������������Eʼ�P'���-J^,	�[��{��3�>� �ﰛB~Ǝ�>��j������3���E6,��h� 'C�;�-�JsT%����'�� x;pG�Ϊ��7U '����W7N�� !Q��ܪ��(veR�2�ω��rˤڳ
DL�V@�{ ��O�6gU��o�T@b sB𸖴�0�8��i�E��� .���
��P1�-
U��FI���7�/�8O�t�} �1�Q}����F
�<�x�{���cf�aN2�.���bJ�-b�*�-\���U��BE�5oI&$�k#�"u�LΥ��*�K*JMl�x�� 	y3���Q9:>�d�y��}o���)A��u��7��H��s�IJ�u<�M�D�k��De����28��J\X�.��kx�m�P�����ϝ���z$�`dn%�k(��D�	H'�/��?6o0*� $.�تL�D""��]�	I�� �Rz�?	Z�U�䂪�C�:7asU�����%ٕ��U�W>dl�u�~�o>�����,�`�5Օ��ĕo����X�	�o���F��a��DWe޳NCs��%�ߦ2ҶvB��y��}���K�m����$i�@r��A����hA�Q'2�DXI�V������������kGLm��e6�eACm�3�a'>kL�@��UײV�P��z4 �BՕ��@΅>��xMf�]V�^�9D

��m�M���՜Dz~Q�g��+N�tz 9�B�a���J>KM��s�&�7	��ܛi���[yw�$��u�qiw��6�K��7�,���Y]FQ���3͘�`U��'�H-����ɨ�D�V)��Z	�K�/[���r;,�_ɂ��*a�	�X	�xN�3������]��Ү��m���5:z3͑�QE�l 򠆝�Pp1�Z��c��s�<K�E:���7��$P�������kfY`�3[�$-�L��4����v�:�Z�gJbZX.�9�
0���쯐�S�j>G�_8̔�Nd��H������]��v���%�9(��%�!P���t�9#��DiqŸ�;r|�H���x��o�<x}u.MkZӚִ�X�!@�ִ�5�i��2��N�]R����=أ7�l>�8��f����|]��7`�**h˩�^�I�+R,��.�����zǂ����U�u-��� ����2(����ǒu,��(6��^�O"�օ��e^Ж�8,��J�l�Bx$���տ�X�
ۡ	T��Lg��*����B�}��E½��g'���
�Z>9=�Ϟ>����T%�"�eMk
�*��tQ�IT��Y%��zl��˛k�9���ш`,�z�>�  	2�u�:��n��}�}��B�i 7I���@.v�2�?���_-���X�
Y�ͷ�'��Z �	�d����όvP�{��K,���}kE����u�;fJx�������=�$T'VU���S�,Nj��rP&��t�:����|`�r�6k�9�1��$_��rα���m (@�4����~��ɐ����N��׻;C틈J%�;�� J���d�s���e@�A��Y�����)&�n�	��Pm�PfߦF
�N[P	�x1���4�#�b�udj�d�Rd�W(h�^в'�ZE ��e�v6��cд#6�$"�=����I"W��a��-U�v1P��H�O~ �m#���� ���Zr�@��g��u6��؀���k�[fc�#5�G6c��`UE��u�����͡�7�ք]@��[JV��V-�1Z�W$j�
�12��*��(���kp��%��Eɺ?�SN�Ĵ�ɜڪ�����Ʈ��mWe�Aԉ�̮K��$�WyW$	A�X�2��u6��Y1�~i��(�'n_E���8-�
��y4��2K�#�vSŉYI��h���}�S�S0��¶�Ŵlbh1��6uQ�!V8/���}�EN�@��""$��O�	��M5`�Av/�)�I�n��r�*Cα)��XI�0��'X�8!a3�1)�dxy!���� r�e��s�Ʉ�3�}lR��ʎ����Y^�P����B� <Հ9����[(aލsH���.�y�[�~Uྙ����&�TK2����z��{�Q:�*�(����C��t܊��5�3d���X���#�f�@x�6�!�� Α��m��J�Y�n��vL8l��
D�2�1C���g���2�%�"$r�A.U�&l_QC�*��v3�<>eU�B+�� �^f��y�(�6㶢B��V�gM�5�V)�����>D��JJ�����P RſiK�Cӝ�@�}���I�(��λ���^�@ܷ�lȹX@��d�AQ�>��/ݖ���a��
D*=aUY�Ҁ�G� �E?�H"\�G�����a=�/+
��u,�l��Eijm��}���i#wK�s��]xG����I�q�g9�)5w�YU�R��EP��J�G�̃!�]E|V �*���U������X���A'�qzE�zӚִ�5�5HӚִ�5�/����rs1a�Ç���� �g@u>dX�.3�.�P����어b�� �N��2��T�+. A�\\���~�ʃ����k�< ����\��0���� �F��t'=]P��q� YS���ʂ�aœD���pف����s�� ��8!��$G㩜]\��ٙ; ��Lu�V���ҲԿ�����F��fE`�;��3{:f�l�8��8F��e���� 8�P�2����կ~%�~��U���{
�������������S�vY)zy~���;�BAe�.n^|���B�=Mi�h ?2Os�h_<��1d����@����+���d8��u���^�81Oi� �@���d�Hh=��s}?�6XU e�l Si�hDP�����X7�}�T��	�.-`������N�q� ��z�2�]A�$#����G�"k{&��G�Ȏka��C�V�v'���>:�����y+��M�E�ԭEFpT��H�vS�ںE<ǁ�L��1
	��a��c�[#�Vܧ�C-9���H�#��U#	Ѣ�2��� ��
��=,V�9�[�^���c"W�
�ڷܫXY1擐; ��B$�%����G��;HI@玡Q}�J {�{q�$oѲ��Ø�ݢ��C0��5p��KuO@mC:1![�lD���  ��IDAT���f�VSaaGI�&��{|DQ��j?�5��Ȩ2~�׺���X��
91	����A���(�b?��OaIvQ�3##�g��~�ҭd.G]f��a)�)B�@��OD����zt.�<I�Z(*�p�K�N��.X��ع�^3.�tB�s�D�ۗ��� ��f1�r�ۡ�*��2#�*�È�Zu�$\;6�,���&pU$�|b[N��(�01�-�o��0*'M`+Պ[�a�~�BԖ������̮q��NQ���q���-�����Y�?��$/L	H�Vi��0��`*��Y�������dU���1�*�Z�����8b.��f�(��U�Q� ��")��Tï�����
�6U'�i����F�3v|��!w��?T��uYS�������уG����=0�:2͌/M���5P@q�y>̕��l�~��v����'bn��`�4[��D�y���C;}*Aq?B�6*��q�S$f�z��5Z ��'�+ ���)�siY�H��wP������X�V����rM��WT��S�C�e�$�����LZ%���d�l�@����ZZ�\�T��(��Mm�}���$(h�Z��	959��L�����Y�-���x��b�z��Dv�B�@����s��a�zu}C�)<�a<���d,A��2@*nu�W
�P�s2��<�;v>J#`���8���
�3��$j�zM��ef��bt���:,��\j���~�i��P��v�P:=(OVT�Y��t�KӚִ�5�?Nk��5�iMkڷ��s��Xl�a�������2�;���J�ON�jt��B����������W�������0P;����+]�|N�\�APӲ�D�̈́+��p���:t�,�o#�� c���,dX%�K�~ G����l"ף����S�A��Ϟ�˗/u� �Vrvv*��Z--�C�\q���LtVOZ n����d�
@������wwz���ê@������˧J�� �u�py��g�O��O�?#|&�'��^�Xwi��~�+y���!�)�ǋE1�ϟ?g(Ũ�7-#Ëyf���	h��TP�Q����rQ��0�<��8�@'���.��H�n�	2��y����v��NIZ8X�!X�#X�
 "q�J�]],%�w=��G�����������>�N�P)�h���mj�������������"��8���}/���AG�K`�U�z � 	�Pa�A`uR� {+Z�y�h\��1X__x��ޭ����L���h����)�*#)Pe/�� ԣSY`�ĔuɱoU�^Z�����-���&�jل�S����mM�&�+��]�����m��mٔQ3b)�KXT��� ��TB 9�6��tC�1������@K�����,�͑��+Tp�nSC��el@�S��ion9������v9�C1���ڀ�+��%֝DNy����l�r�����U��|M�,z�@L� ��c����l�,	�L-�H���w�a}:�Nv��p�qȩ<�@��Hbxu�]uFO�y��_��{8=���P��P�>H�3�0�cW�8q��(��#O��,����YDb��@B��0����R�1���G��W�Ʊ�>���γ�<�}�i�m��t㸳�!9�p����j�g��ԤqP�X����qg�w��X� ����b����Ai������ӠNxT���ֶ���UT��
	A�GP����VN���zOه����O�%���S�-�W��M��֦Q���X	��j��Ex�mk���7������6U����c����ה*TTU�ۯ���m 1_�|@x�;�7�zWg�_{S�{G��sB�c�)GN�~ĵ��;$BՃ��s��T#����dX�&|fkY�H�����|�\��R>;D�R��H�2�wp��8���l� �C���d�q�Fj��d��A�?���i���Qe�A�yl%���I,n�6�\���rR*\_ˊ�`P,�%[�V_���/����p����G��ZԟW�c�����ڞ�T���$wS�53h����+J?Ȅ�u�6 �P�}�1%p��y��J��d2��H��P��<��b�m����(JޣH�6��F^�T�� !A�Z�
���\֓�|��;=���=^��}���r_{��C�9�(,��EÝ]��Q�Y^	�:������l9��z�iMkZӚ����iMkZӚ�o��J�^â��}] !��v 2�g�7��$F�����䂪,f���\���t3y��}Y��2�����k]|%\&�u�xrzB��ũw����C9��!0�d�hX�dlՑX��a �A�����b���<���K������?~M�(��X$~��g��'�����+.Q�OK"]�MfS���ڨ"���Ժ��wy��t�"fz\�F Q����O��.rd]�l�����[�����U� �WK%�}����m����}�\<��D���..ots��a�� ��W�X�.s��܃Iu��w������vO=X1P�0�`WLR��˗OYՉvvr&�=�}s_Q�ȵ���Y�_���)*�ynV8��$�9�P���,���2]� A��eq�$b˭��լȮB�1�������#X2��X��������,��X[�[�"���N� Ae1�#���jN 	���?���)���+�!���V'���>��a��A�.�%I�l��bV(�?���`�IJ$�e �S׭���ձ�Y�V�eN��60��j�0 ����_^�M�U�x���@�8�����l���,����w����ͮ�I�1�ztzZ:�l�����#%8OJ�>�zM'�mk���-� ����T�-1r�f���w-�Ŷ�։���7m���?��f�7F�Į܈ו�Ei�<wP#EF�༒H��#hn���ҧ��cм��n�>�֜���h_'�בg\D��i}�	����fq�/�֑8 g��!������,M���N6�%�����A�$Ւ�EnɆ��p���R���Ǣ����$ ��(rEL�c�,��v2uǽ/�J��q8����~�Ub�ped
��X��I���[��Y\�f�r����H�@������`uDX�,����̣�Ԩ��1G+#����\�P
�vQ)����D\)�$�y$�c )�/�B��^o�96��T"�ac�{E�p��n���
1d?2�b��/�܄�P��u0��e����`}Q���Z��f�2
�^��2+�%OiO|�I�'*hA��s8�ٗ���=9<z��3ؑ��gNr�pͤ6eR-{��}���JpM���:K$;T��e�ߤ�J���;�'����3}X��*�����/����0�v�Ưo�ޚ��_�*L��+��[-������zm�ْ����u�s��()+��O���<TڔNoF�A�I��Ɍ��K�6y���";J�]�-_��5�+@���a/Zs>@�c�>�(8`VG�1�κ,����Y֍�q�-s���ۖ?�̎���T����z��d狕���b�PH��"���>x=�8"�s�3)sJ,�c85j��$�y'�\2���*<ϣPO���,�{��-!-�l��f�%���q�����=�v��t��,��_(T�\Ӛִ�5��_k��5�iMk�_�����]�����-�\I�j�~ǁ*	�v���W�FEF�g�j:�������g?��G����S,�F7�c.n�r�ߓ��B5�AG���������\]_�|>�]]L�� ��1�B���vr�B��?���S/����?b%���K �:�d|3b�(ɔ"�J����tq���ý�TT ��bs>e�w�ߦw6 5�R�s_�X��E_������6iK�K	^�b0�Ec�����%��JXlΖSf��r+a��U�P8<���#X)q�	{�eJ ��6�& ��5*,��S�>� }3=.�驇PC���������_��{T��G������vC�L�p2�^�C��J��?��ڧ�g@ 3x�Wْd|��Piy����⥎��������/V+�ޓt�q�Vټ��7�-�Ƶ����C����a_u����<ppP���-j�D�ח}E�����b�??�����W z{ݍ�M�����An�ɨ�$�W���k�E탄Yb�����ն�vj����v���+�G~B$��L�a�����Ӥ�z��I�m��8@h*��1���Ҭ4k#�ŋH�$���#K6$W��m�~ BC`�������^e��m_��#���݀�d�<t¦�^��t?I-���Ҿ��G �p/��[��8��(��w8�`T���W� :��2��M~1��~{ȹ(���=�we����xp�ws ��Rװ�A8�B���2U�XH\�;(oH��նJ˄JQ��d��󶾋*�$����u�q��m�>���>�!k�����M��(9Ol6Ċ�:tKn����<֠�	��_�7�<�ղ��,�;�ܗ��<��/9�!k�9#��T��v�����N���[0�yn;����`a��"w �����,��Z��l,�@.a���\��YQ�L(҂\��Y�9���U�*�ȯ�h�*Mi�9��(qHH��̶��zeYa�a�{�D�	V^1�b'�8V�VV]�Q���߾�K�~�\��;$�m�^_�*x6����d�t����r�a�*�hm��򂈠��goͥTQ�9����+s~0��Ԭ;����@��&�'A�t�s@H,`����TF�!�vl85�U�= |7^jө���ʈ>�h�.*?�p�ýsՍ>��N���g��L�)�9l���J��)(B��5�Hd�-����;��h�I��U�e*�����T~��1�ԅ�(��v��9��ס+�	m�P܂�j=���h��:�%��r��ضݧ1^�z�s}>BnsF��0�}��5��O�<E1����0��c.���+2UJ�br���l�MW���l�ri*��H�삢��=b�]5��huj�����"0f��v�s+��\�/>�����d"�),f+�$۳zӚִ�5�5HӚִ�5�[�@` �m�e���b���W�U���c��B.����:�D�wt ��n�7�����	������	A�A�͠mT�A!��j, Atz-Y������ꍓ��ve0R�q}s.U��������a��V*�#�o��sA�����R����f��G%]�K�l��j��T����^t�IB�~��o�'=+~c��,j!���G@40(�Ȫ���6��J�-��9+�a����+�y�Aڨ
�����
�Ԋ�a��Eki�(��$Ndt;�����rP�L����)�þ����e�	��}Ϊ�<�N }�n�>���3�ǇPV��@>@l�Ű{`p+�Y����`�� �Ll�y'8�}��_*\�v'���F�׊�j�v&�ٿC�C�Yfs�z�n��[�����@sT���(TwZetbi���0�A�B��������h�e������~����>]�����z�@I�z_�J-@U!���z�>�)ۭ}��V@6�BaO�x����ۗ��M�ƿ����A�k"0�M�lWM����[^U���3��&��ۭ�灠�X~@������̢�_�Ca'�v*	�N�
�8��q�����ϫ��V����*�uV�W�@�l�Z���IŬ��䚽s]Ҷ�DC�5�o�F���y$ިG�hM��������E�����j3<7�[d������Mͳu���9;$o�4k�8� vf��gW���8!1 �fvCF��[����z�	�h��,���O�ݒ�z��[*��k���,X�QMQ"�mE�T+��NiiU��C��B:�)G�9b�]7�����&;�/���k�e�� �xf��3#��Y���)Y�M�*���%#kE���A������̱+����;4�����y�ZϷx���mbw�Ձ���U����\zE��<���b��J�"#u��>�̍���b9<%�\>��c*~�w��v�ʠ��]y�	i<�[ʵ^1�4�iMkZ��zZC�4�iMkZӾ�UZU�|���� �A^`Y�D��U�FT���t���f��@emХ��>�i$�_�L��>)7�	�f�������H>��S],���'T���C�Q=���?8~d��l�s�]��s�g�Z���GT,@^?�12�)?��B��؂�1lR�2�/H�A���e�-�	�0�8,��[ ����:�:D�-T_V�B�R�Y߉D2��.ҡ�5���W׾ N��|���|E{�T��n�/���cQi��DX�u,�5�tt���şA(!�T��-�4����'&"��ѧ���#���8T�����Fm<�XY���k���}
�ZZGYr;kQ�ba����ҭD����x���Ip�/Ym^�Ų��U�nM���[������~_�OG�*�; ��m�_ /��N|X8���j���
 ߟ�*r��S��_�}�� ( �Q�v��~%@�5Z���^uL�}]���U-�������*�i�5kb�O��ngm��
򿬧;�֐m��E~�k5d��xM�����F��[6P���{+	���|�޿򏟧�xrb!k8��\���-��V���}�c$�W��G y�����yvsߞ�ͩ1������u�h�Ve�6y�P(Fq
�%kF�a��S�ܦ)�UA�����k�2~���V໶l��w�\��X+P|E�<�����2�~6(<^�����c�����9�+ӌ{��v�����>3�&+��Z�p�nQ=��$r�XnF�?[%�a�e���o/m2�秕.��x��z$E�gD�U�HD_��}l�g*XV[ʕй�f]M��6��(��ǟ�0���x=�ڪ-�'�Z���UTl|��Z���!\w/���J�N=I���
aC����ض��V�s+��2Ri���5Ӈ��pU�6[��q%T�D�T꥾�Yg4ִ�5�iͭ��ִ�5�i��Bfk��ʗ�U�"�KY�|6�'/���J�7���wgg�vQy1�E�������_77_N�5���X�]�:\��ӞA	2�/_pa&��Z����r��\�rE��G���.s�%��o�"6��xƜe� �
3�F�:������A���-����F�^�� �!��Ќ�0og˺ؼ��E�/f��}G���"^̟>r�|	��Y{�}�XL��L�:��+,.b'��s��S��E˕tڦl�������|��o�Ww+%3&]�/���_��@�=�/ �ٰ,J#셥�Т��Z0�ٔ�lg��}���!�����^��q���%Od�Z�=�9IZV�Z��-�J˼���\��k ��|'	���愿��mc^�k�k �n�4���6�`��aր�6>c!ڶ�����O ����?w�Z �������mp�x�y���x�
_���w�&m��Aw4���N�W���U�Ǘ�_k|1�Z�v�emug��L��U��+���wݧw*���w��j-&��喁���w2aRx�o�۝��Mګ?拄��j�U����:��7!�n�Ѿ����qrK��S�Ds�ֿ�d��r+�����u�ʾe�Pn�?�����/�wy'٭��s����a�ի�=_l6��w>7��Qb[Yڶ\�R�ܘ�j-a����Pn�#}���*�bځA`�BdR�?iKz듷U�~���m����m?b�X�#m�P8���)ɍʆ�>ڮ��}&/-T��tZYaö��~	a� V���H�M���jY�>q��1Z�r��HܽԷe]ݺ�G[[�g��V\I�JX{%f�r�B�8)I�J-1�M���3d��Y�%3�%<kÚ�{x �ٕ)e[Y�iMkZӚ��mҴ�5�iM�ֵ�����>$77c�|������/������}y��ߓ���t��/�2_�t>���%��Þ̦+ ���I]�Ky)Ū��$A������<%�0��!���h��奜��K��UTB�U���T�w�I'��)��>)+V�-SY��gRQa�%-�*�,�  ��吺�]�2�Xx/Vf� <TN�Ϝ�\���A �`g�V��E|f�{�K��lh�Г�}��@�%�����DLP`�R�g�~��+�-]K��46i):y�Ge�jmg�q�}Ǫ>xk��$��N�e`���CL+Z��j:1on�m�1}�L��d1��y2 ����'�s����I�s;��@�����<�*���:ߠ���O�ك:Dd��l6�j �PT���ɓ0>�6�;<���7��K3} �oȏ�T"�������n����;���%A�f�uL_�x�K�W*��w*��������-�}�۟��T�L)�o�Q�u���F��HS��k��k��K�斺��6�u�Y&��ϭ����Z_G��g�m���\_�տ�9k����������
vW��T[���?�O��r&d���>��!���=-��)So�9���ZT��$p"/
�7�%�q�ԋ<P�QEz�-@�IP�������)<� ��n��X�,����>�o�(v�e|�� (>h�tw�ϟ|6�g�$9uiK�S�� ��|z��TÆ,��	<á�"��z���d�7�A���2U5Ɇ��&?8��o�ެG�-��6�S�w�;T}�UUw���+O�H �/h��_�@�' ���PK�/A�'>5��o�{3oޜb���>k�s��-��=2"oFfپ>�;fn~�^{��I�g�_�iN��prWmpC<3��iq�<�z��ZO��{u	�4(qMZ�����8��W�>̴1�l�@e��@N)��HUмw9;ӥj}��]}��G�`� H}��G�&j&�����c6�˫W����xn���<;��K�O�L��DNNe0��1�����񉜜��$Y�FJ��������݀U��7�aT^Ƀ�s��#������痯MBZR+��/����>?���5�c:����C�݀]�шc�de��AB	��X�⽯���b�.�4P�x�Kl]7�J��o|�k���ߪ�Yy��Ŕ|
�����!v����Q�d�W6FD�-P�P���ٞ�s��IIh��~�2Y#3w`o@��(~���K&���m}A�4��6Yc���a� ��P����|��>��̫A0�yDbRmk;0�/J-h�Ɣ4[f*ρ����W+�dRf�z75�V����FgK��uն+	x��������z��u����Ƥ��;��w!��ֽ�&�G��f ��u:��+���;���[�����N[�sL���E��َ�|u��^rh{�gT��N}�ڲ�]��m���g��=W�vrC:N���D[�gt�h���}��~[����.3�퉴��VK��Kt�y욳_�/��q~2���~���mc�̘�Y��5�����X���lk��{���D��ZmH�$��̡��p?��������K���o�U�^�y��@�eA�o&�7���X�ߧ��
�n}-��h)a��-��[P��(���a��Z 	~s]꫱;�]f�7���X `r�gv�9���
ҍ��gt �z�E��x�B�D��5�23����{���.�����t);(����?Ѓ,�'*V�ڽ(����[�� �<An1�ryfVw>%��裏>����@�裏>��a��u��gA~���8Eo$�K��ϯ~�l	�O��cy����DL�2�]Zy)_�O��v2Y�s�M�	�H^����H�`��_\��<@�������<W��7��p]^N��g_�� ��锝�y�{��Y.�h�����iq�I�3�D��~Ld�YLf+&��a�_�۟v�Y��Nñ>V���s%9`��j2� �.PH0D4#W��#�bŔ-g�C�`���v!tVJ��`,`� Ա��TY�ƻ0n�\z�����,2�/H�yo0$�K{f_寎��I��\0�\��*U�2�fL�����K0V�dQ,ȂPa����0RZ ���9в���P��k��]����a�2~^/�X�ε��Ic�"j�*�ի�ju�µ�ޑv1�Sl���Y���H[5�k?��s�b'��t��߆���T���H���X7>���Vw.[�r��6�Åg��w�����q�6Sa�5�=敤���H�K���7���g�����,�K�P�x�W��:3�=�. ە)��9���fc��u��5��-�no�ƺ�������-����E�ʤ�6�9�������U�~���A���c�o!�����t�<0<���b���Y7Q�f��b�5 �Q����v@�\�i�����/_�����<#��Q�"��\�o��`�����/�̬1�����1k�Ad�j=�tN+�K*�h`3	��m�_i���mG��mʳ�
��i�6:'"Z<."2Z�Np���tTk�k>��V��).Y)�>�u�����dc��5�`�ʚ溰rM?*�V�S	��b��G}���F���G}�q�X��;�L���@F����b�`��?�x!y6gq<I"y��9�Hg%ñ�  Y���Ix
�����IY���^y�n��$MH���9;?�h1#E�jv����/���$R�?8���/.�2������?J�rz�X��]weQ��O�����8NTf�X��L�(h"�d�H��5���[F�M �8�v��G"��JOT
�����'�C��� �8���۟���J'�B�ʺji�ה�'&�Y^��S3�W�n	bJR�)i�n>�:�?ag�O�s���?�Â�潗g�48��be# �a�OC���	-�Q5!�P@�[�QV�����{o]�SM�bD�<�.�-�>WXۢc�����Q�,��n�n�����(\�ڿ����UDV��yi�Ű�tS��c:7�5`��Ҵ��
=7>>�9]��~O\c[Я���ۂ1��竎׵����x�w�6W]�ۃi�s�}�-�վV���t�huq����p�K���TvN�L1�eư-v�A���Q��q�MZv�n�o�ߒ�����P��f�Y�?��P��k�����[�.VM�aی� �����Y��7|?ெ�LA�4k�zfօ���pmʰM)V,���B;�i�FW���s����C���e٫,�jBVI��  �Z�Z�X�f^�t >?k���1��o)������N�
�pT�����S9&�?<+W��`�@�k��z�8o3�����`%�Z�d
J�V���KF����{6v65�/��t/�B�裏>��|�@�裏>���U03�Y����$�!�2 �?b���穜�M�ȹ�������W&YZ� ��ѓG4�C����L|,�	�KG�����yݿ�Oe8����rv~)P���2_,���726��@N ��/d6_ȷ�%��'��8��r~>3ۘ�p���hL�M����x�Z�P��,M�8@8�!P�/$e 	 � ������?�k�f�1�t���k�o��M�󨽚�yt0a�!��s�4Pf�x aA`Ì�4VO"�Z6� ��$�  ��P�`�( 	�Μ��;-!c���Ш���| �OER+O�=�ah�F�Q�,3�KJe��.33'I!Ǚ�3Ή!e� �̦����J[P^F����I�!AFQ«mq��b��*�U+�T�u���GR7FWTD�m�*]���hq '�IZ����N��Ck�w�QP[k׼0��kz��6�d�m�/~�M�i�������+Qi��n��-�����c�]�W�e���h��}�e@�qw�ˠ1���v#�|sӕ�F{��<R��aǸ}�Uw����d�z'�d(�מ���X6\�@ܰ0P+;���v�k���]1v����~}���ж��sѫ��/Z�=��;׷g�Ok�ς5�t iuR�~(TVk���ϗ;�]- k#Xՙ��k��$�^ל��u����(��sՖ5�7K�����<���^�X���w�މhm�]�k�d���5�oEX������kv7p_��B�Uf����}��g?�U�<����~�� �����<�z��_�I24k�T>�fH~z��س!�,��*ǚ���MFfq`�4��a0/�g�
,�Ri*�	�k��l�p�IZ��c�"���*m�?�Xs᳅5���cT�+`���*gZ7M2e-Rm8w�I��@X���>���[ ��hz֣�+O��缴~o�*{UZiU���@�̳@H)+�uhځ_dQ�<֒X*ɬ� |U*�{�r�l`|&ԏ���2�� �� ����G}���'= �G}��ǽ	H=y^��;�!(��4�.�0���E*�uq6e�&-L6Yg��/����#�yr89��� �y�������I���!=<F�r9���z^���0�0	�O�^���fKy��B~z�Fƃ1��_���g�-K�����\� ��ɘ��@�
Y,��*��K~ ��3>��n����7:
�(���l	kZ�ȋܚ��s����G`<H`�=<�Vb���L�8l
�HH+���f���G2&�#�N ��!�YT�MHq���Pb���h]l���M^�4�tA�����r�r{` A�"���\D�_���� 6�HԥM�/d<�H2���L�0@7	�E��$�c�+CQ*`U�-��U	�nl*�^-%��J��F�zS���IE��� �?�����J��b ]��� պ�Ȃ�-�ō���6�=�Ғ�P�k�d5 �W�ۢ������̾Qu�w�5�fmsm����e�|��W6k+Hb�.X`�v�=��q���&/��5��z@w/b�~��^����� �Fޘ#r�uLs=Ǚ8�t�F������e���;HͿgf�Y���rr��F���k��z���b�U+��*)���.c@����LT�l`'m��L&�߯��e��@8��+�
A?hy�Y�s�c�����b�Y_�A��s�sYHDf]��_��5�K�vl�K�Ĳ�{^��r��Y�����X�裏>��l�@�裏>��W)#$�9t�I���s2���O���; I���?� �l)gg��_��S98<�C���K���$K:_�<U���X�Ifa�t��p�Pb��X���	m��//f�f�K��M������b�.?�
3�2H���1aF.���H�k����xrr�$mz9m���~�P	 L$�.�C�&�  ^�c��0~��H�Z줜�'����_5��dA�� ���VƄ+���)�
,���&a�!Q ��VA�]}����(ZL�kpN�@PK���UAڎ����vĹ��ra����H��ڜ7��^%������<
JEX}h��RY<&���|Ziv4��*N6�_��[=l���M\�ˎ��"��tպN�K��>dl�겅Տ-��d��c�:�w 2,�K2p�(,��X{o��h�kY������.v�]��S]�����&�ݽ�� ���D�&�㯶WY��N��}n���4�mF�M$�v��d!��T��8�򔡷҄���h�ݽ�6<��fY=)�c���k� r�춹ZW�ͫ�W����f���p��@����2���H�}��`�MeF�cl�>��Y&J��~�ڬ�JiHI,�d ��2?��y�=b��4������ޱl�;_�\N2
��C���k(=��S;�����sS_���29����7n}����9�`���w�7�[V�e�X)Nbe1��ȃ׃!F�<&�ج�8 ę�ֺd�A�6���y�Ȭ���_�<�?�����G}���g= �G}��ǽ
׽�߮x?�_��}xx$�����&�s��Lf���g���KY�3����'���I�9:�����D46I�RQ�
��:�;^��A./�%�C�In��b>S��B��ȼ~p��Լgi^�nzn�10R��X�GLF&i���eE&�G󅔾�uY���j�.�ڈRTH� �(�A�$J�����u#��c�2�L���aSp������t�]�n	�QTS�b	���N$fΒD.�8��WU)�wg�p@a���^��W(8�plx��7z3ǁ��b9�2{����ON�����,����e�xSu=f�� V�G23���V��8�5��G��\�J����2+݀�
Em�ܖ���bᕪC-W�
P�ا�t��'�p��m��{8������Wlc�+S��ض���{�r��;d�����-�Ŀ�[���q���;��������.�\d���<v��m��
+��.��Q���0���G>��^K�;?�M����{�C���\y]����mZT*��>V�WmЩ�o��D��W�W�	�=�R� ���zdv`���$_�/��>h�������k�d��՛���}�v~8E%���d���]�=�a4k ��j�#T#����_˚7�$�{�0�Rԗe�\�~�����w����x�!� �֙��˨|E�k�R�"������9��]	g��dߥ��p?Z̲��M��>�裏�2z ��>�裏{GǇ2�d����5e�,�G����i.�˔RW�h ?�Ï�����Dq6�w��x��/������N��K�����ⵄ^"�陜��� �䋧_����r��B�m �.�J^�f�9::��Ne6�˙�~9]�x���L���|r��+�c�d� �)�P�%	t�!uȂĚ&���';��z��
T�u�<"H�8!�0JFq�"m g�f�$���;��e��cE���:U���$�&��	���nC��=�P�/p( ��Ȝ��x �t.�s������b)�ɁL�ǔ���8!�ߎ��Xy|U�&�(�I����¬^����W`~��X��*�cG����$����\�ZH!^�ۋ�P..��d9�_\\ȥ������1�X"��\N��cw���?^���#X֊[��t��w�T�[�ul��x`|�q��.��xH��@= ї���g Ҍ��)�g�y��O����7��l}��s��5Y�6{���F��� �����;^�7�\}�u����ΰ2ZW�S8V�6�~�1�v��֝�Y#���:k�ּa��yG������z��!P�2��$���#hb	̿39�x����ˌG�I���B�Ј���.� �Y���J�/����b�e�n����_%����8��hQ�5`�@�g٧� ��6I�2;��j������)B6K�L���k��z�`MZ��бFc�^)v��DA�p=,�sɋ��u�;��\'�'�uO�q���G}��YF���G}����ɓ'��ū���`���=-ơ�=���8�NN�Q"���N�/gL2QT����$���'C��ٗ����w��2���իW2�'e�b9<> �^ ��!; c������"�O��7o�9����t�שzE�(�9�!�F˭1L�}� �@��Z5���` X�c����$����o� �¨)�R�������3��
Ƃ��p0�\q�>V�rT(�����<Y� e�x��aj�mH6
�{vv&S�ה
�0�,�4JMb�,*s��	v�Ր*(U�;��9��%��d�P��,����Z�O�"3c4�A�4iX(�)��V"�9���!%����N��(��O��/̹ �4ڄ�����BS�D��%E���S��oԿ�R��T ���6	�?�*��jZ���'�^��Y3��u|�c�ԉ}]�Sl���=�����y��w��A��;,�o2����HQm�A���o�`x�pfՐM���{�o�l;M�`�J�]�q_���}���o8w��m�q@����{�װL�3�����|n���?Xk�a���3Fo��Zḧ��������RY.\�\\L��/��l�/�R��(E��\
XH#�~v,�^6,d���#pҞ�)���s�Tiq��Q*��aW�����#�
�ߕ�@v1A�6$�w�ͱ��q���#��;����y���&�Z��	���j�yΔ��ł!�q�UT{^l�>1�H�=2�;�����������J}��G�U� H}��G�. j��RN0���D�U�����u��XFc)+O�It��G2`�>���<X���B�0}��3�*�Rb�!<9�xG��dK��\^�z-˴�,Y&9�S��l.��R��1N�ȟx!N�y���l6�A� ��n���0��ٞG�($�R���Kʜl�X��:�b5/K�a]�%� �d�-=ɪ��C3G��봐=�e �9���>�s�)�U�},%ϗ�}��h%{��cd�[��Y�*�� p��C� ,H�k��">�����`��d~rJ?���j8�kMh�`sp���T:/��9�����9%{�c���(
eh�h82��/�%e.\W!�!aL����I�5ހw`�C��<>>���|n~�W
^����ʫ��U��@� Ȯ�Ӷg�.>���D���*Z���I��W�g�%���}@v�������u��"����wD��>�Q��&�� 5�i]4`I{��U鬶�H�wa��l�KPڒ�Zc������we;������Ǣr���0��̄[I�}ࠉy�^X�8]w�v>�T�7?���ί0{6�o�=�o1�z�S���7�4M���G�kp�����L'd5��-�S����j6�p�=�(�˺�l�k�Z��YL'�߱ؖO*i�l1��K�#:d��#h��f��̬1z�#Mv�+��	��,�D��Ϣ�o��@>�Ypf{T�sP_��o ���;P����w�M0�
鎣���rl^	����>jX���o0�qm�a��W�>�@�h�9��������yf���@��0EG&/8(��7C>���@�裏>���aЧ_>���_�㯞��y6@� ��Xf������Yh��=>�~��|��L޾��墠�6Vn���&�HF!o�Dԏo��x|�d̅�l)GG������0���wv�N~~�rS<����RW�L=?�Q�f��Nd��2W�j�Bz�s�K����p�r2L��i)�~�HU�ʶP����}�KM�3��#�����`��S�ʗ�C����RF�����Waƞ�:JwE�_Ă8(Ԕ�8f7$�d�)P�')y��e�svttl�H	��Yi��2@0E`��1���E�ۮ͚�X`a,�������&���*�1j>]� 96#��@�L������p� /�R돏y|I�9&�a�3�L��L�rzr(ss�Zdu��%�u%�h��
k�=�-���^�b�	��z�D�	��ڪ��^0U�\Ow6$	XT�����7��������u�;���V�P|[���z�|ԫ�(c����u���}��!��|�ޢ�z+i=_ez��
�\�ݕ��kP�+��w{�k�Y�B}��_mi�v܄I�����)ų�� �M̔=��0m���і�r� ~�YIFG3����5�� Q�*�s�RY� X+�1Mfi)�y]A���1�xD��~l>�Դ!dh�(G��\�A�/]F����xl���E{0DD���С_�QJW!5pLx��m��VQ;����/#��Y�!W/ݪ���90�k���D�Z��B�dq�Xx\��g���cU�S����*�a�s��8����#�6CH��� 5��lq`�����?����W�G}����= �G}���GJ��<��	�ЙIb��T�A �,�TҜv�R��dF(�ϖ3�M4�������W����?Sf	 	���Z��8��d���P^����y�� /2��.$�L�����}�L2�0�,$���e\:<4c&C�w�Sk:�2&�H�!��GA҉�>�D��9�g @&J��2�催wF�$��́�9��������f;'�	;ސ�#���2���y��pb�w_���'rj��ӌ�A�X�*�ŤZprf��7�&�C3 )��K�4f2>�x�99>��6d#0, �4s]ntG��9F��R{ڵ	 {�\D`�
���kɭ>6t�1A.< �@��4�1�b)�E�m!S.r�}v}�!�R\B�3�W�k�b4�ȁ��+4�	}h��H�� ,�6�(�E3o����8N��Iam���;X!�v��]m����J�i�@c�]�[��~�Vo�-�o�m�	�n�-��&��~�u>��� ���OW^o�W0n�����VK�x_鿼-��H`���j�ɲ5�����v������r��t^׮QO���Qke%sE���RY5��?<n+a�ՀR��.�Uv�-�E�Mu���5k�D*���U���h�����Cۛ��9�u��&;�NA�c���vz�Ͷ;�}m��]Y�����5�O]�����:���T��]��m��+��&I��1x���u "���1�1������l�#�m,��L�O���ց_�� f���_?_�׆��uE�|�����l��ςX�{��ʾ\̸o8(��97롱Y�-�9��)�g�3�oZd����ڈR�5��`b��C��2�~��ugl�I`�b��u߃�c��:���uH�<��/�r��̬Oz�����(��%�Hd�2C N�u.E�m���e`��Y�r'�/s�)��S��.�]��s�9�(�c�����s� �|��H��
$��~m�(���SU��� �{~@��j�M)��M/���`[�;�R|��54��X�
��WL��<Ϭ�=i�/X��Ϯ&�91���9��o߽��b*�ln֖��ab>�)pg������f��7�>�裏>>���>�裏>�M�[�&b=)2 (B�)*-�1߫��W��2i<=�0���W�'"����0?��CM}T�m0��(���7�d:_���9;��T�"�l&�z�����|Ai��n��ԟ��,;}54G���M�!�G ~��1��9��!r�,R��,��O8.gެ�6B	�\^��( S��e��`��a��<ɹ�~v�ߎ��$ynp<�#�uW"�.�y�����<��7�Z�¢b5'�.�(3�1�yl�,�yF��0�am��Ѳ�D^�?�<�W	�$��R2Qf��UP����1@���jk��&yΥ0s�G��

��;�?���\/��K���_Zk��і�n{��)����O�6��������5ZB��ގ��-,#g����r�k�
(�������6���������^�M�i÷Fe�:����7��
&)�A �G�φ	��p�ٵ4��)��Ԣ\*ȜF����������Cz��}\[Mg��u�RX�� 1�u�J!�?H�z%�������'h�!��Z���8T�.@D*k�q�(�7��_K0�W@��U���~#n�)�(���\����P{"9��k2O��J��E���O�H���.���ec=`�PZ���+�l-�x��X3.�f����_߬+Y�2�XJ׵WVA飏>���@�裏>���<:��ˀ�(1��"OU2��)Y�b���ЂD���$.�In�y��D��'���;n�"�л8_���2�����@e�,lM�/������7���^�l^�J��B�bA��,-L� ��ײ����CC[��F�+�2QȤ-g�ZZK�Zεyݒ���$` ( �|�L
t�����A�Jr��(䌿Uڡn�^<�F��t��o�� (�׺�sBY�X�f|lHX���TZ�c�ٍW����sR #�h�}�$��.�(Ip��E�J�tA���h� 9 �0Khz/S.�̑d��&��u@ 
@
�E�����,m�g���U��Iv`Ԕ�#ˋUe�_u �$��Bm�6{��FW��=����_\q�[�"�Ӎ]��)b��E{������]��s�M�
�^�a�Ǉ���Fe%�Q�Ű�vN���>w����_�}�� �]���w}\|�{�v�n���>��c6���.�@����<�*];	�	��	*5Ȯ*�'���oŹ���2�������/�|��fn����?�`ޟ��O�b�Y/Y!ٺ�eF�f�6�y!��0H���6��5�.�Y����)ǆ�S�t�@'��a�`ԑHh�ؼu���h��U�kr�G��zw�+	3_�]d�Vn>A��)UZ�w����#G�a�ͬ��ذ.�#֫�sf�>Lh܉�vu> �����r�$`��sA�����������>�裏O(z ��>�裏�,>���A|99y�F��]6�*�P2�����p(�������82�[.�����gI�G�D�˄� O�>��耯===���sɗ���R`��s�OgA��8��5�U6
�p���e�)��EtBΠ��\��W�C�~����8$�`v xY����Y!����jf�Q��Lf����0	����隆��v�q@��$8�)�" P (�9H���Q���]�1��B���<��,2�6��4�W�
t�3_踃�h��J�D��q(U�	�r�ݔ�9�sxL�''��5���B������0%l�(;H��eR���1�f�ys]p2��ڂM��{g�[��2��=��R��ױgߖ�ju�o���1�㵻��T6e�����
۷�Þ�to����Ħ{����${K�ʤ9�c�6�L���X��somI*��p~���}�Ʋ�ל#z�p�+�~��|_��j*_��G�6tx\cD^h�f9�� /��#���y6��DH�C�X�.�0S9`Nb֟֏£�&֍����'��fl��Wm�K����p,�F˂rz�Q�A�ìm������E�d���B?y�h�*@ؾ�zV�ʝ��� �_*۷22�Xb�Q�-���ϸ�q2J5uw�,��V��z| ������@H����e�0֐���y�؟o	h�!3|2�~��/����������}��G}|�� }��G}܋�;�3�%,�CH��M��<���	��S�8đ�9���$3(%N qd�����g�\p���=K�G����7���&������B~z�B^�|!LRE(��	*����r���{:T�["�X�d�K��ҷ���$�%�>�\�b-�[�'�!Vr0A���0�c��y�i'�R�)�7�	V�) �O^��>�OrrȂ=���e�D3�`��!_�ug��"+4��P�$� ?�~)H��b�y!;�<hk�c����P�9�	-$�0g_�Lls���"���	hx� �����)M�a�N�� "Ã�VR��2H��1%�@g����gf����(�@�z�+v^�ZĻ]�*$���}��>6��ȇ)����7��
�7Av� �,<��S��k�:�1�6u�o�����F� w��$��i؝ �����}�S�?�h�9��'E%{TdL	L��\�������`c�$���D�:�c���� x�i9
mb!|	+��x��(�~��[pM��,��ٖS�jM�ʲK,$B�U��-ӌ�G�k�l� ����@C��ڄCyNxi�}6s�=���ٱ��:��{]�+�K��k�^"�3�`��� s��A��v����S�������a�k v�` �b	s�����-xT�9�� K[�/;<x�ͲM.u����7�w�}~����A���I}��G�]� H}��G=��R�	RF�v�9�`A��[~��Q��ĉ��7�B�<ew^2�$����t����9�]��3y��-�C������[��6	Z)#0��CJ��t~��Dh��v��'Gf{&�*e:�r_,��3�P6B���D*����.��0p�86$�3�-ϲ2<o��q,K���Yј��MY1ʔhV������m���G�I�)=z�f�q���r�x>��]�|��H|k&N�N�E:N�*��I'���ͬ�� ��%+U�f��1�l< `�d�x���y�V�
 ��i)�an��{���^m ��^@�x����8�(
����i��+�ϳ�`�/��2�����V��|Ӣ�6���v ��e;ܵ|S�	q�ؽ#��A���d�2�o�e�i�v��>�7n�P��?l��\�k����Q�:�o�Tu�c�\߄]������l����}ӽko���9r&�p�(�_k�6Z�!¼?��z�Y�К��@J4������Ěx+q­[��7�. Y~tAd��c��тr�f�A)�LR~�,J����B�f�ǰ�CU��am&�y�sa��Jsb�F�K ��X~de��� `�hB<o�X�����X
��㺯����ؾ��.�C�пk��\s�}�2X�q�1G�8Ն�k����nך=�(��P���4�;0�ko�s�5<֧f���5nc�Cs�>�����_����������>�裏�&z ��>�裏{�INQ_�#P|�W���DI�J+�Q)CY���W+5�(��q%��Ts�d6���K���r|r">1�3�2�N/)y�D�7I�8I��K�GM�t�T)��l�׿��|���r~~aƚ�Ż���;)�%���5��� (�{���|1�4[I@����z�D�'@I���Ҍ)���5I�߉�[��*��x^��$By��O%X�,�b��d$ʦ#�h�_BY1$�>|�*԰�'@��a����;tRR"��Yn�PL����02�f��1�E��.(�J}��0��e�V~� ��C	X0�7I��L�e���X `�`x���%�
�͢W!�XC���ﾕ��D�ڰ�!��SP��*���p�{�Gb�s�n��& ȾT[����h�oC��u��p��	��(����_:��J_n��������x]Ɏ�-�H����S�]�]і��t��P[rx8x�$�?\%�FRx��*�	����l!�l<�V�[��@�JT��#��H^�b`�:^u
X�&���D��\V��� ���E�m8D����k
6g�-�k+HB��"1�Z�7�Y� �P_5���4p��EVe�:0��б�û�q�d�wo��ì�+4���|Z����:��f�Tj��Ih���h�k�� 4�2W�WKƺ4�B���4kƌkB4�Я��F��@ER������v-�a48!=����X��<2�=3c|m�t�o���9�����K}��G�E� H}��G?��"4b!��y'�3\B���[� 0>JK}G�I	_��YA�*�l���/��˟�ʗ_,TG�$��˹��]�'��R֪,}~y.�&a��� �k0$6��ӧ��+����Ͷ��w�d�X*��_aR����5҆1:� �x����;$K&�HpK���� ��bN�G^��q7'�<Sj�	0��Ghq�}i�&��@ �>�)���LQh��%�*��$�� �`�y�MC �(�e���2u���06�
2Fp�)���X���Up}�0-'hZ�M�5hiǱ9$��I���a�P� �� ~�C ���Ij�*k��1?V����vVn �v3�S���	�n�bb�>�Ý�����ی����~�Y+{^���h��x�������g�=�m�M�dWlB��-�\߮}�3|���}��'��_��[f�6_d���'��8-������B
��$�Ve�X,>(�YW\,�
mlq�� jm4�����l�x�rY��;����O,j����
Ԑ��+�Q� \r�T橰l`}/}A*�����TUհM�	��ʿ��{�Q����k]G5��ږ�� ��}��}���&�J=�-����(!�6��F ]�����LP*�%5� @U4a�f�T��DI43�V���������L�h1�=&������ٴ��_���������飏>��㓏 飏>�����~mR#�<_2�����!:��2�� �=0	�p�ȲX�����T��Zd6���K���S�ĳ�?����Q��ɑ����z��\f��#9=}@��(H<0��b!Y�2��� ���X��巿�N~������I�
��x %��$�Ui;
�1�:��Щ����DFá&�y@y�ԌRH�f�I��0���#��a�7�����a�P�`�^6r_�I���p�`$�b>_�S���'�������� ��n�J.�L��jb������S�#����l1��R��� 4��T�&��*��/1N���1I�m�9��!�����Q.��=#�^v����b&k���,lC}@r�	)j����-sq`�������$���^�]]���"�&��F��Wɢ��R	�ME�
���iv��I52*NӃ���+��%F����������5Z�"��zo���ת^/
m7>��ZǠǶy�6�wM��cZ�Y� �B�<�j��Dܼ�B�rk\�$���1�w��ER�\� �m�w�2����r�1b�US0[/̮G�Zo�{�ͯmϭz��n��qQ����H}�s�������$1t�p���n���hغ6�Ъ�F�w��g�}�b@k�ԥ��V0ým��Up�{�V+@��X#��A�k�y�����U��M��߿���>;��߶�m,�}���>����X6��	X/%�/����Y#�w|�6ܮ�3���`㈓=��b6��4뵃�̺��,X�����E��~�kYdK�z�0k���/>�	y-ng��ĉ��i>�h�����W4��dY�T�6qwLA^�\����1�a��$�ߥ�O�f�j�~�6��{I�������H|��@��2"���3U6��"����ԱY���Ȍ.�f�<Of�8�g�a��f� `�� �qb}��K0�Xߣ�&�w�����Ro1~-c�|���b��h>E�o�m>�#`��@��KY̧f�1�ӧ�����C4���cs{���z����x�~YM�^{ ��>���3� 飏>���ޅI��d�ԑJX���$��<&��z��Q ~(�ғ��W&�{ɤ��kjz/_�c���?rxt������û��L��&),�i��x$'�����_�_>2�W-�ť�f�L�aV	��I����J߹�]|�7�?�-M�����96t���.���@���s#�3���8*5��HɩL�������̲3�ƣ�$K��[	���4�n�I(���	>}=�X�>�h��2W������R��
{�+�Pcn
Hx�7Hwez�0�Ln3-(��2���8���k�^F���0>|?����_���SO��+�T֮EW gǩ�����A�@���4i�G��kF�7)�n�oZ���=Y�5sx���c'��t��D�[ Ɏ���*�f3�����o=ו����� ���w��ʿ�ئ��L�����X�'���޷;?���}�RqW�r/v�-��W������r{��Q��sX��/(�	���k���|����A ��d�ʄ�����ŏ�!��	�� #re�PF�`A��`-���VS!HC_mb}�A�4߭=���N&��Q��[̱�Vm�@<˖@�MYq���,����` ��wX'��"�,�Z4��ei �*�6���sB��>�[C0��6
|�p�qL�M)`o'1�8���ʔP�u�e%vmg��zXw��&�ʈ,K�0?/Xۂu'$�jm���S���-_>�B��yGi��� 3Þ���6����W����������G}��IG���G}�q�"`�.�� >�E���$|�x����ڃ��
tjL9�dR�`0�V<عW�00��g���`9�����C99~`��$KKf�����tf��c��������'��G��٩N�2�^�@���WԈ���T�L'"��\n$�&A��ϡ��&��9$�����Őr�!�U�v�$�@�$�O&Y~�Z�0C����8A����V�$�V�4���%���&�Xy-������TN	+ !�]�PP��ݧ|�]6F��'�MqBV^'����6��-�s��J7��R���fl�+����{R��`,5d�3�JE��0>����=�P�X��E��?�3��5�Vj�	-p��G�[�v�&����k�
�^�p���ĭ=,v<g~"-�5��]��e�}�����xϢ=�i%k��{���m��>�m��5>w�ɵ�0�O5���Ů�n�[;M�۝��ƶ.�n�>c�����+�[�"��=�n��M`�u������,�	V�jL�|'..g36rp-!b:"Q�	�>C����hd���.���0��s��Ԓ>�"%�X��*i�d�Z�Q���f_҄op�.yl���4��8\���P f��G�u��x��\_��7^23<������zXk�V*+����[1x�e*������=h���@R)�A^Q#�e�ʪ�
���p�x/l? �D��W��g��~�j�J��<��,�����U�� �� �ᩲ�a`��c���F �pn&���S��˧rl֔��:�`<�Q�c}h��#s��3<�>�裏>>���>�裏>�e��a�)���B�J�}��p������vɅ�`.d��z��@�yQ��۩I�t�ڹ�~&����hD&Q:����w(��7_?��$4c+��;����7o�V��t8Hdd���s�%�����jv��9Ov���~4QD� ��P ��A��hd�����ozo� �b�&��[���W���;��35�M∱����ɵ݌�7�k3J������i;rj�9�Έ��5a�\P0����%��F�"@諦t��� �˓�'<_Ht'��_����Lg3�O����D�7��������Ur��δAb0��r��~{n���������+�>�G�{�kƮ��>�G�z0`_��+1Ӏ �}��V�[��~�&gպ�֘��o�Q*��o)����Ao���Jt�϶��s�67}��?Q+��IU{���D�>��>th�z%��B�A��yq�]�`��5��!��`�� �30Gܳl	<����W�kh}մ�^�h�H�¥��
X�@�r9';k�/,��O29�%o��>�5�����T/6���̺Ĭ1}�~c+?�+��߅mQ�:6yX�B��|��7���`c�w�Ae�W���^+���{�"����	�J�~�^a�MeM�s�b�E&Jaט��2Y�gM�V X�vG�<�kz� ��* Of4֡h�QD$6�I���R�)������ӓcy����e�^F�	���|꒪�F��j��꣏>��㓏�f�G}���G�83	[�i ��ꚲ������U���$�E��d%�8Ij�&��zO �QCq���$Ue&��I��J��v�A���Ņ��3�$��x���h,��rx8����BC�	G4�R�e�޽;�����.T;��}����Tz&ܾ-H��H�{Skr���&�(.B�p��'��_$� J`�NfH����eZ}���x�P�f��0�f~�$ `�A����`v��A"�̔���,�LgRY_)�i"���e�Hi1t�eu��(
Hf��k��4�v8gQl�e�]����s�A�,�h�9=>��~�K!?�x"o߾����=H*^�3Q.��i��]�95�=J��)
( "��
۟���"_}��� �-�xk�m��!w��汻,̶�QĻsɩ}���'�c���������r���x��i�'>���~� ���u�/{y�|�����k=�v����XA.t����5�/�*��C�,�a<���F�1(��~@�7�?x�r*�N��h��]X�R�X�䖽�+<X֬�R\R�V�5*U�շ*XMoFiA�`e�yX[e\��08"z�`,��BƔR\f�`Ȱ��P���{ʢ�z�!`�f�̲�u�X�!�������� �J�7�@C ��&$eXX),\Vv ����뱴�ᅅYo'\[�߭(}6y�lgO�f4?��3=�(��)����<?�f.̸"�ށ[���f�?͹ rrx$_<zH_���#���3�ݱ_Uk�h��K'0��EY~�7�>�裏����>�裏>�E����E:�w@�@��HLT�X}%��R.�L�`���oA	+���ə�E�yw�0	q�������'L�3tAN�@�e4H���H�V�yZ0�B"v܅R��u��]h�pC��Ę����Ι�a[ 6`ƉC���,���,UJ�r�r�	���=�T�֯��M�_�e�@c�Ü�`T֘��b�ն���H�;T��8�Ū��K)�8��KEp��qI�B	-Mk;�a*=WV������>�q(������B�~�T��D������n����w���?�z��@4�C�uk��7���E��NPZ�s�@H�[BqM�?4Cb�����;F�׽����E�$�}��<3nk��o_`�w��ږ�iwZo2�v��ɱ������
�r���7��˷�o<�-��b�g¾�m�ο��z�ۯz��^D���K׋�S�� �k�x6~)O��������6i�]�����ɹ^�#�.$0�k��|������p86���M+K/�|)"�a��9�Sؠ��S�:&+)�E��*P��D��QA b�ߣ��&֝�#�j�^�?���Qz.�Q�qgf}���l9��<�(��o<��>Y XO�o���8�T|%�E�EQؿ�ƿ~n)��]�XEъE\���4�tn�=t��4�({9�>�"DA���k�8�L�Ѵ��`,�b���VU��>�|��u5ن���#⨤�lv)Ӌ���˯�����ݚ�򠑉����3ט�g����G}��D���G}�qo����Z��& ���+�p��X��u��� ~�0����ӅM�JH>a��#
�"�4�ۧ�r%�y	1�2�W�ޘ�L� 	c_N����1;ɤv�N>+1��ɬ(��V~!����X��e
�H��&�(�#�$�3aGg^�� �$�g	$\�>��
%��%Ũ�\��E��=d�j��^㽱\�j�n�I�Y1
�x�o�f�0�T���"��z};n���	ti]jjY���f�ɀ�- A\��y�9f��bc�̗s3�y���2_�(>!p�@�^�h��3l�[Kty�Z��f��|��+x�� ${�C�ec�!�=����Ɨ��@�;�?�����-L�}$��n�Ym���������S��\��\&�qȼ8=|��} L�Mw��o00�&�B��^˪�C�>n~�ܻs�ib w��Q����}X*X3p��5P�L�� 
�R�+؃A1�"Ϋ���Z�k�|a��3ޟ���>=��Ц�/b�?�Tby`T`�z`Ԫ<��VF��؆]����I �����בz���R9��ш�B4=� �V^�Ռ����k����t�j�,�6=ެ	<�Mm�Kd�|X�5�͂,x�^�����Laל��>�(ba�>@�
���,���ɱ��~nQ��o'�;���"�J��y�{��0�F��Ωk�:88�5��X�哧��᩼~�Z޽{'��0�?��li�{i�4�"�w���裏>��4�@�裏>��葙��p����4��5 $�H��P}"�&C5��j-T�X M�8��y
mf�h�< Qxj �D�~`��>�H�]k�g��`���+Y,ϙHA���CI~�[�d�LtӴ0I!<9����I�%aR�Ķ��w ;�_���	�G�NI�YW�$���t���IMBX奂&��߃̗�[�9��	:��D���� V@��Q���f�c�~р�ˬ��D �����d�u�1�\�QO��2Z��``Z*+���06�k"����&걕��.ΐ&�AlNb%Ǉ'29:0�4��&�N�Q���<��WE��soY5�� d(�eᒺ^ �V��;�ւ&�
Ή|��v�k���;����~�6��}���s�}nÞe�J��*:�ĕ��KŢގ�d��>�k$vhN��1�g?箘H���ߋ�|>���]I}D�wm���>a�+��߸CY�&�B�t��������>q��w�aב#�����%!ǂ:Ǡ2L��0�=$��������
V`�u_�'\'�d��Y��o狥�jm"QB�����aֆ����9/��JY8ǺUIԘܵ�����H6F��+:���U����M3벰�:���b�c�������G��Ե0�W�V����h�S��V7R�Y6�
���B�h�a��C���8&�)m��i5?�dm_"j2�Q	��2J2�wj�ʖ���
���<?7��H��p��'�#�|�'w���3�D�9�(Ѧ�t^�s�0��/��Gc9:>R)�(��hH�+����X���[�����\�g�o���ȏ?�h�ܬg�Z��H���^��H}��G�G� H}��G�" J�����Z�C�Z�!t�e&k?`HaفI� i���0	�I�J�K��\&�d�)�&YH.e:���!͗,棋���\��L���<�//MrV.�| �Θ\"�C�`
�~]��nBޞ���hH\U&i��p̡I��Ut��EZҗ�2	_?]���Q{����-=[R�����#U^�� �M��ͼ,A�2^9��>��Ő`�]*CE�$ɐ�Bk���$��D�_Y� �������W-�al�U+��(J90�+�'�B���LW:7�4�$���l���:�S%�"=�ؖ�@�XF�@�A�� �HLF����p����>���/a�D̛�v���du����xĮIʥ٘9W����z���ٷ_��T&�F�Q"q�A:.L[X����'ŷ��o�u�(p;I�va�1f�Y���X��r]A|Ә}�Z�l��x�� r���sk2,��VW����M��u�i��_9&k�퐁���c�W�Yk&� UJ�*��Ԙ��,w_��׼L��1�����z��-2h���+6Yw�nl���x�*+�T5�L���~�1��<o�����^c���͆i�um�([f�иWĵ[�1��������L�;�������t��fm0��*���Y\�"+Tj3��ֱ�;���������t��{�ςq�v�X�Q��V�`w�������7���{�&���>�g�1�npk3��绨��j��w�&>�4$�^?	�kr������{Í���� k�lޞU�eІ�X.eV�E�x(Qs�Xc���P�j�3Ț�zf�k�B�`X�Y1�:��k��/0@�f��H
`B��#�RK���2�)�5LFx�؞>%W�}� 8�&�R���Ū<�`0�a��'�����ׂ��xx �ш�X|���2ȃ�c"E��iQ6+'�16�c��>~��-ץG��r|r*�a��H@�/x��u}��X�3y��g�_̵��l�Ds�b.��'\C�����ج9��׵�Y7^^^r�+��xl61ks�ț5��4�fx�-͵r0q�V��_�{k֠ʢ������/������t*f��E2�'c��]\\�����M�N��e&���-_=�^�O��șY��̺����|��P�Gl�RV�ޣ .��G}��yD���G}����ž2L�kM>U�X=$��Gw�dh��ArS����S�MS�8;��$f���%����`G@�"3�� 
 $�#�2f�ar5�����5��F�������#	�o�ő�1�P�$�g�o%��f[��\i�O&�O��<��qF�st�Af*S�0&XP����
"0Ts�s�-�&i�~rdT�6Hޠ�tO�VԌF�&O�X]������ 5����"_�)R�P�1s��d�@gK=Y����ds��-6aщ0�(�|;y�D�T-�$�؎����I�E�Fʒ�-�ͪ��q�.�r����<�u��ŠN�˧O��gNpn1�jG�3�q:�fal�^�l��sy��9G������D)-��R�}�N{���w-���!����.�(�go|�xWX6ۙ��m�Cө�e�����uѝ����Z�(	u��Q-�;fWk����<}`�&��~?��q������nhu�߫��~�����厳}���j���A
˶�7�]����TY�f0i�c��k~}�sݖʂ�j��<��*TړMF nB��6��<GM��P��9j��o��m���~�5��,���t�����(��'��*�u[rZ5�̷��(���<~����A2���y��+y���xf}���c���3�9#�*���;	l�"-t�j֢��6뜽� kD��ɀ}������^T/��O/$5kkό��hB��d4���H~|��if�r��6��|>����<4�{��HFCQ9,έ2J�ˌc�g10k�Ԭa`n&֜���c�?������_��/l�ȕ�{���RZ`� t������o(c�k֓�#���ddƋ������u�0��m�glW����ry~P��y}��G�I� H}��G=�1O�:�H��x@�� �U�J#,M���.�v�͗���r~~�DI$�j��d
�P*,�[�&�`��C�i9�Ț@ D����<cB]g�MeL\K9;�2�z��zj 9����9:�2���xK�W^0�C�d��P��|	+��v�h⍤��E�\#vfsd0'`h�/K	�B�c���L���$�����ԅ6��"'H�.ld�Ѕ��.0���3����p�!:��_3y���	�՘��b�%�ŏAr�.D�!&	b�\ޱF�l����4? OF����W_���O&�^�D��Grd��7oefl�:��@��p8�FI;���o��?��sR �Є^�I��
�h`>q�D8!��������	t��`�y��\�m	�C��+I�,��g�ݢ�&ɩ��7uE�o�M|�L��5���Fև�������ۊ����.�����fI����w3o>D\'/v��w��{.��.�g�F[��9���f�uk��=����Ɗ�\<J7��j�.k�t羢"S-f�� �2TU� �B
4���($� �
٤t��+#�6���Ei��D� h�m�`?�f��ۅI2T9V�����Y�R����s�5����M�k�R��ڤ�G��o����o��o��BNN��~���_��Y;Z�Et]�1� �Ǚ���u����\\�U�H9k�Ib��cB����S�dʴ������"9}����L��t6�/^�b����.�2�θ�<pX�ӕ��+�����\�E�t����#��H..�囯�6������7��G�T��~�������s>_ ye��قMNO?�gϾ�SsL�A22��CJ��f]�א�C_���i�5So���z�V}��G}�_� H}��G�(�|�/D�I�	�1�r9g�?�1���5;� ��'�9?ɛ��ڕ���$>���#���%99>U����7�'��2�D�L�rY�ZZ7K�;�y��)Gtٝ�Me��4ۍ%��B�D,���m1����ÇM��d�5�������H0�du�2@�`{�dkLg|-@tޥ&��8�����\J�9�_P@��ƏD����#��o����珤sZ�L�? �f����1�>c2< S��_<=�Ǐ��gGѓ�:�G�9��g�իW�?�A�|qa�R&��$�!��3N�f>���w�db������s3'a`� ����ƾ����l�J��t�z9�<�
�^f�!��NA 3iJ�U�������/��bkԼ`��L���-���z�q����c��=�M�S7G�H�}��N�i��ݸ��ʎ"s��B�۟�m܆Q�.ro+��%�6Vžl��_wJ�u��b�@�҇�d\7���\����s�wq�]۾�2R�k��~Ck`��־JrU�6���K���XܬO�aH�?ΏX܇,*^*�w�6�����*�y����ʠP�>#��}����l�}�#b�͜��k �:�\�5aM�99<�/�x*�oߑ�1��w�|#�~��=���%��������D3��䏇�`6�Iu93���Z�ˑY��~29��������1MW�T-C�n{����#��u�я����gra������q@��YZ�5�M4�)��8���65�OHw�AD&s����\W��8�_@��4s�u�ج1GXC����V�l���&�	ׂx,6���h�5oI�w��D� �Ǻ۬	��F,s����TE��X�裏>����@�裏>�����+%��)�L.�F���  �2����/�k�����s�ta���MR��x0b�Ч>��������.L���d
�<�t�e�� a0&`�@��߼;�^#�#��>���OR,s�$�U!qIP��Q�� �����Ƈ&�E��Wj2�JtAo��B�?.�z���p Cs�W�K���6�Nշ��C���%�&8I{�F�L�c��&�L���V�t7���T��/5�M⚕,`{������`�1/�Ԯ���?��_���{vE"Q�� ��`��Bc�Ϗ�������ß�1�9�9{ O�<����?"�ݷ�$�����;���sWB���y����`���?�Y�g���BP����îU[��< 鴃ɐ����_@[��.-�xMAƫ�D�=�	���E>g>]�b�.	�]�뵛dU�+����@ܶP�����2x�G�{Ӥ�i�0�nb��q�{\?�-��R����+�: ��E�(�->��g��t�v3X��^I���Ҷ�ذ)���6<���Q����C���R~����j+EU���Xg�l�M�s�ܞ���<�ViЪn5�x����y9̽�/x|`2F,���-K���߱��M�dɑ�9��X��boO�-�����O�+X�NN06h�tWK��陪���I�����ϭ''+�x<N♩�j��D!�?����zm� 0b��X��1AbԶ��g��?(�S�3��3��t}��cM6se>gخ�?\�_Sü;p,يc�Z���\x���C����mt��p��.Gfj��3����c�����|�i}�kSۇ�ٜ@��O���K.^�Y�_躯�/��d.���D��y�s�����q�4�C����s�W��ܟ��F�k3]����e��>�K��RZ64s�����X��;O�9cY�Y�Lɏu��Ne~t��mu=��d2���2�|Yr��N2�^bmHs���ȼn�ޔ�!�b�!>� �!�b�!>y@�
V�� ����kK"{�ɤ�k�w���z��dn]\Hj�Ǎ��l
y�����_���m^2�������cM��4�B2��Ņ&y�L������+���e,k�7��I$�C�ŏ?R:	z�0}�ͷL4�]B��Ry���fK��믿���O)gg��[��3� �4�x.�o��o���\^�x)�6��#�N���@~��9W'���(�TH�`6�v3�f�hB�
*�n{��. 	`�-2_���/����&��� /H�q$L�!�yH	f4�D�����%��љ���ל0* T��1J���M�2�#������������Ϸ��e>;������?�O�3�u�����g�?�����I�x�Ƌ/���r�s��ykr
7R���XDe�q4u$O����''�,W:G5eɸ��nEǦ�
����M�����;�I]ꄿ�d�����.�s������?��ѩ�2xh�}�z:t�|��w�������)R���0��,���~��9|�{�i��}<@n��%� ;�= �2� ���ǵ]��
o�Ki�[���/��E�"�]q;�4�>�=�k�m�5'���m?�5�_��<��ӫ��r���&���H߃u+�DS���ܼ>(�*X�Ñ��L�ݽ�n�ؖ��\�*��K}��	�"`�B>�<L:�4�3���N�<�ͫ���T�u�p�t��.];c����dk�ؤ�$��	e��K�^^��t�룭�����6�ۇT:U����vվ� >�s��Y�>�Z`^cMiV�`/CV�Z����!Ǝ񆡱~�Tיc�"c���fsK�9K�A�����14MF��K�b��C1��� �!�b�!>y�4Y�:�����}G�B`����Մ�x0D�2K:'���Ov�e�0^\��xAK�!�<#CB\G MÓ�����f�f���2�L-�f��_/b��c�z�!����_<}�:R���ׯ�0/�K�;c������_�����̏O���sj ܀i8��x6eR�����Q��� ����
 �d:"��l����zs��)��N�_>��|*�qJVL�������9I6A�9=;���?��!l���e�Ǖ,�������8ދ7f*_���:�t�Ԓ��?{����Y�tD��X��VH2˳�O�ﾓG�N����S?z�$=M�}����S} �mr=�Hh�ꀿ�V{x{\__SR��읍��&���m���m����R�L����V�Lx)�V�u�Wu�Q|�Eڏ]Ċ\g��d?$����R��x�v��{�����_:8�O8ľ�L������ݝ��8��Թٍ��g}j���3�>����_?�ݱ����#?�����@~�������;�uysKz�T;&����}�����-�1��*�ۿ}!����D- ���ǽl�-�_�5gDfo�kŲ*T�a�+���S�?�D�ht����+k�Om`E$�'�*G�0(z���d6�����兮�W\�4:�<ې�Ы�X6���������L ��}��P�Sߏ5����r|��/���ҫ/_� ˍy���}��*���!r,�~�Ӊ��t]�몭�%/6:�-A���<��W�w�G��S��@F�=�Ƙ��k��x���3�Mbzفu���� S�)0�)3F&sh~�<��\]�d���,�y�ҵ���:�
c��A#g\�Uz.6�C�����s+b�!�� �!�b�!>y ��a��� ��B��~K��@��ؿ���lz�	���]B�����U^�|���6���J�B?:�㱬Wk��'x�&M�rq~.o��@��I�|6��щ,W��\����K� ��ђ�>�e�z|��7�{9��0E�c�������O�����Y��f7���Й7c_F�� �=yJ*>�}��a:�N5}������5��d�^I�����tʳg��{��LF��qu���/��ۗrP0��\�/�d��.���z=c'b�Od�d���h��6� ńu��$�	 8:vHa�e��1�F��"����@2��D���R5M9=:��lS�|�q=HN��C�^%�v)k&�УN��^2`��)t���@a)�y\��d��ٸ|�F��|h����a[h�a>�o�ǈ�i�K�|��9�Ů}���^w�� &Tz��%�'��P��a�I���K�����>��c}�C���;�������y���Od��S�m��s�����:x�vϓ��+>��7��� q�{?����w�]�?0,oeVy���������F����X�Z?e�=F�hbah��^-;�3,r���f|�c��̃
��<"B��i(l>����IY�Ip��F�z�3B"V��v6Ԍ2F�-+1,��5cR�}��Zɤ��^_ɏ/~��N�&�Lf\��Tk�k޷���[����8~���Sk�]K2�1dk��n`�� ���gŖ�֥�YJ`�� ��P&�\��K\�_��#�(��^��<(R8Ct�7����s��XS��O��S]�MMj�4�1�E2H�b��k���k}8��d�E_DiX�.�1��>� 1�NNkm�\��mp b�!��m� �1�C���|u.GM�g.h�b6�
�&�۲0������M&Gi��6��{{q-ϟ�������+Yos��g�rM'�1�d��fR�g�y�J�0A>9>��l*��\���'�^t�Ց�K.�u%gO����k���y$���H�Q��~|��Ņ~^�?�XE�Q�����9js��O�����.��o$��b��/�ʱ>f�d2Մ�Of��t^�r�������c@b��`V��i@ �����r_�?Y�����$�1�}���\\�����x���	�!�x����^,�	��a��㗀���O?��q���,
(��كb:�Oɗ�|��4�q���H}ghA_^^rN� ⾠H�$�Rh#��<������U���ެ��Av��X�d�T˥&�'��`�������䋯��&��=NK�uܶz��+��p�[�l?P�yHo+��
��'�_��ผ�A��_͡��w�H��)�}m�C�g��}��}_��s�k�>��V�Ɓ5
-SزXtË�,Z�j;qxN��k��v���`������������}fG|곃������[k�u�U�_������~������{�����({E)��η�����q7�������x�=?���z��7�-�e���[ߏCL��
��\���.��� ]�ԛp����I$�E�w��{r�Uu��n�������M�����{�C�]r���}P�����쏫�������ߝ�������k�:���{0�GX_a���^��J�av����;t�Q��(	�X�c)��k��.͘�����7^�Yg�cBcE�5m���Bv�~N���^ 9����};Q�6M��M�&5��"r�}S� ֽ�'�3]�<z�륑��V\G��,���I^�����d O�4KU�#�ֺ&��f��Sy���t��T��4<1���tI|`MI|8t��Ǒ�E��N)�ڔX_mMf��t@�xp�mٜ�?�r_�]��ǭ2�'��5������30W���c����v�c�	�V4��'�!v~b�!�
r�A����L4ؠQ��۟�g�UԲ?j��T��RC1�C��c @�b�!�����Yo��d�iԨ��`��.1B���8˺Y�����=?�X�ͯ��Z�	G���[���WPO2s�q�.9$D`��یE|�OO��@Ԓ&�`�v��AǢ�kۛ�R���I����`z��5+$r`�4�=�d�K���h?A�Q�dT��&5��,Ph�zyu�������;pc�#�A�����]q�Nٖ 	��Н�t�!��G2�:mc׺���Ȕ���_��/^R/���j;(�8O�Ac�L8Ou�H¯.��]��:v9Z8@D�F�	�#��3Lx������y������\]_�{E��
I�F2���Ņ<���%ލ�a����6g���ӓ�G~��Cp�iҮ�Q��(�>@l��"Ӈ����|��}�����9�/5��Ϲk���I���������1o�{���-��_x����oߣ��	&�s�X�� ��r���T�������������r��ک�@{�1�+>�`����  ����~��PB�i�DH���C��� 0�f�V�b7�>�s�u�d�y�߮���mH)��!YC���~�	r��a{�.iY ���Z�b�T4�ELft�8a��:������l����ѱ,�����!���|&��Zk��d.��=e�Ya-��\�I�c��C�l��&�:`�~A�5{�b�ko[� �]!��؉G?��!�?���\������eg:������/_����
u�)��x��&�1�{�<����������7�_j}]D0~p+!��5.a�x^ю��C1��� �!�b�!>�Xn֚ČM"J�24��H���e��;�ߙiB���GϾ���Ml^���bv��e>;�b����ZJM&!����3i��r~�x��H
M"����y.k��l2H��` ��D5"Pr�����X�1�l�?��R��ɷ�^�В�zM����z��FX���\�W�h?�\..�r.�u�H����� ��DF���L��̉%���T�+G&n�$��u��>�;\Y��d����_�I;��ׯ�E���s ���U9�>��,�#K��������W�/8]�2A�~3�'�K��m!᧟^q��ğ���f��57���9A��#I_鼏F_L����Zӧ+b�҉���<��c�fH���ƁD	�N�+��~�����`�C�����������=��Jb��)b�3L �����/��߶͝�ߟ���v�+�,���RT~�^�y��c�����}��o�>�}��� ��~E`�~ؽ�~���}�?6��9n}�
n��k�w���	�� ��L���>� C&6�Ժ6i".��a^f�r���l=�A��, +C�j��q���[ە�h��d��q^p8�R����YU����F��s��!�EA�;7�HfH��H�e���5'g9Y`>`|�W}-�I�����L���|�!�%%���A�&�� N��-��cPx���7�k��t\�7�D(�ぐIj�Q~T���q,���3l�v��I�>:!C���?��ִ���@�VωI�/��T�ӹnkL�H��h]�튝'� z}��L�h�	x�`�W.v�gC1�C��b @�b�!��,�@G^2��NF��dL��P�H�dl$+�G�|�*��7�����o�?���jK����Nc9�M4��犀]lH��=},O�>s	s%�톯C`}c�]X�v�ITh	p���-�$�:& !3��u���7/$�x�� 5���K��Z^�_H���_qd�}�I�f�$��b��ɑ<~�X���#�|��C�	x��7O$�$2
:����Ӥ���H��=��&����H��"��1C���j��x>;&ӣ��;�/0I|�hq�����{yy%o޼�����S�Z�u;���(�BbM^7����+y���q��Q��ރƑ��,�Z���J�	�/`�Xb�ɫI\ d9����q�v��-5,��9=}$3M��+�"�C6����C��?xa�v�QNr��Rݫ �tU���#u��>�k�c�ۗ*�K�%�������P�U����v��h~�s�>�su���\oݜ~��z��?O���_;���ȅ��ˁ�U�^�1�k�]@�����̹+:�'��XA��y�5l`1ibE|4���S6u҂��Xuk�(a�=��c��{�k����]��1
z�􂯂�T��6;��{Sp�Y�E��fC�-��0���ד 	�(�u�(��A��N�2ӵ&։��B��Mɱ.úlj���vҵ��\߅N��|O����M��G������J��~�!���<����8űHM�,
��E���������5���� ��Ҳc���^4@kd`��g����cQV���l2?��/�X�� @�} �{�B�b�!~1  C1�C|�X�g6����Ս%�^� +r����z��֙KP�.f���8_�j�IQ�LVS�;�i�8�M�\Vc}�l&ǋ#9=:aҹ,�d| ������dd]cM �(���ϖ>0BRM�JM��VA��t1��&��V�l<1�Z�h�	���յ����t��G�&�yWW�iYC�X_Ƞ_]]P�	�_|)O�xF�d��8�J)�iѐ�Pi2���)��X�W�ބW%��K���LnW�g�_YwnY6���k9?��x����-3��d4i�z$a�IZT�89�8Y^�Z��իW)��LhᾆR;cR�����&��-�b9���Sl-�^.����e�әnob,��j��F�`�T���DZ7#v��Yd��C|4��{�����&vA� ��ҝ���{���D�vjx4;E��ü�p�G�ύ���/L>t�B�A��m	n}��SP�B���[q��wIy�����P��f�yM?��538�|�����$S"�^�n��]��oۺ�}U��7n�Ԛ��~�x��{�^�(c-�A���`������y�x�����lLџ�u��Y�0Ӷ��u~�,��(��F�[t)���,�p큵�[W1Ä���,���΋�	�m&�[�`]���XKھ��gN0���.䤦6�����k�����uRB_H�����=R ����1�~�6�2�L"�=Qp��=�v���U� I�na����3%��aM�5a^�$~�^�y|r&�Dס�&�Q����HM��$�jǨ�W��'��c���?'�y�T���<�n'b�aoK�!�b��D �C1��<泔  ��0�v+&.HB���L�?[M�R�6jB~��Z�bxh�� �ˣ�S�(��(դ�o5A���#	���"�"��0e�Y$fЍ�؍G�y��2֏�ͧ�,�Q�����(�0AGAr��(��<z�H.ϯ��w�w��g���׺�#��X�����b����BJ����LN����Oٕ/�,[��-��+�L�\���~���sH���������WL�i���}h e$��K�.��i�^�랳�
��`f,�����͚ۀ<X'EP�JSp�4��N粝�r��ȅP�c;i����L��� �# 0s�(����f���N��8�XI�D̽z��,, )��4
���@���TP�8����&yu���3�~���H1��n��y�S`�%�Y�Co���	o���Z�u�f�{F������� �<�җ��y���C���)�n��<�Hm�c�S�R���9u�4|l��_}���f��Ep�{������{�Q�|]}<iE嗊�뚟~˜�;̏�ç��3�FH ��o�bw�D�5��;��M3��V(���KⱤ "�4'������n�� 4*p�t�"�F�>�^鍙f�lH)�J7�ϗ�)�:����2W�ia��#�1�cDc
��	��t]��uc#QY�aL���i\��d�5߇��1�C�� ��o]ǖUق+6Ͻ��>'��x�f��Ʋݩޯd��ź4�5;�ٜC7k����+�T�Z�+��K'��vPpކ��k9c|��kD0��8p�g��e�}�1a�ˆ>+���sD�\W�l"C1�C��c @�b�!���a����5��6��h:�@�V�t�2A���-M^F��&���v��́	'����Vg�r<?b�y$��~�X�*G>yr&o�\���a��a�a)M�NR�16�4}$n��@BG�h����.���W_m��Ꜿ��܂���4f���h�	_�q C�N��GO���{�K�O�H���{'0�Ԥm�r�H	5��Ik��	��ȵ��1#�,	�>���ٳg���4Ki奢�v&��Y�fƪ����9� ?p�X'�h H�&&c��d6�a�㧏�{�C��1-�H拙L�2I"x�,��Q6���=�3:#�O��o�,�$ۜ�f Pby6�Sc�WK���Kݘ�8Ph�������ԡՇ���ɻHI�ee�����O��x@A̠�C�m ȡ��s�������o�'|N?�j������n �(�����C^'����,��|<d�: ���#�c�5/8Pٵ���S��M�w|A�3 ��oo����s�k��E�=���}5EGF� �!�cn?>5�q�M�hY�{3�]����n�� �Q�N��
�X������*JH���,��LR�<1�ǎ�0lM�!�G�2?`B9W@0�y � Jm����\em�%)ƺ�K����$�c��d�d�7ץy.��F�Ӆ�]if9�c>�� lL�"�xa_i�ZcE@�R��/�6އ5)��l]��I`�cut��s炞c�s3G�3Q��>0�X�c�5��B� �MihR�`UOt�^c�X�!��S���1�u鱌Ä@ 컾����F[�w�&�O�Q�b�!���� �1�C������V����/Zb$?m!42]��tΤ���G��I$
�����:�,��sy��-;�a~�����ɑ�t ��2M�d�	Ғ	de�
����,$UH���1�B��m��1I������=y�W�[��3g<I��&xq<'C#+2hu�x6%P P�Z���Ĳ�I��c����vK9,� k}d�rx�@��ICL��P���:��7��!>3
MZ*�6ruy%�Ř�#!�*�Ir��=�j���=��f"�e�>^K���l2������dv@�� ��1����)�%m�^�/ӱ��k�&gUI�mYx��&::�lMh���Sd�T�mLM�Kaa$ߖ�\��*����8��YXzH����C��9�Ͳ�}6ʎ,�}0w�q]}$�l��?� ٿF�AW@���x���`��=d'�a>���C�b?nA����]��t�[�dQ�����~�Y�~���,���Xt{��8���& �3��Y/~ @X8���=ƾ���ă��� �����뇿�����uw��@5���� 	L댼e�R�
F-�$]5�����1J�uEt,���m��VA�>�2\h��5յj�����Ī��v@ l����c;�F2w�����,6���E�x�2H?e\;3��,+�D��B��)��kB��☺�_?t�FYBjvL�f�` �7-;~��F����K�9]�e:�Q�"�A�"8���XםXן��������R��n�Ώ�� Z�QJv0��
X�=�6OM��-Y����uu��/k�G�d��5`wc�q0���np|?j9�C1�'� b�!����*Y95~!˴ R���2K��'������qXl���G�̶L\�9A���7��]��n� dz4�)X��2�y����f���d.ۨ���F./6�ݔ�h�e<-���Z2� �Ia���� # �F��L1��
e��Dĺٍ����l1gG��x�"�x2�]u��X0�����rj��3oܲ�R`�L&ǒ,"M�8Y��� k���$l�D�2�����Woe�d� �gSy$ t�W�+�� `Y./�TC�2
�MNpf��)��!c�.E&Ρ�7솜꜀	�"�H��q��O ���KF#��|��,o�S��̍�a�>��B���Բ��<����92F����Wd��j��a����H�)LC5�m���Hi�C�q���xcJl�l�,L]��u�6,>8�}�@��ɣ;J�x�*���j9��Gw�j�۟�����P�he=�vov����HW��jz�t5,�Xa%�i�1��J;΅��m%A�.X�@�m�x�17��N�7��+�GP��n�<�f�`�7��u���v�X��эZ\���֣E�h�6�}��!	��I��݋w��=Y�Vn��e���Hg�Li��s����V����}!��]a�I��1��Bz�*?�C�����{�/\[���4�羇�m��|�U�X7�i���GsX�?�v[�c�����=�t���8P�{���n�]�Gc�EE��޶�s
�a��hܽ�=7����4{;��P �ʖ������IƁ����kۃ�:�d_2���гF��^�}��eܿ���]���E<x��j�Z
�߿w?��Ï?8n+({I�.��_�F�/*JX�jcq���JbΎyNDѶ�	#��s�5"�3����vAS�!�b����;�d����Yg��&��~
�1�0,��]��mzt`��M��
�uh�۲��-��`��?z��}a�4�����B�Y�m�kGcE�h��������t���]��@ =�uƆ��tΦ���ȃE&#;��X�o�2M�x��ۤ�u_�����G�b�����s9�����9�[�蟩�y�?���<����?�߾�'����rz�Țn�	��
=�l��I�tĆ)=F�+���:_�<MM*,�̌����y�um���� z6Eޞ�&f��B�b�!��-� �1�C�D!��Q��o�A�����$/��t���Պ�h@�����rI��c2�ۭ!���^ʛ7oh:�@�u�^�lq�3$L4t,
�I ��e[�% <
r�#&�(���M�/�|�K�P8��&�G�����h6A�7���Ì"F�h2��ZM:�,�s��䌅~�/�'���R�����ǭA��3��P�cvL��%p=�0aO��!���Ƥ��I�G2��
���� �.`r\/�4Q>��,Ć�I�&���@BNX�x����@��x<�qNu�g�X�
�`��u��$x�n�-���(��>5��kr`��x �M��d�P_���(����}�<tR`��.5��2�ž`���B���ߦl�q�m!���-��ǽ�￠������<}G��?��]1�"tN��j��U���k�;ؠ~�Bj=@�dd��X{�:脇?g��ؗ���T �����j���j[j�Fn)�G h���A�{<��+�~p-�q�5��\/���0�n�7�uP����2�ڧfx�����w��Ѿ����%�v�~�ۄ5�s�I������{������3�e�����[҇fU������cz���w��i%S	�������0I�L�J������EƵ 4Xef����T 9�Y!uQ�!z_]4Nj
�j�&�|�"JgNf���(ʊ�WX�+� ���PXS��@"�c�\��ߙ�O���a]T�[8�9 Q����L&3c�nu}�Vc2���rߗo7-4�8�Fx�a�)��J3��9}M8�kK�TX���k~׷n&���G������i�]���lak���*b�/y��@�]o�#"D8.EY��4+�Z4��;ה,�!�&��K�y���`��c�`[�yQY�Km�e&�*P�b�!��7 2�C1�'��rMH���_���#��/���&HH�6������B>�b+Ui]��Tcr�-�y��9x|LӶ����o�5�$��z��ܚt���Z�������4QҎ�fG{d	o�J�L�6�]s��9��P�#����$v��G�Dl��'�����{`ޝ I,Q�PYG�7ׄ.�t�Ii��r#�I��Ń�)��"��&���F�/�ۂ�F�6�f���<y���!_���}�٫'�%�&+Pr>)��؏Q:ar�1���O�����uGI@��z�S�hе�R1�҄���1�o�fq�25ޤ�n�M$��81i4$�[����%�&�R���ErL�?V�.:X<ɘ@�su��>Xۻ�0h��㏸������}�a�M����b��K�z��=H�c�5:W������X����Ǆ,���b \��Nб=P,�`�m��Iz��4���1A���v���J��6���}V���~����g��*	Z�`>�Y���/pu���A���<�	�@�`�S�s����؝������r ��� L��wo������]��C���۞���Ϳ�����fڿ��bT: {w�ǀ��o0�A2���6
����`inH���%h=8v>���w'u���;���O�ϳ���������ջ/�V�o������Wo΂ޫ>L���-����q��o_X��~7�n>x	y�_Wi�G���y}��K�0�K�RxN׏(���A:��s랜��u�V{�)i�Ϲ^r�v�nꝽ���v+�ab�ᡘ)n]XÖe�u-�B��!4�w���k���$��3]�-G���?Ù��I` O��X����r�~s3�C�Ǝ5������(�� ��t�|I�y��N���~m¤5=	�t��t]��/>�����x����:e\��&w����gt�iȱ�V��K����%h��`��`�����ϭl����C1�C�b @�b�!��,�o���i�3�T
��W+�������&��(��&|��b��)2M�j&k��\��f�	�T�=���p�'���Nco<�@��B�f��fC��tb�XZ}d��jC��14	M#��KW���`�����ҽd�X	l�
4���w�Q�]k��M���0�T7Qf[{��0���8����:�M33�}@�(xLo$�yemm�4��C�伨8_f��а�K�M�xHF�Q�S��}�G��/KjGkb���ɺ=Y!q�=�b�c&sm�^U��c2jPX�q����5�����D �Wcn &5Kh:�q�C�N��Ai.'�ga���M#1I���J��w<�}��6����e����E���`�+����{Gf��w�z�UqG��MP�kZ����/��F�]�'���\O���О!�}q{xЛ�w�����q�{��O�]Y��cW6�{�Cž��m۾�+�DwO���y�<��������A�w�{=>����=p����G�ִ�Ybf���3ǭA��N"��,w[ ��X'`���}���~h� 4�uF��z���
k3�& ��p-�� i�c�&�}xg��a��;��C`��i:�42�Tɨ����m��� �J|�
 �r�
� 5��KZ����N�Y����� @��?J�f�O� �ƉSb�P�!�\R⵰F�b')�xI�5�=`�I3���٘�Hu��]:1br_�31f�	?S[x���m-�5^���B�!s�����A�H��XRԺQ�6�1��l�a��NF8����ןCA�!A�!�b�!>u �C1��M��\A^���b�|��%�Ɣ&��I(ߓ���ך�m�q"!��8�ӓ3MG�!�c��GO	 �8I��u�e"8�cC��1_�d>�H��>�CM�PLgjL5�� d � �,XЬ1q�GҚa�̹-�%��J��x��/�@�
%tRoC@W��F�N�����2��|hE�}~m��$^�x!O�=���cJS�gc���V�����H|�>}BP�cQh��e�0�L3�Ob�ԫ벬��Y-tP��'4�d� fB�C�3�Ld!�;���L9��Jm�2a�Ϧ)��,������1� �$Ѥ�JK�/	;�Bm<z�@��9��;�����lhE�=i���ݣݿ|��gT�7O�N*���n�]��~��V��n(�����l�*s��u|��ߦ����k��M�����y�������֣C�7�|� ۫_��������Ʊiv�켯Z�Oy��{�<n�s��"�'��`NcŨкw�x��
�7>���wmg�/������Mv�>���_��j�`�;�����oc��筐�}O��[Pϐ��=�����׶��4;���k������8=aw���yOD���3pE�0ڽ>����W�s�m�(Kek�������w�������CI϶�y~��#I��F�\��,�e�5��L��<���Q���� �\o�s�Wc�f*�M%��E�v�Q}| �ot1�T*غ�D�ɘ�0t���:l]�x�a��efL]WE��Tb"W�ǜ�Wc2�= M+��uf�QM�"4�0l�<�c���Ͷ� �33����Wut�:��?Źp�1|�����"f�Sjky��.�~Bcz��3zcC�G������뙤���]<䒨a�U����jC1�C|� �!�b�!>y�������k�."Y-kik��F)�����RF]d0;��^_^�6�yaĢ�d2j%�,B�d��N�,�ysο��'ɋ�&rN�ɱ�� f�.N���;U#'_ e��.�*����+MƞQ��f����Q��Mp&[]c A�K�+�:��D|�D�o2*+Zs{�=��#�+��� lB[�}�r���Ͽgr�t$�x�h��d��G��7ߘ�&�!�`Ɯ���^e�|'�MB����r]��Ԁ$�`�@��0��xa�N� ������[m����ǔ���E��8���9={$WW[��L�k�	F�B��qYoJz�x�<`����(a�ct�����)��;��ō��O����0|!�-Z~�@ˀ	��S�W�3�N��jg��wy�x�k���"n)�;&�C�z�о���dkWgA�gF�����}��y�cB�9����HAz��]~^:+x���Ky��_=���y@������s(��Eﲭ�`�a��j��(��ͧ?���&��C�_.�{��q��Nb���pd,���Dƺ&(j��b<Jɳ�LG&s�+N{-�V�C�&�S)�(i:0�'�6����b�y�A��E���le,��Ej���Լ�"w���C�:�0L�}0���tn��q�봆�!Y�5ח�x	�[rMUs]��>�<z�%�3����ng���II�����>`-I�H����QGB&��͏5�`�'���C@n�IK�D�[����n<��Qэ��S]���=��E�Wm�[[�dc%e����hX��A�C�4E���������-�O�f�]�C1�C<, d�!�b�O������D��#hCr@�6$x�uF�#$;qR�Ya�HQ�ry�����ʛWW���k�$:Rv	"�]������=:���0��� 4��WגW�*�������{����R�d$#$�!�� Q�R0"��&q0��+'�P5V,-+�~�4,�iaE��X�r7���X�v��7��K>'��:C�b�_��%H��Q���
������CY3ϷRj�jr�8�db�A��E�F�3N�h\	6$���qƢ����X�x�L���f�[‵-K|��6���r~!;� �<z�H^��Fr����������X�eD��RX������wMcTҶð+R��]���=R�{���
���������fDߍ�?�+��J��;��g���ʛV�	A˖�>qW�61�~7|أj�W������D�c㐜Q��rye���?�Z/���)��,,�0Cw<�V�=xG,6ӇA��FWUS�og��e��@}HӴ�F�}���{Ѓ]	���ΕgU?�<{��۶b��M{S��g�fow�������#����{�}��^ͽy"�_NNj߳�c���������~rD�0m�j����}�&c͗���y����������6�7ě��>�W7��wo�>��g���g�z���qC��~��n�QC*�nޅ�HQ���bI�o�S���M5��-�9����5�-q��Z���ۤ��.Hs�(D$`����v'͛�7z�N~�	������RɈ^d�['���2���c\��T��y�~����j�I�6,��Y#;&�4�e�m)���1C���O�_%еolco���O�-[��<A�k8���~de���y��E�l���U�����&�Tp�?zLyZ3/�8>�ÎǶf���ޟF��)���4��L&��%Glm,�B�GS4������!����[�v;�_WF C1��� �!�b�!>�X_���i���r�f�W]#�*��OI'A�	����O��"����ǶWK&h��	�f���b�ύ	��)�0b���F!�~�x�ɘT�Q�ֵ7���Q:sE�a��8&��H֌͐���iC#!o��7��dG��l�mg�$��Ke$�H��$ sܾI ,@��X�njj+x ٷ�<�'O����g�<���2�}�h2���8b1`�^��� ͔�2ߏ�&�q�aǠ����f�;��v�%�]�Xa��
��1'�6С	�v#e`�:4�g�r�Q��K'$lc�кB�m%�"�\_���p�c��NE�hC�=4��L�QDm�����v|K�йy�~H��_,®0�A�}��Fv����e��_ڱ�=����v��s�# \?�u�W�/��m���?F�Gи����n����Ac]'�4��k'ET9OψB��6�%ҙ�?l���2�cq��!��~D�y����}�)x?��sc�����g�}��ܾ/e��逰��-z�i?�;����v��챇 ��߿�ޜ�u��A>��g���Bw �A����?�>&b��;)h�p��C@4EL�,8�k�ҡ	��R3��"k^��!1���[�?���HAԮW�6$83!�C6�<ۛ"�_š3YױD�����Ŋ$�<�E�%鎯\5>�(z�Pʬ�d�z4��K@�t�=3���{s�}1�5���ґ�kay��w��2ɪ���������X,y�����: ac�����0�ˣG���'2�O:f�FcS�طe�uldic��SkB�6�2Hsձ5$a���s;hz	�^Pe^ ���w�!x��)d�!�� 2�C1�gh;9	��f�W���/����|�e�N6$e���>�eQ}1_H:Nd���F�U@��lo����j��)�xbE�L��A�)G�\l^!�/��SSF���BV�L�#��,/�'�F���4o��X���G}�ȼ0`(���c�6�&��iC�
��������h�(2�s�8��s^�Uy.)M� (�Lg�l6kv4nsMB��˿�����O���s��n�`�(����`����&۴`����2�A�xJV�t1��4�K\�$f�u m!A\G�8��0�N�F��� �i`)%ke�Y�x����~��ӳ�Vvρ	�$����ݛ�MFVP�L@��Zf�HN��4�|2:���닗���KY��q;*�X�<N�ӌv�S=?ꨤ�f�SDn��]���>X�#���K���u�CbBJr�_��C��싁��n�صv&�8� z���Q]���ͱu�;)����Xձ4����X�"(=TV�6�q;W��KWxAxMn�L,,��P*Н�[�<�"W�6V��"��'�aգ�-��;���l�=�/EW�4�J�����(�a��Y��gC^���޸�G��DGV8����w�7��_k��D�6W6�Q{N���\&ib@��_��Qc���"a��Y�d)GGn?}Gk�����Ǝ%�q� h,�ƶY���D�+
u�$d���<������	;�p���c��V�CVd,̅,oy�������1Oj8�X�ds�V CEQw����=d�� F�M��>Ď֯���g��k������z�;�Ь�Lbl2�⼡�^W����>Uۼ=V�l���Nḅ��Y����
�<�8��y��뛜�p�ʾ�\k�X�M+q�?o�Ȯ��1Cpm�=��-�&�n�L�ij,�$��qU��g�u&Ɣ!
9f2K0�?��M�f��8��p��}���,Gaw�ֵ��Yg��o�{�~^��Wk�T�_<ӏ��~�}N�J�yP��$�t�0^|o�\��{��/q��k�a~?��=��i�i�'v�����Q~o���'#A��&'��d{�v�$u�t�{̿.	m.Ѐ����~�ǌ��a'9��{�C��x^���lx,���8�]�s�{�5��u�/��}v�t�(p���qlP\�:��G����Y��ۿ���s6�@>	 �H�_~��l�����Oryq%ח+�L'��Yv<���ۙ��Q��~׫_�5g�������k�\��&�$��?�Zg�O�:6��x6������B` �!��~t�y�ݹC	��L�ׅ�{s��)�����^Ƭ��N�#���75�@��<n�1�&1ɬ���L�l�ʾk���Y���h$��̎힅u�~o����s�F��ų?�?4$�<Og3�q��_,����mM���k"~�U���z��	�w|L�+����Idk/�ͫژ���T���!�����	 �uJb�!�� 2�C1�'���B�خ5��P���Ȯ;�2(�C�7Մ�
�	�</�A�(N�$��n��	���>d���r-��Lf�#)R����\��L������-��ӓSg��3�c�%���1���2�dM's9���T3M�XDoN��������@�-%�P�t]y(�F�M��$b�k~ �}�Ay�]Yٙ;"�C�1VA#��Z�(R�3|��0}GºҤo�Y	r�8��5��� ��z�";�=�M	4��ФǼZ����^QE!�Et�ti�0�vA�'u�!dm�*�W�{� ����M(ƹZ�I�����c��dd������Ok�?arXad,�L����7��w��l~��gu��/�B��������4���d_j�뗵B��P\�(��`��p�� �HW��.o�p�b��B�(l��(�m��h��A��Io��nX�BUC��!�xi��-Z�;���雧I�ݍ���9���u����@�뚰�yl ^&��%�X�aQ�
t5	���#�Z�P��D��;�Q�$`�]P�]q��e�H����m�-�[!݊ǘ���l�XEA�E���bh�㷛W�u�;g�S�
됾+��
l,
��a��<�*L��x��S�v�6Vg�6�_|�|����t�y�"�;�a ;�3w�
M3���d�9���1�\�� �U(^׵+��1��jf(�%q{��q����TY�4�j�� �+	�|���;f����~���[O ;���,�|���T�5�9@�yHyB���{El�;�G�ҋ����'�䎉c��l��S��Z�� F�_�����u�������s޼���*��1��0�+��P��u���-���c�q�`�w��{B�?�4�ȑ��~���=@�NB�k��5i��������@��E���q��2��uP;3��]��!��p��N��m���<nDq.�dR�>�/"׸<8Yꍢ�<�����1��P~�������q��V��hM$���{#�|��o�u�{��/W�.��q"��P��rWu�X�Įe�Z6����O�6��^�E��^��o���Օ@��s��6��d�f8����_y��� {Ur} d>]���s�����j��[�a��  �qt�;����Ɗ/�[�ץ�>Ҹ�ߛ�v�k/�Nȋ'�����Z,_ll򮅱x?�Z��]`D��Q�X�F��8�*ː��tľ#�a�,�zo\�I�,�g�<ͷ[=޸�v/���~�;-B�uygt�Wd�H!�ng
�v6��y����
�oךp������ȼ��i�'W�UC�I��� o�9뜮u��M��_a��F��5�`�O��3b�!��� 2�C1�gu�I5��#AA����P;9�[�6�qa���*H���hb=�rq��\]�H���!�0�?(z��'0�FA���˥�iB ��5�$���E���KY]��a��B��$�
�'�{0�6�t��� ,�V 
�<"���W �t?XTt݅I褙j��[P�rU�Y\G�@c~|�ی�nA��,r3lO̰=DW4�HKW˥�DyM����Zm姟^I�c���+����J�����<>=���3!�hMg<r�Ƙ�f4�Y�U�}"j�($� �_���ň:Q���{��ؼU��k �q�[0��z>l����& D�$��e:J��5;�G#+�U�P��ǉd��&}p,���'�JɕU��Щ�W���T�w#p@H���]t�.^7\\�I}:Y��5��oK��
|�c��A1!ۮ�zU��[����1���wmb_d�UW��� GW�1��&iZ��G"mW&�jUe,��c�; � 
Ι�d�<k�@2��q��׽�id�`E4��7\O,�TVH-[�n} Vly�/�����'����zeE;�L̀<_"�YN�� '�h$�n[)��
�A�@|���W��;�Z���>�Z�G�X
tC������X,��Ƽ2�/��q�'mi����ڢ��O!b_Ԍ�\�6p�ܱg�𜭝$`m���p��>|֎���;�_�����LtnK��"��IwI���$\��p,�T�y}ũI�ᘂ(� ���Fl�1�`@�w +�5V���_R;@��}����� h;�Mv�u�
+��f|_��L�*��9=C�C[�R���2 ��%P���@I��ߍ��Ɓ ���{qd��cٵQ�xZ#�ژdjw-�+�K@��!u$�N��[��<2 6�=/j�L�[ �ׂ�[�q�$�a�Ү�PZ�����O��A�������	P<�1�;6XdW�s�W�MҀz���G�5@C�����9'Qm��K����W�%s��ؤ�ЙO0����	8�k�Vb�@�~sԍ�g#u������4d�t�G'c��-��!=$pז�ój|]��պ����o��g�Ƙ1�nw�	Z�q6�RӓX3`9/��+Y�c��*�I��wf.JB^zW��������lM�5�c��=ѵ�(��Ņ������_�0�Ɖ���ȱ�p��G��b(���p��"l�}1����{������wj�#����>�:`�ȫ���<�@�ݞr��q�&3
` �Y�$�������?�?��$;�¦
7o#]s�[�a���4`׸kw��7��ɚ�Φ��2�Sw���r�N�@�̝����|. 4�C�s*�����:���y�qձ�j�,
�ZR��}1�f�����E�f\{��2�rn1�^b,!�^A (=>��`&2�C1�o# d�!�b�O�ܺw! ���Ssv⡓պ��n�Lڐ,ǚaC*	�y	�%����Dq:6��f�I��0A���rU�rŮ��h�\$��&>�^�b"r��͚	�,�u���������K9==��\��L�d$��T�+P:MeR�uo�4tf�}�m_,b�/�s�#�qj�Q'I�8�|��7���#�8?g1�o�ްr=}0k��1�p��8��:%Q�,�J^��R��+M�/�,�(��oI"�����������wK�;�E�A���u?W�w v������vK�Q�d�u�;w5��s�;��� �l�ë%�SJ`��ԟ�fȲ��`��d]\�q[�X�����/����:��=��bM���}����T��P$$��N�����\Ɋ�	eM0V�1����F�ݶ��g��D��Sf�n�e��"�D�8�+�7u��ֻ�&� �ǂ�x���6h�� �R�n��x�l�k�wD��)�τ\�ۀ�Yh�{CU��ޫA��O:���w�]Q�G�u���Y`A�+����!���R�-%Z�g�ʈxy3���P�c��N��ƃD�C�pZ�US�9��l�r[�Nݪ���9����Y2��滑\1�E�?x||�]�;�)K��e�����_�??j�����QQ�RvE��ֺ7e˜^>����?���skߍ���Ϗ�F�/���B'Of]�&!�2dt���[]Y�3���$T�Fq�u���� ��[���y/�i�'#�.�����+�p�(~��qH�W�@x%������z�r�(��]��P�܇D�5Ų]n�!�S� 4��ıT(9t~(�<*+c�-���G�}�r�U�<y�*�>W^�P\���b���{o���$=���]wx{>�c�%��"h�����\fBJ�pF���3;����I���R�:7b۪]1��}����Ag��Ih V�؆ Kw���r�]�XG����uv��L8ր1�� n���VB:Jq|�v��_��	LRM(pWd���{k�qݮlX�> f9�J����B@c�*~��t�7��P�wH����u�[�������|k*Ǿ�ɐ�z��^t�Z�A9�^�Ep/q� �m0�Bä�}w�����q,��)�L�0&��`t}��˫�^o#���v0
��*'W��x0��7*o����j?��+��N�ߡ�osw�A,��ֱ��KQ� ����{>�jh�����o5�7ĸ����[��f�v~�����������0k��>��H���/k6�DzO�ch.�z�a�&OU{�e�>n�g2X�;��=��?�5��j6(�ۛ�z�3��#��v:z�G�{5qlr�'��K��4�h���5M��fc��֭�	�}�����il�O�NZ��GO����C1��� �!�b�!>�@B�.£�\&i�B蔚�I�̌E��b7,��-(�o(����xf�Yө\^\�ؔR��RLHq����G2��r&���0�%#�/�L�~H+e�KVSMs�r�B��Z�&�� �"F^�Lސ�f��Х������t��]�g��[���B;�Abv f�5��jЃ��g�?��|��聴
�A1��_���53��䚸ϦӖk�.	���{*�U���5��)Y*��
Y7覜N',,Ե/���k����NV��̋�
�5u�!�[7��=a"�X3pRS(�4M��;C��g>�`��H���t����i����k��8��*�s�������'�&�W�/�Ug����Ӄ�ߍc��8o� 0��Bbil���?,�5��y��֍�[���Ѓ!8�P(C_�"�BR��#�߾`�ܝ�2~;^�O�PB�/y�>A��꟧ܘ�� {����Y��������5+�&3�g�< ܱD���Ih����>9`�DN��(����������Nǜ[x \^]��(������<�u��J �-�X�t����b>�D�;�ȅ��1���惀���X\��4�)͕�[_ _Ķ���İiH��b���%���q�dׄ�JB�|��=c�@�j��Q`f�UPs�ɦ�D��=v�YZu�28�Ƭj Zf<��/����L`�u{�t/Y���x4�Y�4�Wp,R�JF�k^x�Qĭ���&�������kI&�֞���k�I���>�dQ]C�E��:�y�L2�`���+z�I����Vh�`.���9MӲ'�9䎕�ܣ
������>�NbcU�c�N�ȼ3�x�ȃ2�ctӐ8p��UO�� X���5�f����w��&rx��� j�<�M��]`��E�쏟Y'�r�8��;p�դ��( �9�_��xM4����������a�7�Y�l�*��: �ƍ�+,�$�� B����E��+����b~�&�'��q�69�(؋�Ø��� 0Fë���HR��j��}o����;�>{�7k�(�{�����9� ^3��;��~������݇�=����@b��Pm�8 ^Z�E��gYA�fJy���u�m`�d&[�5�})�|�9�s�,]WL�s�O��g٩������x�\����؈���4G�^nҏ��mµ�$ЂȘd��l�?�B���\#8�׍V��)h�Ad�y�1Kwl�`�F��}���߅`����kiU8����I����;�,���#"�a k'40�X�1�K7��lu��(0;>#$�z,o�~x����;��];t4��9F3@��g��驮/�R�V��j���R�<�y�'�>�P�%�6d+Vl��ڴ����b�[��~�#�u��!�NIA�ܣ���1��kl�!�b�_u �C1��e��	
�''�̡=>��t��Lf��ºkٌ��mF����7��B.:�Q��5=:�Y��Q�����VU+t���%W`9�Τ�k��m"�5��N�u����M�Y�&\`b,�����4�o<��1��7�w ���T��mD��O�`3v���&�c�XADH�泉|����y��߬x I�0�����9:6٪�llE�\�	s�NA��o�z;�͚���q.����:+W��{�����v�UVLB�:%`����������E�:y�8R"&`1)��26��[m�Jт6c=Syy�V޼~���W_|AY��O+��X߇��D_wʂ4:���6h�#۱A�,��Y[�}�'���꼕�4���cv>���<@��d\��=ߊ~׽/R���E�]:�U��(�zE��Q6/6ru��(u>;�B�'D)'�����}'�;xQ�"u����v.�h���Y��X��q+d: �X�ۤ�F�W�DM�۫�\^^�|��Kn;�z�Y�B�cH�HF���c�W�y}}���������E�:�������\F,8�Pٺ�o߰H���c9��t�~���D�����13�kw�����x�������b.=W��d{�݋��<�_|�U[T�E\_̧�c���x�\���b�>jǼ��_{�c̮��mb�Y��}Ž'Mg݃.�2���ܔ�����\h�C�LȒrs�B�"p�M����,��ucWL&�y���� b�> P8J��Y�����8��c���\_����5��&�)Yb�+��|���������K�$,����:��|4��j�������E��������__���꜅̣�9��U����=�h8#^K)��)֙��F�,�'�������:[��\:�)0y|���kp�����C�k�ݝg<�B5ƃ�&����η�d1�k ��j�*Yn�7���lf>Rk�Vqޡ[ ��{�I�w��w��ڞ�H��ؙ��2��LF��O ��Āc��2��W��y�Z�3��\�7:��c������������1ޔ���.��5�"��.Ü�w�]gU������u�z'y0�Y�s�8$<Cl��d6wsif������b�ƬQ`��eA+��Hܴ눦��|�k�*h�} �עj��Jv�vk�˿U�/�ځ\��Xi�^�IdRx����׃jY��e`1���Eu��	�?ʜ9@�1ݸr�;$�(L�y���yi�y�̾��D�������W߲����L��c�����&�������� ,M�
��V���Ԏ�5��c�}�H1\Oa�k�(�5�a\����U�+Y(�S˶�@4�����G;�6�>z�:�hIvnݓ���+� !�<۸��9��S�&�XI��^������ص��6��"ȓV`��O���}O�Ǔ:��|o�'�H졈�'�E'�����O�6<��d��� i��I[�ܭ���(���za��9F�K��(�89�������A=�k��MZ�@��w�k����1�C�ۊ b�!��	04 Q�`���0(g��&�M�K)6��A���Yp�KYg[v���b
�(.���k�TA���z&M��b2�//���X���Y�CJuzv&ח+�1Ht!SVH%)q��"ID�	�
@��D�v��rH��� f�h�.ݺ��'7I�	�$;�	k��K�뢷��H�,����d����gB*�c|o߾��&���ٱ�S�!�[�	����=t�7͖�����7�O���	�7`����r6�[.�cgb-;�HT���.
	^��M
��rљ��`P���c���0۲b����L�M."�x6��W�&u�m�H;�I���9>{$��?�ƨCe�ql�N��
8!������w�I��i��YFrd	��"==��r�r�{{"���Dv������"(T$'�yx���3�����0��2#�͍�����3?�Ғ2FЂG�����<�$[�����ϲKy���4�**S���䗈O�z�7������;1�����8?�����C��I����1�Ɏ�ӟ��Fy�ܹ���%o�L�M�b��ק�z�(��'��mc0�q�亐L�Y�"ʟ����A��l\B���B���f+ERg�8V0f1��N46�����Z@\��`�!�.ҥ�g�d��ϒ	T���vp���\!����;Ӥ� ��P��q�]����h蹢SQ���Kd��2���Z�z6�k�����~�>��33��$�TJ�u�����E)9�P��m�~�A_⋃���2'.�R,�ħ��l�YN�q�9����v@������Eg1P�������<���FGDV���`�%}�ĕ�Df����y�p&R�XD֢�O�.����x�^IQF�K�?RA���Y/�un��oD�2f�4eo��Arrsm�r yY��L��W댫�g�j ��VA�ME�\^2!!Ҹ�EBD�S���G�Zr	&�e����A�+Y�F�.�bb2I���B �]�%�hg��c�C�R�u��>K"��Z�����ˬ��?�X��ƃ���=�"�����̳zf�ɚ�r���	ځ��`��a������s��H�� ��5�Y�z���4�e�n�%	02m2��6��+d���/���G��[��
藅�%2����{��.��S�`�t�Yf98�����]�����ɻ�LU��l�{�B(_k}��\J�>;�B�{Z"��4e�Lm?�p�'���������99"
��V.E��,t�%[���-�W]���Hr��<�ⳗ��qڳ��Tb�1���p�̮�A<[߻h����ryH�l���%�7)z֏��}��Z?�d!���P�)���b^\g)C0�,Q����%7��هL��V=�{���ӧ����#<����w$�Y*6x7lϹ������(R3�e�C�ћc����*Y�3�i��
�){�RI"?b�$f��W)�,֨�����>�"d��DA�Ȃ�G��������Ņ;�,�;k��{.g"6��T��P�ϼO�����L[ �
	�JR�S�W�_��>Y�O��
{����#��MY�S�1Z���4f���}����p(O�4�J�B� �a��͉A��<�z&���"jmiNfN��˓P�c����OP&�Rً����,m�GI5�y�"[��<��R��b}��d�6eS6eS6��l�MٔMٔM�w/''�t�������DE���0J0�E�1�|A��A&���"`[�����X���WK�Ӑ���*���^W���r�X
��;V���~r (աp���B�?::r3n;_��_���d�|�*�O)#���������K�>%7�T�>�����!^<>S�H�(�T&�+EEsp�8 ���B���#t��Q'n�.`,(���t��y�R�u�etH_H�1"����J&��e���K�d��\�Z�Qg�+��2M����(n�]��]~@���9���* �|�*u��r��f�����=���7
ȈY�n�wV^�ީ?��{�r�r��4b�K���YZg����0,s2$����V�ϕ�i�%m�/4'��C~��Ѳ+�̓��0�6������^��I��V���ߥr	��4��e�()K
� ,n�j8�/����O�L�Rԇ`|�f�~���A�=R��������&1�v��01�l �(N4�'���̫���kX�'��"i�M���%Z
�s����H��O�}DC�#��K�H��>[����Cy�f�%�ׂga�H� �(������<�!sj��> �:�k�����G�DD�j�*1:������Y�A��y�9t�i�Y�����Rf.k�����q��y�d�z"q3u��b��V: �/��� �%C��,��� q*"� ���BH?{���\�H���s��\���y��/K�� �7�x5_K��6�*XmF�~2�ŃJ 7dV������ZS��$������B�_����^�,9�������1�~�1����莮��t��	|7s��1���;�q"����;F�;1��d#$�$�#�'ۂu��n�v��(x��)�<�� k����Aڟ����~�k�9�sE�w[C�|��ݳ �� �]����s�:�~� ,yfBo6s�'k�F��� Y�<�����byW=k&� $���zA�ΜPtR�	2�1�-ݕ=4�5o$�U$)���Y}N���A����8��D9a_R��̠m��*���H_�~#'��~��U���u���j=��g�Q��gV�r�yy(����$�@�6ϬD\If����y�}t���=}B�x��|�>UE���q|d��\�i��1�}~��.�D�陣��i���x�)�dUP�kŞݚ���oMT
'�<��ѣ��(���c-�j�×��&<��˰�/�F}'���[��k�z�y�k]D:����Sp��!&'1�f��L �b̼���I`���D/ZBİ�y ��_X{O��?����n<��g�=c�l̜_�Ļ\�\���m �S��J��#�k&�_)�u�-HT�<{s:�����)Pw�b�2*�soA~Z%��+�}���t�g.��g�-Y�+I��I�ф��i8;?�^�R���w������8�}l�q�d��bA�R�{U�,�q�F����G9�q�)��}P�➵/m�?���<�lʦlʦl��M� ��)��)��7S>|<�����ɉ�8�rO��؝��j%�} ��t���}�r8};��4��'A��J��T�g�v8&�y��9���]c�P��04m� m��F�Q�ً��j�R	���� |:=����Jxs�k߹СPf�+�8t�� ~yU�f[�*�!�`�t���~�υ"(3�>Q��E���a��A�l�����N'�����6�^\J�Y��4�A'd����Dd@���V�3�jS�ؗ77�r)K�#��X�R�  ��IDATyyB��$�6���E8��du^S���ݭ�Y�:��!�4��h��x4�|�H烃�ж~^E�R#��j�jEI�,�I�u����m���
۠�A ��������0�Fs��G�����������Ք������а�(W���7�V�u�� �ŝE�j�Ƌ8����� ��� ����F��+�� V^!<&���l�h�uhd۸ ���9�[�6�.{e�]�ڠc�1
�꾀)�.�	���Y.��Z�A�4�O���^�å5 ��&�͉�v����#u�QV.��ZF�PD�v�J�=�����@�V�!��7 $��e"i:"���(wT�:��C�y]����%*ʶX��.����"3 ^�v�g��W컪���}h��8��lE�C�p��Hvľ� ��7�(���Q��D�Od!�*�d��8��R���j�io�V��`� ���J�T+E#jk���	ͥ�r@�P����бz��qN4e�?�'�^G��>�̺Z�*� ~��ȯ�]B�uGF������J�hʛZ�֥��/����|l�z��mo<К���q���4�tm�N =ڱ���*�4�VN����g�@�BN���*��ȴQd+Ym2�<�m�
zY�de	"��[�����6����$�L�n.��	!����c�&�\�2���o2���dbk�g��We��Σ�/��#�ԕ���2Jڹ��Ga;�@��&R�~���,��.\��Z��DT�i$��*��g�,2�ͦ��r��=���:Q�{� �%'�i�؋�f�#n!�<[�됱6���0�>�,�y��[h����U��o6�e�e�Q�a���f�|$�4�����_��ۻ���9Ad9aY�l vQ�(��Y�|��2$���.�d��'C��`�21P�w�³��ms	�:�+'���(96q@�}�괰�~7�x?k?��f̣��@ؚ�v��d9]�i�3�
ԭ�x�0Z����h0�+qP����O��ܥ+E�Q�����2����HF�r,ݫ��+���������B	��;XӪ�4��7Zo������ 4�M�m�`����ţ/ja���/��*�Gq�g�BY�k'�
����b"��3i��R�{7��3�d�g�}dE�N(N$�ec��7�A���	�_�{�$����?��ׯC����ۮ]ÞG̟��(����.�3�k���JU�� rlHr�Fa�=�v����	Iq)���H1��y�Jx)5�`6V���&��c���E�V��-KZ����9xV��w�\fm�J2�s�ux�� .�]�>U��(���-8+y��E�L��SHܟLH��= �.�����L�/��PRQ�R��~yqM*��^I�#C)��6Sv�2R�~A ��+�߃���R������;ûP��E���t·�Kx�����p$�:HIe��L���.d�,��	&I\.roo/��y���c���p���'z�e���A����ր�v��Y��j��������RW�"��)��)eC�lʦlʦl��D���(�#���_���������}�)�����9X,�aL��G����[�æt��M��%���"���4���T�U"��\��ap,���ө�:|��Ƴ��AD�ժ�0��i R��.?�!j_�n�R������Q`�M��2Qϱ^e�{�G@���O�{r�	�C�ONN���^$=��sɎ����?��B�&�� ��q|,� �m�석����#���S�J23���U�#`��5|�p��|�>}�{;#.//�PG���1vxu@T��T� ����>�ֿ�W~Bd޾��5�c;�\]��~����Kp4��P�>Pl�Cy3�skg+\]ߺ� d��st���d����k�ТGN��$�Q����Jx9$�G%�+�.38�e��Y=".�7�#]��j�9R���� s�6���L&�.ID6H��9�w�߸�.4h�G�w /$�޿���}}v���?`��T,��is�਱��:җ"�;/O��`��Y(T$e4�-��������QLm�*��x&7��5C��W��"��2f�!_z���S@tԅ����ӯ��xM��vߘ��kM�Et΋!7hG�N�?6�!8r�R�&����y:�-rv�^w��hud�fQ�%D��z��XE����mQ�����RE�f:w�EԹ/ɧ� �2и�!�J����Y.a<�*�F6��A�N�"@�L���'Ѯ.'U�]K��\���HR =�ӱ�%��5^%K��e,��"����v�%	I�~i�~4o�+�=V��_Ķo8x�,(�cf��Y��u%=�$u}xJ.#�(��1C`}�$� __�_��Һ�Xil�����>V�k��d-��/����u��3��/ id� ݈rF.Q~Ni��K���IYd�X~��gu�!�WTu�Eٻ�k�#��l�38h�F=���/�����g W��}RXia�О�,�X��r�ĉ2�l��0��`���ڀ9�!څk��4A�D��FB����S���ܚ���Y2�f]���'x���P܋����5��Q�M��'�#��Rs	!��~5_.b�eI��=�Xe��Ĝ��s�Я$5��^. ��P��� ���s�T� ��%���v�;��3�4�؏y����{�r�eK�d�^������r�H��K��3��ʥ��A��b  �cI1F�G�ϗ3���4�ꚻ����T�T�^��M���kؽ�~�y#��M�Q���˒`��}���:���{�e�2U�D�_.���Ha��*�l5���(+��������r/H�<;E����t���*�P�q�L��2z��QH}�jE��dw�*�pt�0<��Nϯ4N��O�R1��'��%o����:�?W��2�K뒛ˢO�d�撧+y�B��o��Uk���]�=c�L��3�Z��R]��Z�,[�N ��h��fl{��F A3T NY'����z�V
H�ؾI�T��3�5���g�ekg��b	iBIY�1��Ƚ�5�E�j4�n?4�U��ٳ��ێ���=��$mZ-��
1S9(p�Z�3,2=�N%f�]���vn�=e>1X�&s7/����e�����ܙ}~*_'�;�����	C`�h8�s��ō<�g,�<Yx&U ��'�Ud�oʦlʦl��g� ��)��)��7Qno�C�]��,4[����V���ͺT��E�6\.�&�Q �)r+ϭ�y�H�p�����FP7���k�s�  �s��$_��iy�O/��(߱�At"��ɴ.��������vD0
Ѡq!�fI`�k�� 
�V�ʨ�z��V
4�Z��p���=I�#e���'�ߝd�M���{Ն�Q�������=DqJ^]��~�r�ڻ�f�����$%��ҒG���w�������?�������(�:��3&�|�,nܛzD'�"iZ�J8zpF����8��3�T�}  х��<��oH�@Aq�����wwt��-@�2�-�<B�#N�pmcI�������~���f�e�d���<X
.�XCtm1q�� q���Z�K�>��Ȭdc�T��Z@��_��At@e��^�.�����O�V��������� s�����7ww���%�[�� \�'�%S �DJ8(��I@Z1\�.%��HJ$)`�$�����x���qK 4�S �����=B�V .�йٜ��'����5m-D��R��6�ϥ�cc�#����2[��-E�+:�>&���%�>�2�Fˮ]�xty�T������6Oz��"������~�(�k%bQ��3e���B��fʳ�Y6�ÉI x!ʝ%���:1��@(��S̉��� `��`#�(S�@A� �<!f�
���}n���g�J�=�:c
��1$U��U�K���D&]eJ���e�#R�yN��b�ܮ����B�BT4e[�*���9�%�L��?HRBE��hTͺ���8sd9s��"�I�"� � �J6 � � �d�y�Gn �9V��4�e���sO�CԿ�$�T����������W�����+
X-�ߊP��L�?Y��u�n�>��w9�T�wh�V�
�ےt.��q�!�T��ED%��rI���OD�&�2��m7�Q�j�aI����,��9S9Ĭ�T[�=�>���Ϝo4m�uz�&�<Q���@d���_K�^Zr���\rPA}��+�LZ�+'ʐ���rS��D��
rfe?BJB�3�b��,b�u����X\�/H��B�,�F�8���^V�{���R �����^I��$(>.�U��ȼ�OK��cc��L Y,Ro�*[�[�Ƭ�1�y������Kd�UԦzV�#�euH�
��h�e����ɴp��f�A��%}����,��r%���j���Ϟ=/y����j�p4�+�'M3����ç3eʜ=M�c����b��R|n�i���])�I�3U��`_j,� ��!"��Ƙޯ\�R����M1[��uE�L:�����k[��6.k"\D0���n��%,�ɒ�:K��Jc@>MIEYhdI�~��m�@�� �Sп�)��#�u{� H�1���+�zӳ�
N^D�^B�D��m� �a6+`��ޡ�sճz=�[��<�Z��#onn��0�}��a���5_Nmޔ5�xN�z �������)���k=���xmu;=+�ŋt�|���W�<ڷ�������?�5Ǒ%+��t�,�H!��W�r�{���/^C�Pa��I
UI��J=ȄԳz %������(�"R��'�����{�����W���d9��*Zx@S�� ��h�<d�J�4�����	��)��)���l�MٔMٔM��)��������p{{%@�/�!��&�Y1��90Z,����D@OQ���#�y/���"8Ыo���T�d�$;��pk�IN@)� ���J�"(ȶ�N��*�]����B��J�&��ù}��gM����T-�ޫ��s��$#����۷���?�㰍�ևO����VK��Ib�~1�Yx*�#�G�u�������鋤A�D�Vhb&9��K�����h��.CفJI���5$�c ���rHI,���P�3�6�����A�7��$+8hg���#'iO��LEdJ&RX p���E>j�FH�%I?�����#�(�ǇH�R���/��cA�	_�eh�r4�V���=�e~x�ƚ�'��gaM�Q��3C�$(G�U�٩?R?D�V*�6��x���Cx����;���~(]BC޾���8\\߄~�I�������[.��ײ ��<u�!t�C�(��9w��Gk\�N�n?ab}~a����5Wvw�a����wc�,4��Vh��(�0����Z��X��k�w��9�߷�xpPId}���2�V��P-���/�+%ל�G�KE�H�@(*
���r���ZS�	��z �K6G��Zq����n�m:��3n���� L�E6R_�>H��iU�	�����MM���1l&J^�IvO|�aP��e����A[h�KS]���`�}_���I���j�ql�r)f eekgs�t�"�����}M�n=h+�u���z}�Ğj�����ѷ �f�꬈�h�>�Dn��Fɧ��z�V�l훁�J�LYx��	�~�:,�sWX�������G�*'��1��:�L��-�Z �	ϋRe�}ᅑ|ЋF�>�W�(wT���X�e.�rk��\WfY?�k=-N*.II�Q�4zg��ڸ6D;�8:��{���ϹW ��@DB��� ���Q�n�O�|��l%�*u��q! ���O����N��
+��3�uC������ٽ��.�G��ʣ�!�@�Ɋ�T$c�bm�g*���Y�tB5��@#-��z��Td��'JH�;y?y;�$?E���Z�m��b�2�&���A��R5�g���*Jb�T��-*��{�@����>{���R�������ǋQ	�V�@���:*����=��3F
Z'�EP�3�
����M��}�v�t�=3Pދ��2Ŵ����z�Y�I��O�ErIr���}��E���^*A�
No�NJD/2=3�4�+z�x��u���1��~
�|��֥�Ζ}o��nC����Z�߾?���W_}��Old�$х�|�QS�e�OH_x��kY����T`A��I��y*<o�_E�$�� a�3~��ʾq�N26!b�E���$g���ʃHV"��i���x1v43��Dʎ�	�����e2�^3��~�O��?�<Y�F6��3�<��i8�}؍�=��ZiʳF�(d�+N`Z]y�#K�,?�/�o��P����ޯ,�K�"����Xb����=/\���=~���>�}��sr���B�4�xw{GD���d��μ��Dz�P�n1����M�:�9�ҵ��5����pzvac���y~���3)d��֞t��E{�q��L�Y\��G`�m$3�#���=+v�Q��emuh�=����fd���P�"9Y�RyA�g�5$�x|t`���c�g��'�1�}�k|^��-��)��)���l�MٔMٔM�w/�0[����.4[���*���ڿ������R���r���½ �$7���Ղ@9 $"?s�,����+���'OE����MW�e�����h7����]'��Y�to�d�V�Fs'�ZM�w���$@�-E��0��3���H�x���:��D��\�Af�h�ۡy{{�z�vௗ*���<<	�~��CE{
C�r[�n��أ���v�};���~&y���'ӥK�k�PV�F=��\��R����' �ȼ �b�p^��^S��;�ht���U��Y����AomU�v�v���^��n�ܮ�F�*D��3mc�F$��i.}�,�bp���;QҡiI&*�R1K����r莇��#a 5�'s���*�\L�(^�v��B�܅A���iqm6��YS֠kk�iJ9����K�E�`�������w�w�>�������0E�>�t�A�)�~9�X�<��<�n��pN�ݗ!7V)��L��X�.<�Y3V�$�O�&��9��?��w�[?�R���w��U ��;2u��o��r�P���݅O�>H&���t?t{�pvv�#`���RY��o�|g������6�w� �3��:f�����6�2�z� 䈘�}�УN��T^M�f+Ԭnn�����.��Q�9�Y�ܔKi��U8:>r��� ���E����"�& ;h���\�}7O��f��ul\H�hgo��&�J����՝��'�3������%#�o�L�A��W��ص���v�Զ늀�; ��܆�7󍱤h��;��a}s}%��{NB�L�B"0"��a�t&��4�+��V�:@���ǽ�M�ögɑ�e�su~&��v{K���zڝu��u���$��UE���Fvˠ7T]���Z���ڑ�����Z�޽�����Cغ6�5�>����L��"�����Z����7>/%0����u�y?9)aC�kO����YJڋ��HE�zj����F��h������l<�x�^XJ6�Y� �!�{���0U�H]ك+��d��z�r��e�^���s�|����/�"�$��Z�d���|-)���GZ˹Ż�[_k��0Q�d�@�����߲u]F������BV�I��ڸ����o����da1֊��HVN� ]x-R��`I%Ҿ�h���:nb�ok!��$rA7�����-�,�7�[����!p�>�\�P��s�$^S@,2eqޓM��$�r`��X��n+[�	����d"!@Ҵ�6'�7g&���������{�51�tз��=���ZDG����VCk�k�A�g�E}��g�`届�s�ӓ�2[�U�3R@0} �]j8�,k2:���?�g�~�Ztks�y����L��w�Ë/��%��e����᫧Ol�ٽAȒh����f#�̥B��{�!|��[Y���@�/�@����
��ao�����ɣ���+��ێ��u=��	{s�.4n	�`Ow.��={�l&_�b����Q�P<($(��ݻl��v{����F��qp��}�L
d��?��ֹ�P�1:���ԥZ�R��vsK��R���T^
Y��Z�����}_$C�:�=m$R���C��Қ�cc�u���������L���5�?{8k>h���%IC�y؛��[��w�'2Q�?��}W��ao���"��ꩍ��pb{6�j�6�lC�n�o/|Q��9�wO��p����{}���1�[�\�k���Ϝ�X$�����G�����=�u��k5>K����(#��cw���T2@��~z�/O�2�y�
$ekow=F7eS6eS6�?v� ��)��)��7W�9��������f��4v��{P�H��"D�\���B����<�b��z��� ���P)�th��"�>~k�m�-��$t{]��N]K;�$�y�w2ڮ��^'�� �U��@^���X���`����0��T�㩴�9@7�0[���=v������I��:pN��:RG �ܛ�?�8��i���� ���3����H_�t��������I��r?��ޭ�B��<�,���#�;R�������b.SI����*ү������ X�z�A��ە���2pF���-V1�Eƹ���O�K�x>�:���\�j�f�D�#���)�����s��o"�����ʥ����ya�����pm�.��a<9PA��$���e�����>
�$Y��ŊN����`m�S?]'�u�e>Zp�����_|!#O ��o߆��k����çO��㍷���߅�o�
������G'�������:a���o>����Z�ݒAq�22�^���Ӓ���K�N�x=;;�_�*����A��Gσ���o�&�`u8�n����1J8(��<c���WF�ʚ��j�L��d=���=R= c߼y#�/� �@�o�f+�����'��쁽�k�E�)��ݩ���P��xmmmL"�l��(+e4�T[_n_	4B�	����L�� C�R��-Y�J��y���@���g �zB����^U���	D�d~0y^,�^��3�f���6�ϯ��v���cOق���?�t.�i0섃�}�7����y"��k��17��w�~�NQ������W�7Np���k�e6���H�����}]݈DkZ��3��U���i���x&"SpL�����9�z�����/��P��ux�ꕌ�<zhs�@r�Y�u�.����R�uj.���zC�0� h�@���/YS�#}�� �A�߿Q�4k���=[O
$|$�����Çw���B�4� �L"�_Y��m��4���Y@���w����>�R��~q^�~-`I�����#��N}G@�������Sx��I8yx_�����͝Ӏ�6�v�����E�ؼ �c�«���/=	���s�c��V��so�C46���_¹�/��Ç]����̅��G _ekc���^�wqyf�6�l��ce�@� [�쇟��P�Ǐ*�$��l[�Y[Y?X���|��iho5���g�=:�����(�i�����*�.{���t$�ncgic�n>	o^��=S�{����vM�"�믿��6�n��_��`��9���/�[K�9|��I�ﺔ���4�[���E�E8�q��rs��<⺬cM�u�?tℌ�����g']��������~m}���sc�־u�d�@ҰOt;�i�a��(��T)�Sd��p�=�1ȏPr��R��4�\{ݿ����m8?�
{�����+C���{�WY_N?|Ե�m��|}������m�q9������Yws{�9ryq�9�8�w	�������)UE�*�?�|�g8)��+m�.	ҕ�n`<�³ݝ�Ϭ�3�Yگ�M�Y�v5���@k}&�S���"Q�O!�	�$�Ab"���Oz���?�������5V��AJ�"�fc����H�U��M�7�H��	R]c{&a1����h<k=A�rV�m��4��%�E�e�MF�m��!8�|���i���U�XŬ��c�ZY��x�j撉��I|o1>���f�ܰ���%u�{����)���ɣ�����s��2�V�ϓ9��ZY"�kAVvG��S|?ҷ��䒅U��Uu�ggڿ wv�W���-�'��J.ǙD�7���Uo<�JEy��ȤY�4����T�l�e�e���)��)��)��ˆ ٔMٔMٔ��[I

�H��� ���+o:{t�V�2�aww'4W��W���C�)"��,sO���v����Z5�r�Vu�)�� i4 �|��U;�VkE7^����VC���9�Bp}x>��uEBH�;)��h�C�j����O�����@�^�+pH����`o_�Ҡ7���$4�w����MЁ_�@����߅��LѨ����v�'���@ ��9H��vd���$�3��O�~n�=��'���9Y��~n����p 5��N�� � ȼ�媤���"��
p�#g��FvP�٨�K�n?�«�_�_}���"@є����hٽ<z�(���������ahUka{o+4G-v��;@v���MB��PѐAYy��8�D�f�WW������J穀�:�/V_d�N?��痒˨�ɂ���ˉ4�3ϯ\Gqx��4�b�#_H{����H@]��TFϻw�«��_��`,��ap}.�H����`7�|y ��Q�%��߾wם��_�'�Y��̇s����*�]R:1��`�8bl~�{e4*�;QD6�t6���c�?�?��� �R�f�GI�����<�����ͮW��������>Y�5G'�a��
G�{�됡�)��ЉRo4\ ^Qǘ����j�v���Rs���^�޽��?�9��NV06W|?�;8�'g{gG 6Q��?mЉϷ����|����?�v ���]�����#^;v�k[D̗"�ٹ�	���	�����|�K[�l̟���641���!O4��������A�Cfɯ�������jW�Y�˛[��l������Kd���ڌ�����������l,? �nz������e�, )��o_��ϟ��^H�Pn�!!��;Zd+l��(��ز�$��������_<���;�|�����	 ¬3����+���
o쳬W��? �A���2�eM+J)ywzzn�/5ϩ3���˹F]�H�@(��Rp�փqx����_m\U�ǯߋLϦ���K�=�����������=������d�5���_�/?���?��ޒ���m'�^݆;[�k�~?�zi���4�Ӆ����ߊ0�h�?}�TRc�c�����/�䥭�m��Fݽl����Ov�g"@X7�{>�i �
YFa� ���O��p������ϕ����Ӱe�cE{64���e�ӳË_���ݫ�G��eքW/_k_�n�������M5���ŀ�5����/»7��g_�\C^�e�?�(k'S}=B�3�G���˗�������������/�w����x��&��`��� �g�N��ޮ2Q��޿��z���Se�V�Rs���>C����y�t�����~P���'O�į��dY��P�kc�m�i�L$<�mI���g�:�K����.z��P@�p0ѳ�x:W���a��z��ﾳ����J��ϴ���ps���v:9���?��3
��>z�v��z�B�g.���P�>>��}�V#8����i�0�gHN�;�觔[ܿ_$�{Ɣ�]�#�;�A����٧w��/2c�w��!�g��0A���7a��~AV^IdBam�g�����V���N���_��±ի?i�_,���{�u�'�.d��1=+vnu��H>F�>>OƲ2
�n�4
�� ��X�왢�[�
27��Kt!P�H�$}5�t}2R�ݐ�1�+���*�2Ӊg�ȣ����=�H��V?��Ş�Z�����#h`6� ����5���dI��!o2o!�X���
Q�bP�~�^�p�ݿ���A�㑾�l�Lҡ�!�r6u�?y�
�aL�c
IU���;�n��d.;I�YZ�"��)��)��wQ6Ȧlʦlʦ����������p{�Y@1��ާ�C/J˞����4{9�gK�4���P��V ��{�*ٟ>���k�'ƒ���,G�.C]�z �d����?h��V��v ���X�D��;4��� ����#c� �N�'@���Ǌ"}t�8|�_�''�Y�����pg����� �.3pi��ьҀ�u�߳�����0F�~/��LQ�� |0����;F�E��Vu(���u��i�9XJr�`�t u`��T�<�d���&K8���u�Gn`�j4][��S��S�N�`���Q���CI|�ݽ�S�$^)Ve�Ox)| ����'G���U�8���Cz���b���](c{���&D�k:u�x��ֈ�d&TX,#h4Qv��.��P-Y�����ɉXF�"���e.rib�A$#��K�U�XP`������?:�~�tui{�Rv�9���LDb�;}E��jUDY�u{��x��B� �_'v��pc�
�$"ZɆh ����$DS�g-n �q�3_<~���k�kZ�/"�w���0�>��)��&�h��
O�<����YJV��d��
�}�1 ?��,�#��ȯAH"�ထK!An)�s�w�׿��Q�R��W_}-0�@������l� ��}�x*��D@�\Z���8f,m*�*��d���wL�on/m���׫U��{*e��F[''S�t� ��p^��K������ ��# BɄU+j�ݽ�p��N'7�+�O����$f(��������g�B)�o���=>#c�tyqf��1�������k,����c��{t� <�����Dz����6���귝�}eP�e�|�$ĸ�$��f{A��^���HR>�j]�R5�mO��J�8`߇�Z�Xu����/�kH���	����h�T�Rt���%��گ^�ϘÕ��ML��?Q�����>���M��Bw���x��_������ebզd�$u8��NW�J���I�l�;�/_�AF�XN�uV_}�;���e+��Y;��"O���pSd���]�/"��k����'�k綫l��v�w�^���Kxl��Z3��.i�HA�1�}�Xc2��������r��XB�
���h��G6�E��Dcz����܅����aཛྷG"��s�D�x&p����Ӱ=�y�\��L�����?h����PM���7g�GC{��)�ͺ����Zc�����r���6$��������]��>{{q�ϳǽ�z�ퟕI�ػ��Ԙcl�����A���`u ��z���e�3h�䙪c��n4O!�ӤN<Ҹ�^V_���R�嗟���YYt����d�)0>:R����z#�@i�뾳����f�U�� 2�.�'��{������y��P�TWV"���ڏm�#��o{���ke�.&��)�W����t��֫����~'�����.k��V���$��\����"�h
��K��}�X1C�,,��܂���D�9��3�U� �*ҿ�,OH�;���:�g��ZW���,&̽/ �!(Yȕ��8���j>�
��^��[��-��/��ƞ{:�gs~�T������b��U��l��B���az��́�\����ǃ�:A�V���TX��Y�z��_�b��d��á������YVVϾk���r�/���l>����qD���؞���c��{�f-���"��Y��-y`R&����c3�0y';8+D������x�)�K�{�!$	���_�kC��yM�\1�։76_���Q�٬"�
z>+"���RZ�6�qM`Ԧlʦlʦ����)��)��)#��t��? �4��P����!��% �ȳG��c� %�s8�N���3�7��ٕ$W�|r�:�CdS���99\=���i8*J��H0���v��c�^�*�p<�P �Z.����^D�����S����p|���U�29�W�{���D�ف�L��H�\���ψl��iA>!�����pH2@�~�2������h�v:��X��`��Ah"�{H�� ��H04�T���+;��1؎�I~�u��f��,� Z�8�0$�$�ϔ
nv�Q�d�2����"�1��c�=:>��eh4A����i֭ݚ�-��
�Ns����������&󰵕(����~^_�����a��KC>"dbL���R]��S�2&:�PZ	pZ-Si^GvE�^��I�$� BN\L":O}3�� ��*�YKȍ��B;��� �H��B�#]�M��}Nu�=�B|� pB�*& "VE�tRtn4���;��7o����#�~�ltg��� ��2�z�<k�����c$��;9C�9Y�  ��-��@����g��R6���YdtE�7m�����5t�D A�H����w�N̜�d^l��ecs��������[י/q\WD2�Cɽp����&�%�9�Ѝ,3�s�"�
ʞ@f�Z��t��D�Q�k�@;dL� #�߭��NA�����?�/B.���ߕ1��w�	���=��=�3�1>G\ �v�T���=H0@$2 y�v�߿����@�0�!�h3��\���n��aε�O�d8�K&������ݎډz�_C{��٩�զ�'c�Yk�)�7��0�&���[���Ϟ��/_�g���e`��56z������������Y��� $��=%I�A�B�,�.�(B�����e��J�l�`ϥSn�����m2���߽�nm}P��5����J���=3Ǒ��۶���KU
��	dz\FY)�*����SX�����!2�׹O��NY{ ����	 �L�^S[+�zB�	p�̻����Po4���!r�/�.ç���I�ʐ�K���20Y_�Y�j���@d9�K�ۮd���[뿺� r�Ѣ}�$SV�t<W�7�,+���嵵�V�E͉__ކ�o_�<^V���a�r箫�Lk��U�%KE��9��������JYRsU�j���4��R:~��B_����CD��}�2�2���~XH5��?�(���(dYA Ō-2�v��Ɍ�[�������Š�=��Ǐ�t�ds�l��������h8]{�A�\i�ݝ{6DF"?u{u)s���Q����ɉ�sq�)|���կo�q[Yf{�*(H�ղ��T�=��R���h��e>-gKk۲꾴��l-�KI�^Z��v�__��9��+�-2��٩��q�:�<�<����㒖��xh�Q'J�����<�����
d�,���������k���a �/�E`�
�6[���m�`u{""I�P/�`��M�7UdlX���Գ�c���'�H;}|���ە ����ڣ�����([����J�.-xFF9Jrf6ޖ�b�)�O�󼗖]�**cI��I�D��z�*��E.���g���-�N(��(r_da����FQ �f\���Q��c�����Q� ��$�I��䵖�	�qr���ź̼%cc�k��\
B�x/���Y�⤋�;�ͫ>��V�]����{*�s��}6-{V�*f��m@�"S[!�%f��"��)��)���l�MٔMٔM�w/;�����޼~+�������v�ʳ(x ��`؁����u4Z�;\G�2�]�
<>�ߓ,�T� ��Ɨ �0�Z����d$QE�):1�4U�{ g@%��d���{�� R��?~"	$�8x��}]3�.`�\�F�
?���aX�9V�FZQ=0��**���|~@s	�,F�!����!�<
�a��b�Qt��d��,2���\�Nn�&��
�'q ϐ8 �H7;Ezb:w��,'E��*BǾ��$:37�-7��ρв�U���rVX+9�Ұ����Y���*!E�0R]�֎"����i���B�� l��OF�1Q(x6 ���B�M⑨�lH_̔M��'���
�+{�4�?�f `�ˡ�\V�(�LQ�ei�j�D'�0|WZ����L@�b�X�	��}(�}4�C�ޗ��M� ����V�R�K3��>}�b�W��D1,��3E����L�
�B6S�U�����l^����i�wu?�[ME�C F��=<�|��+����\E]n����z)������������� Ֆ�|�3�z��g���C�~�� �]�
����xZTV�X����H�I�v�	"u�兼t*�e�k��c� �c}�� WY��Ȳ���xqy��[D��B�� �Ƴ�J+Է"w����psy!i��� 9�g� �b���[ͦ�%�Ï;;"� �%}"��M��B@"���l("�l�3�:�|�s�:=���e#m��Sg��G��~�����T������7�adkR�V���M�� ��G�>�pB_�*=����I$�n/.�����s��>�-E���t$!������o����||�!tm�޶�-��Ŋͳ�����䁒���M��l�U���m8��ј��=Q��x�X߸,�"ԋ5wUk�|����:?��®W�����w}|G���(����v����w޼|��<�X�!GJ�e�]D�ӿ�7�9�:�V[�����pz�>L�	�@��Ik�7����Ӛh�F��H|� �+Ҳ_D� )�<3 p����v���1���[��4dq�v����i�H�U���'��^/�66Z���y�"?{.d�d�o5�~4½�������o�;��-M�֖g�X��P�L�ľ\���������/����=_�8����OE L2dr	�s�'��V�)2r���Y�\_�L����u�KIo����ߺ$���Hdi�����uӃ�2'�G�c ~��jؚS�y����F��gD�@"Y(�b2�R�*�5 `rK��0��I���?�X_ڞ�Dn��N�1z=& �#�@�	�2�bFƪ�~�l���k��Q���D�/�a-%r��jFP�d�1�\���c^�Dx��yy!9,{��L{ �G����(b�lUV�.��%}�*��(�	���RW�\&�Yq��r٥Lm���A�o�>�ǠD�RY:���S�$���\U�}I̞)�/��r���]8;?���D�=|p�w�a��"��
�G����2;�i����(���a�q����!:�:�������N��s�e\$ٚ�K��tR$Y�=B4fV��3�߳���d��b����d4��elԷ�kQ���Re�(�b�D�>H �J��q�N-�� �ŭ���w���ϋ�����ϗ\��?�&�3�{
�!0d��M��j��C�El��}B�o��MٔMٔM��(dS6eS6eS�f��hb9�w��)z���x�X�Vk�&me������d�1H˷|�d��ޕ�����a�W�F��Q߳�T@'����"��-E�v"C��l<	 �I��yQ�2�ǵf�p �:��-ES���`<r�����T�#:m��q��2J��� J�C�rY������cI9�@�H
��D5 ���L�7;E��
���=�DT�\�S�Q �6��j����\:�,3���luOiꀀ�K׭�p��O�"]���L��sȐB��G�! U�`��_F�	�G��e4b&��������
 +�����`$�1�~i��	�/����-��2J`y�"���"�Mʒ�(����y�,���2E��:���t)�7?HK�s���Uȓ�%����H�!��E�ƺ'@9����Z��O�0���8{��^ūH+ܿ��2MV��(H.hɘ��Y��P8�w��{%���� $�3��͇�8L�S�fo7��.�v�����3��}e"�0��T������p�}��a�H���������ͫW����N!u� u�9��-��[��p|o?L�pxt/$Ͻ���V("�V�آ}�@Y��r�j��g
��/�� r����1��#G��a/��{{�ׯ/���o^
@Ttq���F(v�b1��WH����,&#e����"}+���N�9��|9�8c�q������p�������K��x8[��OH\F�l8�|�麐���~2 �\�/4"��x �^g���]onI��`gO:�x��z�:t��P�l	���X{g˞"��!b�[�ag� ��j�!?�����\^�̕��!s���J�M�S�w�z�������A8�x��ӷ���y�y��SM�Zs�����Y[���^�g?�%܌zQ���s�)�XWV�̦��7D4ɓS�~�,��* q�?9��ܓ�H�'���v����<�>|:=�Z�޷#P�h���@pW�1�e}���ݻ�����~�Q��5��6�V}�?l��V��W��3����2������ay�	4eKN��O��e³ΒɅ���>�c7||�!l�ϳ�O!��d�Ml� LCx!���ْl#��Γe��L�g����mk��b^.E 1�w��乂�m���l���?��>��2{�������*z�خ�8�y\E�j�:q����g�i���g�d+� �:��uxw?�Z=h�Ȇ�~-�;H�;V��`���b�p�Z��y������������H�1�>�D����/F�:�=���]��ز��ի_�y�ߑ�X��c�H;1�  jV�V{7�����ۻ;���~a�-�t��!�[�R�Z���(���!��zD�ӂ"�NA�[m�x�Dc!�e�����R)B�Ք��[�,��ҳ�D~,��f>��H���|��$)���M�������+Γ��M�	�������ư~Ҿ��W�{X."RP�4�W�^���9�/��;�};Y_�,�5w�$F^�Y���;�K&q����x"�o߄�/���h`��+�k7^G
�ɓ/CÞC��)�3i)-+��,������(-��'~߉ޟ�˵_���<��^������PhG��:�!����ZY��Da̟�胔�l��G�>3<_HjR$E|����,W���H�4�g,��'@X�*u���y�/U�*�sl���jqd�SyY�Z�ԳBE�ȇ"�5g�{��E M)�F��E'�ݳd���)��)���V6Ȧlʦlʦ���f��G]���:ڕ�"��u:��
n���{��*�ЪH/@�I?zC;R'a��h�_z�DKC�ܜ�q*r3R"u'v}���}��8�2���/��$3&���P�	� �l�u� \��Q(�(Bex���/�;;8��\����tVM���F�9􇊎���4A�����[R8H}A<<��{j[��<b{��)߿���!�e�N<Tۣ�.	,�=ь2�°?p����ba��#Sy<L�QzQ�Z}��rK��r_~�/�'�a��9��t#��Ѽ��w r_h�_\\�][�;͘�c�	�S��}*@L��vH_I�A�rg&�!�@wc<_�2;8ϑ��	Գ�l'4��ރ,�d�EL'd��h��4U�"A�7�wa.`)b�(}t�� ! 5�kS&uXΤ-_����P�dC%0V��!Ofjh��ܰ6����`YĐ���d0�,>,�J���Ѹ�iﺙ��~3n�N��2eHR%�!){6D �IN�d�^�	���Wk�<sY0� (��Hm���r�#�k��m��`�\�LZ���]o��n���u�+�H��Q+�L�1c�0<" /��e���p<q�(H�z�H���ͣP�Ƞ��ݑV��VK��;��"ٍ�"mW���&���Q�}Pg���zE�Q���,��	�-2�h��纼$"�O�\*غ��6k��`(o���]��%�]�1ش��6�u���ŧ��UV�ȼ��9�{��T��-�ס�D�f3�{�5iV�0�B�ޅ�����	�v�m�����[mICq/̧�2 �z!#WIn�k�B1���)
�Q����Ξ2v��ڔ��EuA� i@2��Ͱc�����s'�K��]��9h}�-�}���DfD���Ç�6�x�A�n���t^(Z��@��1�w��ϑ�2�VE� �yNNqlV��^�{m�\�c�i�}�4�4N�"[�Zj��U�˒uÓ��#��m,��p��$�:z*�����9y�2������%�#���}|���ݖ2��'�=�?���Q�������;��f��w`�~"�j|K�ckK�*��+c�^����l�4%ǳk�4���[Ҥ��k9�l8O"��ѵ��l��ڞ��[O�Ī7*a4�+0 Pte�i8�(#t=�X+ho�kg��0����׹ؘ�+�9;�c�^u9�=������n+�?��`c�ӻ��̙kZ�Jv���LY��[��^��Tj-���=��i���[eű߶0x'��t�d����� S�V|IH)[6�oD�ؿNd���﹠�"s�@W���R}a&�'7x/�������������1�l����B���%e��9M��k�.D�f���0�m�f
D�(�m�z�?���_��D�)�b%B�GR �p̳>��~G�D��}7Y��.WI��g.f�%7��9%Bq��������und�>���O�nI�dX0`_���D"P�HDd�5�)z�Q��
�[�����B)f>���<�y�7�?�|QvP�&xs�	�,f�f�gW��GH���#�,�,�L���IT,dيoσ�l�s^����=����B����b�Y� B�&]��/�D&��Yi�\�lYȴ�yY��$_��׽���3wWe{���g�N������Ȥ|����K$/�?_W��V�Y!?&۰!��)��)eC�lʦlʦl��\�=��k:O%�"I$;�!� O��`�  V�¿�A�$��pvz�.�� Vh���COr6C;��dP����k^\]�n�+9#J�ÜG�f�#��냓��)�M�r��@�ģ=9\�QU��U���v�$�U�W�����*<��Y����4�eB$�j���O!�݀9Hw���I�|6��0�Pd� <�	�y�snr=w	��7�|~����t�w�7�~G��I�37%j��ڙ���}���yj�c��	�(D�F�l�e�� ����ۗ?ё+d� P���r�@�����y}�b����HDbW�ɌE��=��|E1i�z�|�t�2G�n��~�5�B�?����ԕ��rIz��G�7Z��*@���O��+��tNJq�t82e� 
\]�ީ�#��D����a��a��G*��sev�" b�P����D�R�Pjk��P@On��L�R���� �R���t����xX.�`Q>o~+{�GkR�������e`^+�����x 	9w I�r�c$��I�im�T�ȩ�6\�<Q��YC���hO�gh�$�.J�~��k�B�Q�y�O�Za�˰��C��^��!�����9�n�R逖��%�}/bM��P���h�,�P��D��*�y�A7x��3c��f�NU�$�
.(�|n"��^73�?�[k\����H�.ܛ�2 ���~�䒔Yj�?urs%��U�PO���Ks��<��3Z-�I��� ��9h?�5/��F���L�;Լfn�8�(�x���V�K9�v��M}ڗ�>P1���5e��`��6D����"<�"��Q�A�	 �-9�+�cH��g���W���t<t3��g��X��F �	@uѥ���G�/��q�	�ƞ���ek Q�<D�W+�ꃈ��\�G�3f�K�:b��oE�2�E��{�(�:���ߏ�����'R|��SFE�&PQ�C��Z�2(����+'A�Sd�D5j��e__��3���W�Jj����Q�<�����M��W��	W�Χ $T�DY�tͪ�������3f3��6k��*
 A�'S��o�9�狛	�ճ,,>Z���"�S�~�� ��9��pM��OȻڑ��g��ּ6uS�,�/h�ch	0�؋1�<��i�Q娈/� 耔!�#U��.��\$�ܦB(I�~��ȷ����Fb�S�d�>*FX#�f�#��(�`U��u��u�~����O��*�~a> �c�׮��"RuT̈�.�^�*��������J�^W��#s�r@ޕÝ�H�^BR�U%�9�U�Li��}7�}/���6$^��Ĭ�������v�X=�5J�A9�5	�	��@,�&"���s�x�����*Bg1Zq��ً߁IXF� �2�7��ec���s���1\�eow"��K�9����B�ya�1Խ%t����7pA!	�B���[b��>�Q��U�h ����rj�C�;�c(nq�~K@Zވ���a|��z�qo��6{+�â�̾ʾ����,���caC��C����k���m����n�^�w/����_��yM�:����a!�p�� �r:j�";����Ԋ�壕��o��/���������>���ޓ���T�9�ym@՗2���BG�U��w)UG�t�k]�ڏ�uH׺ֵ�u����@�_�����52A���[�D	�x nǇ+*�w K �R����ry=%03��Շ�HN���Z߇�]T��}W��1pv6���^?6��#�R���Oh�E��'Ѕ
�U?�D~�R�z���<lρ�fed�ց'��\��ӗ����|������᱌�`T��5}���*�Pm_�o���� �P |]�7�n'��
���:�>��>��c�b��^������傖`_�-���߱"7�� �Ba�Jn*>��V> �P�:E	¿#Z����;����O���g�>@H��f6��s2< �R�ih�^�"��j��V�lYeR��a���C4�;P�p S{�oCB�{~� 4#��ۗT�5����'�Ji�џ��*� , H�v�!A&AY5>�h���(����)#V��
B�EI�(0���]U ��5-����Z)�$/7��1����+0��0 �I�ƀ0�Z 2 �!?U�P��\�7��q� Q0� -p=���̯	&���A< Ģw�����7a��୏��?�����T;��������g�fa�W:G�c]g�Ϫ��zI�8�m�b���J@|Qf=OI{�H����N��M��I,7�����碯��C�nFp	$3�2{1T	�+1��{ؘ �}˽�{�B�2���o�� }��9�jT=_Sq����~�e�R������4�	$�b���)\�5CG���2��\�eUΚH޲j��I|���l�E�=>�[7r�}5[.����q��#�D��0�$'�CUZ�=�,NO��|9%!ҳ"�� 0=F����L���w�X�.����RVيk�7}V��V���G�6�$L=�����dCV��� h���4h}@���H�©�V����\ߚR����럄lu�C������Sv����é�˹Y7�Frbn�Y��oؿъз�*��a���r�qy�U ��
�td�m��w`:	m�1���
Ǡ݆�իB�c@�`="��H�|��չ�\�B��c��M�{!�U�Tҕ̇A��R�{�n���S'��b�58��9Hb�L��<�� �`5P�b��7E�s����(�k������b��@�J�,ac�\���1KUr]_��ř\__��Z��`R���G!�A�����O/9��b�r,j��e�>܏��sA����$�p:���XT�U���Fm8a���k�%��W���%��OJH�蔤5s�Ȕ� ����S��Gm��0������ߓ�p6X$�!�]�@%�̪���q�sص?�o��"f-D� /�S��{�~p]���9 �ɔ����N\�IM�'���jHRA-�맩fq�G�ók���5	��SYĸ^��m[{.��xΥS���X� ���<�!�� �7�kT&v?RH�g�~;�<ܯ`�#=���Z:>$�h���JZ�>[ڂڪ齑�,��}�8K�g�V�V��x���bޛ�.:�9�'fW�?à}_M3"4Җ*���Mz���S�y$&�^9�B������1���U�N(F�:��c2j�{*�]m�(>���x�0�ڧ:��������g����z��[����y)����������#螨{��jy���������@�.]�Z׺ֵ��#@�ֵ�u�k?��w���o�B��ۊ����@/�ۀRXQ-�]�˗��o^��g8��� -�F ��L��X-W��*K���3��[�ra^�x*>P�����@�`T^�=>H���:x`�,���,��U���p��?�/����^_�óYm����W������ގ��P�ј a���B>��rH@7��@-/�ԓ��!�|�^]���	
���O�O&�%O����țW���L�.����pGFzLxX�8��e����J>7�e��d3_�Wf�|�})���w�$�w �&������!�bQ/�03��q�|�JxT����9����K�ӕ�+ѷs}�d�ڪuX�������
Ğ#Z"�z�YV-�̊�w9�ר-`�b-d0�g�8�~�|+��~(=�0�a5n�q	|kX���~��:��h<=��m�z�y�+R#7�JgY�S}�svsB�V��KV�;P˸ڠ���4��P�ѾDYfo����V�k��f7s��(HH4�5m8���@Q�T�j�%�P�?���fm������W[��:��j���ܐX���6�5�'x@ҋ�-*�˵�>�/B���-	����B���W�����C�e:���6�#n.T��IX5��)62 � ��3U _ ���dȨ�$�U\��o�3AQ�;$s���l�#؅�r �Qf��A.W"ƾ����z�T��:�h�gVkF��Z��Z���`�k>߮��15A����}��Q�����A�Q]�sk`��;�O�4C��`�^+9	����rh��ST���8����j�1 Me�g���_��4 �E?g%y�9���0� �_�����h����y۷��K�����X,V��}�/��Y\�
$�* ������4ȱ!���
r���I��^�#р�
0�+�A�h�j�o��-��^s
I�Si!��<3Yȁ)���狵l�z�xmI{:'6%�J�{�ϻ�<����VQ��7~f@|c ��U(*�e��s�'�ݵ��(���;KBd
�z^?���B����P9;&�:�`Ňq.0^�oT�u����}�K�:}% ��OF V�̄x�ojI�C���'�������|�>Z` /	 �^�@�\h�<���HHi��H�K X��pB�e����R�4�/�
;�.��Ei9S�:��4-ɿZ�z���템���-!��t3�Rv^����e�Ed*�v�O�o!m��b�be�8��wj��/E�Ѫ>��ƇT[�V����Ғ ��q	EX�3�ֿ�.!�!��B�ds�����>�^�y��� wC�M��߻U.��J)��+5��:_9���~��F5�
��Y��)<B�=,0�0��2˶��Pp�uY)�u� ��p�H��X4��f�{�� 6[=���Is�:�{��TFْ��J��Ĵ:8{�b��TM:o� �,��Ԇ΀�uu��v�IS��s2�.X�q�*o豀ɬ6=*07�*{�����
�������{��}YA��uh��xF��R�:��c�m�1oN�����9U|?
�����f�е�3��~C%6�`��D�c���$ŭ�%8a��Dҵ�u�k]�w�:�k]�Z׺��i��.�w�VTX h10@ŧ�CHOvf��Y%YF ���Rޞ���ޮ��a{�p@dw7���C�]ʰ�3�������b��̴g@?[����Cv¦(io���US�]Ea�
��x�cգen�����=	<��3non����rvzJ ��9����Qq�ǯ���xM;�)�ю���iC59��@����p 2C���W5�GB��������G{����K���1Ht�fǒlR�%=���_��g�����#�W2�-i] ����GU:�W�ȯ��!�% ���v��ɀ������S�r�w ��У2�"`�	������lZz��0��dGV�Z��oy �,�"�Ct��чuT���I�z��]=�k�4����/@k����"�V�:�p/(�'x3[�һ�sT�j_l���2>��s'lE�����<_���T���hp��*V��q��Q^Au@-m�$�m9*����1p���
8���*���,H�cŮ�]h)QJԘ� C�o �x/r**�>�@"��[߻�̺�!����ґ0[R�DP-7W7���kV�N�C�X;t���%^i��
��`*��G$`�39!� d� +�4��/um��)��c�C��`=�r*�@`��h����A��.�Q�:�%b�	��1���(	��4�x+�1T'Y�b�cE�� ��;�ϣZE`��1A��;�i�+��=Z�DV	��t��j��*�f+N�Ӑ8� ,�9+�}*����ҥ��H\�p�be����#@��7-�g����!T
������k�4��lVc���ry�����+
i	�q�ʍν�{$��$���\4�@���Z��t�wM��r����d%�%�6�wI���0N���9��$T�����
G��ƴfA�%������؈�B���4���Y�](l�UH'�����c�� 	����B?f�h�����0�dI��rM�8�j�_1�pM�s�?�:��X%z�\�.��.�mߩ�zF@�Ӱo$q
��*%0�@��>� lB��[���d���=VWSD�A^���⇡�Uc�^z|��k*=@�V�+��[�� +�f� ��L�,�����F<��;0��^bL�Y�q�shTt�Y������ǒ(ٸ(�.Nv�T��**1� �@�.3^�I�)W�m�Hu^�G�ol�u5ӿ�$��c�Ӿ�h-���Y��!�Uל�~k'q��*��������9B�j�ܽ66ekڵ��]�G����寧�����'쐐��y�,5�+|g��v�Đk�xt/l?�j��@eՄR���,���ɮ�ۏͮ��X߅���ف�2��%��6ۮ+!����Y+nCă�߇�iY��$�;Խ�@,���VY�$�MA�}�*�VA�Uv�[�9�3�?�\cE�]�~��M��'�|@jxN�edTC�;�W�NR�"���
'� =�]Z���v�q���QLa
+.�������{C��Uf|?����@�����9�;URs���LIR������Ž�4T�����;�ÃY�6�q��<[1[Q�?��}�_�B��J?������Z׺ֵ���oҵ�u�k]�A����>��A� �^/��؂�j��@�&G��{�0 U�Ւ���>�Ao���g��rus%�U�@�Ýc��;�-N� 퇑l`��V���b���ުXaó�,��V2�Z�^-Q1�Ї����4�j��x3�,#@��K�~ ���l9�ޞ���d�{�䃟�/�� ����%[���}��B6�r}}ðƟ��g���?����������#Kg��� �-�P�g�`�#E���@Vʭ��������ӧ���2�}rx����|���#��W�A�{�}�����o�����C>��3Vz�h�&^D���}�h��{��M&螡�YI�e�1c�nT���vU]m�'j�ͦ���:�e�0���fή�r{=��|E0�u��m� ���T�~ƚ���W�	,(I�R�lz�D�����@�y�`�O�_o+>�P+V%�u.V ��T�FF�'y�(�:�de!�id����U��U���`��ֳ�QI�VY�q;P��\Z,���u�X�y�Ԕ�Ψ���~��|�柑�GH0��-����fjam t�2��H|D8�w%A�s>1?t��M��q��p2r �3V�0G�hU�Z([���u�g
TE ��tM��c��|O�I�����x�	�| ��8�Vߣ?�I�/�e�O��Y�S�j�TT%��u���\J��`(y���� 6��	�E�B yA� 0Ñ"���G�q�PQ8hq��J��2EL���C����eo�����4@��L)6�s���,=�ϕ6`��C�� �������b�
�ʄ�2���\�o<d��\�� �a������(�" Bl�k�7u�J_ _)m�1RU����B58�}=z�gT!@e�db�j6~1̬��E(��[?�����W�9��g�;V�3M�ۓ�9"�hc���P�����D�o���vil���O{�^=V�/�kq�<	�lM���G(\�$X�h��@�U�YT ׍)�`m��Z�\x�-neg��	�� _�s���@���e
�.�ì��>  ��F$�˝�9K2���p��q�ם���PE7!�~�{uJ�
c�$=�8�f����T���~m�: ���ņ���R ���
N��s������|p����>@:K*kZ��Z�+Iʔ�H#M+*�L	��p�#a
5$������EE��Q��2P=I��m�EF$�^ɾ RRuY��Y��T�l�����*Hplz�5�ڏi[$Qq���ա⃲j8�[�*��Wz��u�K�H�ؔ�AE5&� �S��!��}�Ec�`�-��=w��Ya�q��xmm���v�@�$�i�W�:��6$ N3��.D��c�4��8@~a/����h �DH��w�~M�KG7 ﮣ�/���/u���k��X8a�\��en����5,<��h,���P�V�]���ڇ(��=A{��?�fE���ξ��_ �{:Wp^���d̀�i)m�`�l�T�=��ܬ
^;����_ ���r�o�P|W�����.���u��A��R+���R��s�[�?�>8� �6�$��fu�זo��ڈڅ�b�{������e��.�V�pA��g����X(U�^��c.]�3����vo��vn��b�����j gB��C�g��;r��5�iP�%�T6�\�/�dq����K���n��7���p)]�Z׺ֵE���u�k]������`�Aԗ�hB���0H�
�e�+b���L����cfe�AOnn�X�d1[��y2ڑ�`@���vF s�h�q��PƓ��!+J���������C33�q���\�_��$*M3�JG�'��ąAӮ�EY;�ʗA {����#V��n�����L��
P��삶5���O�������?��>���?��|��7rqq*�(�'~�J�|�B���ޮ�W �"��l.o���=�899���>�j�gϟ��<�gϞ�?�D;G@I$_/���+9=9��z����x о ��U�Ɉ�� ]ѷ��b����܆dBQPY�j�P�������ܒ����pL �=��걟�L��:���g� ��V���鉗p�B�NE@	{�������<{�9�sT(0(� N�B� �Y�d�S�{�QE������5�R��D�.@�4��|ѵO �W:�#?�~Z�*+�-D�X�s�'pjꌀ��=�+Wa�di����ހ��$�yQ��w�?�u��*�K��tG�V4���I�¾I�y�ڵ�jX �������� �z�	��U7��=�Q[��&PI[T肸(Y�n[��|ZM��e�4�dgkc!�6�v\�.�{�|�񚒂�xXmm8ܴ�X�ږU���o��h���b�-�VE��a�y�lCX��m� ;��x�Y�'[{0Zh�V��=��|�rGʌ�
����ֿ���L:.�V{8�*q[�*Bj#�/bA+���c�q "p�(_�Ee�U����۬-�b[	M����u���~o���.E*�`%��X�[� ���-t��qk����j�:��S����@g��� ��[D�|���sAʀ@ah�gs���m�c���VUL<Ϸ�&@�PB0�y��6��*0j�����@DP�]{U-$�j�_0Ka`���7n��_�dfU�����J@MҪ|�@��U�T��Ű6�IP�{�1K5��z���[7-8���\lt^X�wQh��$f��O�50�i�JhJM(�P�OEde �X�UA5Z.U`�J̻�����/�Ndn%�SY.CD��Ƒ��_oH�a�7�" �����4��h^��j��1��nn2	VK����G�5uyT��ҡNJ�����t�#�{k-��Z��l��ڢg��Wn��	8ú�a��gE�\�]�R�a�} �������c��;���qת?�˽���-g`� xԌ���-׃�a��m�v�4�*�~�C�B�Q��'�]b�X������	�y�/}Mڳ�k�����c4���ޑ^_�����E΋S�XNG�lA�z�>T�k�\΄Gb�8��h�9A�p6��^�����b�Dz^(@��c��$�艹�i\@�ﮋM����nY ̋�@���qs�w�n���l-=/rs���$�)1b���J��*�J�a,����`x�� �Z9?1�
tXLA���~@�A=#�;��E)8~\�Bw�p�|���;�?�M�~�������l���NW�h5���Z̦������*�%�j�Z�z�]�핼���tҩ?�ֵ�u���:�k]�Z׺��i|����3���BߧW���QŇW<(dFp��=�K>��O��e1��u�\���Bz�;X`���z&��VH� ��H�v����!���%r���d̨H���aOq��5AH<�LjգV]���)��a��e(g�z�m�7�& �I/������8���Y�y�� ?;#�-��~"��\>x��r|���sA��dg$���H" p�77첾��;*^݇f3�C��@�����rs;��h$�QOd��#��P�>2��e!|�����~�;�~���R�� �ҡ�1�"~tt�����x Q����0p����A��pon2��0fU�=&���\�xf��Ymi`�f�5�� �%���'�_����� ����C�G���\���X	��7�웪E��>��0�|w�+�q_��R�౎Fc}����l����K}0�`��`�
u�no�I�=z�� ���F..O���ss�`�V>P��������9�C7:Ψp9GK���5��N�d�@����mY弥eIe���s�ֹ;��ؠ�c�-�@��S0h�a�n��V[Z3-=|����rVMj��#?X]�2:uJ;�������TS9r�ę��n Hk���r�%|�S��U��}���m��&���iSxOF����=���2 ����9�8bf��D_H����� '�|XM0�7Л�6/2�5�����j���^��%i6�:ʅ�"7���=G�6���3fnh���@d�i���o���4V��"����H`u���6�������ʔ>g`Mk�6�$ H����́�|���/�za�B��L�ֆ��u�9��%��!ZU2�@(�`�5�淚�x[K��%���fo&�S���uh�G��ZC�ܑzt�㖳��ߑTq}�U�4����#���ȁ�ei��ez�9歅\�m�5u����W�ۏ런J���ȣ=U���*��$�0gh�e���-��$���������f�y�s�-���q��U�6�����R�՘	�c���-lxln\5ƻ%_pL ���㵡��`������L��]X6m	��2�!�߻2�.á ��f a�M���s�k����n�ll	˶�i'WJ����YY��@��m�ڹR߳r�\�\����@9rɷ��b��ƀp�������G~����H��9�c�k1"��:�A2^:KP�e�C�!��q4���*����΂E(8���TcҒo�4��xW��~m��<�������#��Ïegg��D�-D}��p]����	������gav�	�|f��)L-"���j�Xc�=׷W�b����G����5I{(#�B�1��y�����������ڽn�?:�#h+=�d ��%���{߹��6�#>Z^��f��o(z��r�K�� Ɵs�m��i�%���́kkj䳗P¬�����ΓE�~U��E���}��Y9U·��zo�����ȯK�C�����L��������k]�Z׺��iҵ�u�k]��oyd��o�x�J���uU5ۇ����
��WW�t�� 0@��&�|��W�O�����+� !� w�\P� b��a���ӧO�{#oPz�՘�N@E{�/��y�__L	Ld�A����b>�������]���V��Mi��X D[ ������{�s|x$��D�vY���8;?���W_}%_|�/A?��?ɾ��+= �8'�3�W�r;���|#yV�*�x�>��z���S�k�����	��d��иmxtXɰ?���!���t@��b�Y�$�st�@>���������zl���?���%�. У����W0'���o��H�����nAՍ�`{�XXNv�v�cr=���lT�W���@L�� �P��	^�o@�ʼ2�, �	�?$����d.@i4�xnWW�ryu���z�9 �0�x؇eF4�w �A$ �� ɖ:N��t|tD�avs+��o���y�S?��R�`�@��;~vqN8 �{�;$@~}�����vJ�{˴� �Xn�fm@�f��~X���	���t	Я�1�d �"���AXD��ߙlՃX��r# ���� ���n� �����HȀ�@��B��������|g�N/5���rx�gĴ�I*�oT���0�i�$��D�X�H�B)�Ͻ��,�bd���G?�:b��2V��c�>�`������~j�a���P*Yƭ�`0��>ا���l^�n����Gų�>��$$�:��6s��ȫmAq�.\��#)ٮW�>$�*[�s�2�ue��=��O�&a\[?r��2�������t�p�־}�?�=[4[�wf�QK�!����S���-�ֶ���ۊ}�>��/0���T�s��ẹ>�q#�P�����Ibk+��-ad�ԐD�R��jhTУ����g!�q���X������,j<�1����R�{�g���+j��04X��e��0�Z߁�E+4��چo(3Y�����S����ȁ�-9��ґz�lB�1���H~�ȥ��@��֮g�*1r�l�x�P��)��Y�{p�m��-������
$,��Fǻr$.*�nX,��/e�4���*yO�z��#~�O��yd�+��F��3��U�7���z�{�x���msk���P��x��7�#�N,�]M�/Zu�G��Ue�E��`��}s0�m����S6��^�P�odm�����.��k$2��cF��p�C6�9�f��Y�h��T��������t.7z���ɃX��=��o��R��G}���.��6���ڤ�{+�����}���PY4:�n������O�q��0�[�~Zazf�5��չxP�%��쌷�8��
ޛ�
S
:R��#�
��NS�_iIx. �s:f����5��@�£6����ۙYCq��Sc��Y�f������Yj�;7U�]�g��$	��AOC��N_'M�և�o����Q4�S�ݝn�l�����Ɏ?o�zP��"6���UЦ�d��2U�|I��׿^5��t���[�߹t�k]�Z�~T�#@�ֵ�u�k?���N< ��X-�V��C��E��z����#������k��.��3��|��ٙ0�ᡄ Z�'?6�ý=��Oߗ�H�z��a쨴�EB��b�$�	���l��=�5��YR��,�%LSg�bA��,{Z1|�=�CA����SLx0��:�y�!|n�Oew2�|�����Z�H$�~�������O!�˛7������ݝ�Ϧ$jVP��Z0���@���O:��R��Ut��J�v!����w/�~'�WF�]��=98:$�p�wޓ����|��G/w&#��?����`<��Ϟ92��V�F��pǮ��+�D���,�9		������������^�a��A�I{v��^�-r�J�4!�9��j �:�&1p}eNo��<Z�w3�{8������<�ql����{;��������Ĝ�}[� \���	�@�̓��`�~=�?`������#~l�vuNL��rla%3�	B��yz}Cu����l!��pZW�JD��I���1|�SZePG�-�� =}��������x.W���$D"�e���-dM�����1	T
���>�V�P1����YBu ����qn�hR�0��2p�[�<�+tL��7{�R�|�?u���Ŭ����7�2,����m lT��F\�y\��4�K�ԱÄ��3Z�`��j��*q1 �1H%LejOڠy
PG��{
-���a�V�l ���<D({�,΢�q�x���sj�"!Pn��VY���&{�뺗T��.�Ă�Xw��0��dd��gU��v��n[�l� ^0�3�T�^� 4=>{I��PD���Q,��kϩ���*�AuR���A=Ae�. ��rA�5p��>K;X@5�U��	��w6Y��\H�lt݅q!��)LMn�$j�m *�a�gؼ�#�L��3[M[:�̈����Z��� z	#�U_����{X``�i��0� O�c��	�c/����+i-����Ǚ�� L�H����$�V�\/Q��5Qֲ������I��y ����56iv���/luB�ܸ��f���c�_1&�fz���y�:�-���n�̮����$�>�O�I�9�r�P`G>�%�y�n�G�S�q\�2�\]t���~_� &-�nL���;}��mT�+΁Щ��-�a6?�^�V��� �u�1��̴�#��,����Z[4���A���6��T��ܱc�|�ݟ���8@�����у��N���!�/<��22�IԂ״�x]iB"A��؏�y�9�������`�Ǭ��3�l0kguV�,(�\犲���W�ۿ���E�͓Ʃ�f<���J��gOSڒ��U���j�b�q�Wx�a��gd'��Q	[��q�4#��Z��N�~�?z}i@�h�z���o,��H��.V���8#E�o��⑸��*7�)q}Jl�7�e�೽��q�T�\w��e[��k�d��'�|���(j���Z�c���r��]`c�`�G�W��,��xV��ӛ7'�����ҵ�u�k]�Q�� �Z׺ֵ��`���o���1�Wi�B����VA�J�d� ޶z�_,�rk�y�`RkW�-��޸J�Z�ݑ<}�T�=���y���`Z�$��fMp >ꏏ���?})Q��������X�1
l\Ap��� ?6�h�E����r}}%o޼���>�L@�#�&�13x3���|)�^+W�W�<}������Wrzz"���T#���F]^-2K  � ���U�0�k���l�kS�W�~ޥ���P��������3�g�R����������DU&@���KVm�;�x���*�À�.��F�G��
$ :��]-��f�;�U� �2���
qv*BPS8�k}����`U��v�-�
���DYlm��C�\52Ô(8� � ܅�V\m+��1ߐ��?1� ���$�U����1���0I�O8��	*��X2�z�`�pd�)�XA;��&@�0�8����O�S����+��x{&Yc� -��m*q5�x�k���L�΍!TTl��o�.�6�w 2÷�XT�0i�|��a��*G ����3K����#=��mM6ϡ�T0+*7=悘���Y� 	� ���g²�s���öz��ʁ���B�kAJ�#�\^�� ����x�YF���$45	�N�=��Y��BWN�P)�{�jy7�F	}����i�*V�̍(
$R3s�)TR�y �(��eZM1k��S6e�j�$�'Eq*�������	T�D��	��1���A8a�#��d�tƹ��8���y'�7xnz\ kʸ���oh�9�#��i�$T?�CKҞ��c����7���Z�69����kf8��1e R�����Y��vC�1`�NeO�]Gu^3\��ufQ��	������H�7hbG�6T�$��f�j����tK(�tm#��z6%��*�lND[�7��Ъ��F`�V��ǲK���ZK�Xߙ�j��z����/�����dG�$2}�r�\�5�S�0c��N##�������@Q��,(�tA���FV��zg�߯���w����Vk��9��T�.G��\���ù�&S�e������\�Z�)(0���>�����w�p��Pu�9UT�By�]��C�6���Z:�Rz$�t:kߛj�!��*�>�"���}�)u�m�~v����$��cO+��]���Zu�6���ܟf�u�
�2�������>�>��{�ʇ~H�c�Dz���s�T�����,"GT�q>��Jno�6[KH�[wd�r�-��pB% �o��r(d��ߣj��nZ4b�"#&<BQ��1��T� �I*�Њ�'����n�d��!�,�PL�q@��N����N̈́�1�▝��о����PP໷dF۾O~X���ѣ�H$.@�gڧ9h>�[z\����������("�� i��)�xW���,��E+8*C{���$0OA��lI|�c�Z��==����1��i�e������Z�=]Ͻ��h+i�(<'�O�,hq/AU)�������K����l<���n���_�x���u�k]�ڏ�uH׺ֵ�u���@��y�33@��w�㙤&�P�` i袚k��d1_郭O��Z�r���	@#fn�� ��T�3�0�����/���"��#)%���"���~׌U��{tP5�Z��#�'�6�1�}fL�i��lz>3���|�~��,��|�oof$p 'P�xpt���͜`�f�����͟?�O��o��`G^��V���K��������?x< $Pa?�p<Ga�ۑLF}M��*h�Z�d����	��4��d����C�G -ܾ3�3�^�2���R����F�������OM�%p�EYo�A����<ǈʕ P��*�< �~~~!��T �6M�-�RG�&m�6Nr�|�Q9\;[���ߖU������)�V6���rr6����3t��ua�+j ����?}N��e����<��]��G����)���N(1�k�$W��{�;����䡎��'O��g�|űc�Pt�eS��@V���6 ���%�:���T�v�缾���=�� Yn�5�Yc��V��܆#
�}WM��|P���-�♭�fe�5 �Ɠ��Χ��^�M�U�z�6>�|�a.��9�s�\e9��a�eA�ȁ?ᘡ��ܙ-L�s�0��'qB�ەF1������Խa�`x|���ȑ �q��F�]u���9���Q���y+Ͷ�ߵ !c�
�B�S����=��Y�ߐ�3e��1@N�Y�ǐ������^�$P[����<c@we��-P��[񷄞��"����X.״�K�ʀ�Qa� �̽��9��?�^?�dpG`p����z��ǚمl���f%#�P����-��s�E����� � �\�xl��9�xm�:e�r���T,���@�CY�ż��Bs$J|����X�/YH���}q���`�@i���@�Ү/���!# bFծ��D�.ϙ� ۮ�͗#M[�Ap�rKĭ����> ��j�S[n�6����2Y# ��^Db��1w�ȴs�����˰nb�fa��#ZQݢ�!q�3Ȩ��'��΃��,������g�q?]������¾�Kz�<&	��d����) �I�7w�>x��w��yl �0p�jͨ�\i��$��<��Z�z��" E\�m�[W�O��������4��:)J���4E�]'�%_��&sw�����MA�*b�z��z0�����o⮻��U�7��q]�M�A~<� L�y�����W�����{�yXG��bqEK䗓�����"U� -�-�h*=���Ef]i�9+0�`~�bl�����B�I�6w� I ���޲^lx=�lSrT���8ǼO{��4ec֋�*$Vq}F��0�u,*��8��,-/%	��Z�JQ��0�qf�F`*>�Y@��J�K�>w�cK2ؿmŏ��R�f���?�S���jCb������H<����r�|�ce��9��g$�o�Hf�e�{��m�<A��Ɯ��*\{�$,�e���]tSw-4�^g�'��-�a���߿�Ov �L��K�Z<(���n/���O#���P��u����W�����v�_�����t�k]�Z�~T�#@�ֵ�u�k?�����Rn"y#G����*HX]����)�q"fw�2�>|�f-�J�`˄g��bnv��(sW �G�������P5���O�=�v HC}^�Z�[y�����}�ᨒ�gAm�d 2��PPT�o���6�Xy_Y�*i�P@�����d4����8���=W�v�s T?}�=�䓏d�3fn�o��z>����[���!{雊D�4�rx�'�р ���+6��TV��,Ws�ջ�G�c4������z %H�k����ՐD *f��Lo��/���XU�Ym��=�f 6�C�J�ƀWV1#��6�u4�:�*LXS �B�����\Ǻ�ѳ�,,L�a�^��3W[ޫ��&�Z�wAÉ)��g�[�<�fy�\�e��S� 
}�)�&�*˾�[��r��.�jX\��Ĩ	 ��	mg �U%���� �X������ �8�zSJ7 $����]�2R g�������j�U��b�я�q� > ��PJQ�?Ko�fU4�RYu���<*��A��C�j�����X�+n�����fZ��2_.�O��$Ea�T7��U������[�jH �Py��в����X����G��.�������=Ps�y�8�����K�F�z�O�T !��Z�/ F�I�R�'c���3�)�Y�����ކ>37(�%��g�a�O���K�I9�I���� p��8IeO� =Tt��A�����5\��X�HcvLT)P�b�πb�d ]Y�[��y�Ç"o%�ο~���	���/��D��,̖��^���!�i^���U�~F?a.���!l���x-�HE��l,B�!N-�'�{FPT�]��o��V��ĩe~4>f���U�c_�-���}����7=o���W�d��ׯOG.��)C0WÄ�-TC�����l�B����}�����R4�6�����}@ -�z;�ߤ���k��$Y� ���ﶹl�p'z���w��^,7�7�qlD�e�D<�%��v�V�R?v�T�t,��
ū�k^�3}O��;�k����e/�+a[�}(+���a�KH���_��l���W���a>���t��-����^ m6�Z �"�2<��F$#cZd�}�ΐ0���) {Vz�1�#{�I��k�s�)f��>ļK���lʰ碯(� ,j�XO�V�bj3�F�����P����Д�b���S��Cw�U_0�����`P�[řІ�W��J>����:<�Zk�KP+nr�`r"��{-9�y�<� �9��	>ܩpM�fk+�l��utKh�]����E���fEU��H�V�����s���:�q�UiY,Xk3߄���3}������Pp�B2�L+�Wm)3�є[���v*�K�0&c(is����������Ox������6�q=�]�v�R��Ơ�n�.���ީ6�Z��$�!u��7T�䎀(������8��pDF�g`���	�c8���j�c+i���W4���v^Ȧ2m�S�T����w6WX`����Xg�+��;�ꠅ�_H��V�������������3���@d�$@l��M���z���������}��\�ֵ�u�k?�� ]�Z׺ֵD�*,}4�
��ٕ�r�̅�٧ ��G=�n��2���O���|�#��b��q��z>����pQRр������atz�F^�|I����B�I��q �I#g|н�-��]X>�8���fM{ Xw@��ワ~�K�v�pvO��D�}�? `�,�,d�S5+<V~�|�R.(y ���2d�/�y z��T��v�r�po���?}�G��0-������ ���������ʮ� G�,�3VN�b�po �<����!�X�O
V�Ӓ�1EM�"����}ːvXF�i��X
���� >PM��ʲ`u$���	���U���F����\�X�1���0�Ȋ��!+8�ܹ���M&g��V�gdGh�� nx\NMA?u��$ �����*YQ�T�/�s�ϖ��{�OY�.��0_����-yW�>�$8b@��=u�G �YTm8�q� �ִ 3�
�)���rʊ�22��	w ���� �ٲ�~ϬC [���M�u1	T���T0 N{=�'�_�x%e��w �~a��`$�y e�����(�o��`d��F��'�Nvtl��������2�5=��5TYK���s�?�u�p4��LC��o��䰣�M+3d�xŉ����J���Ik)��W��g���P��Y]�,�Y�/�Z�~4��HJ�s� ����G;��(��\_�̢�b���{x�/O�yW�ڟ�W$A����x�0G0���w���Ndg���n�2Ӿ���$�& ����v��%��$Z�t�x��-ԠZy�}}~~N�O��Z�c�eggryy-��'*�kG0׹����������KO?��~�UI�����G��X���Taݟ���`����#*�Bg�r���X�u?|x̱E����˅Lv��6�g�Śk@>;���G\8ߠB�c���5b�~fF����Oף���Pͽ��	����.������ثG���i�PvQ��൑�ثv���=&��� �}x��y뜄�\��3I��Ht{7��@���΂����Ys-a���}c�g=l}!��N��՗L���>S$�����3����{Y�� ���7Ȉ4-�'����Ρ�Ǖ�)�|�\t>�>�5���eW�׵#��O��R�I腦�S����ެm�
u!��S�X�'�W�cA|Q%�����c�`-!kb4���9�>X�S�C�o�iO�ٜD��l�8�Ps��R��P=},7z�u�ի7z>C���ΟH�
�ͺ ��d�cp��u E���٥���<{���Mt��l��.��.H�8����~g_��P�Ӓ�P�`��:.���*V��&P���������dwG�ӌV�s@�J���@����W$<@h1#����x�s���5���>�qO�=a��c�'�����7,���8>(��n�^�1Ǟu�x�6 ����f^���v�Zx��;UUkY�3|�D���]8�=�1{*S� ����ā�2���fɹ�υ"8��,���\�Y��+�v>}Ƴ_��ĵ��|��I���P��E��C_C味�d����P���Ox-x��|���E��O��5��@���ǀtk�[�5(���"@l6P��HXS"��{!�ƽea$^5��ѵ�;��/Z;޵�-6V���}�Y`5.,ݿ{L���,�
�i��^�

��ʙ��̒&���3[��
U��v��	ˠ��3�8a�RM���۾����k�r=�k�\��R޼�Z�[�K��՘�T���פ�>>~`�s]�Z׺ֵ]���u�k]�ڿy���l6����c�B8�}���o^��D�����G1+��ؓX�Ż{I�����T*}0G�s�Z:�ma :�3	��V�'�i���ýC����A��r!Y  ��Ë���<��PY9�g����J���j]�&̭�� ����a`3��\2���{^�V���2�Z�{]oU-ȟi�������˗:�/{=>X� @|�����>$�e@�zJ�U��=�q��~xx��J!�a�<@�f���WevF�nn+�Q�Y�Ax=�MA���l��c�t��PI��_���R�Q>���к��v��09=�>��f�*c7�-̺%JR˲�k��jG��-WI͐[��몲 PT�CS� 4��1�W�+�7��@9��q�P���2@\�� ��s �R=�s���-�	���଴P6l�L��)hU#���C@���6SC�6���������D�;���$��BdT��|�K @�'.}��7���Ս�����h���G�b�Q�0���<|�D�-~ @҄8Jk�B[� $�����tFPs�u�
��tN*��"7 D 2{���ͥ��-y��ў	ڏ �p� �@�E�z����0�;�j��ذ>�|s3��ψ���e����:�� �P+�YҬ�y��-A�$�ٯ��Y �N����?��很�n���9��[�A�oJ��I|�Sc�B������-e��wyyI�V4P� �j�6O�<�<ս����%[�:�W����Fes�H<HM=Ә�c��qX� �A.�ZVz�K]gf}(��L�1�]��A�_]���	10�P��e�LT6�9?w�� 'Ac���s�p�$��<&,X^�MuM�\6����5|�&����+AlPq R�� �H�9��V�'}=�Bb�/ �nnnIh��	=��Pʀ<A����ο[fN!0X\e�T�2�`b�l[�?�� �� m��Ͼ�{яP�T�F��h�� ��G��&{�:��T �~�F�������7oID��� ��L��I��^��͙S'����C�uY�}�]:������B�)H!�H={�H�9�{֥Y���ÚiZ��n��&�U�'�r��e��~�k2M���U�����_\2[��c��ѹ}qyž�Kg��L"��AO?{*]���$��ϫ���U���푌H˵��8K�B/�UI�c��J�d0��X-�M�k�8�!(�|$�����fku8�ѵ��{�����z����ށ�}��kz�l�vh�X�[P{��0�%�ù���D��V�w����!����;`ÐpX�E����?����s�%2� <R����W��	JM xu��5���(
��m!D][nF�����6S#��=�U9��a��h�u
`�Pc�3�A�<���]�3]�3�N��Z�5|�{�\�m���׺ք�G%��"��|�%k�u�SY�P1�]�Ȯ8��;;+k����m�w�]*g��{���mx�6�ĈZO������� �PZ8:>�����h��p�mk����?ۀ��垉D�`���2���5��~3�������,����DX�E_el�}�����k���X��ޒ �Q�ޯ/nd1;��ש���~�J^�O`ysاp����I{I�{�6z�k]�Z׺��jҵ�u�k]�7og�gr�A
 �P�F��O�M]����z��	@�^����>�T��/�ߓ����� iz��<��F��Ζ���� �	��wH`��������Y�3�`����'C����@0 �����8�Cv09G���U���QD��v+	,2�.��)�>���
���[�������q���V��
�p_�������훂��7�S<8" =�C��E\��5r�f�0�������U����=�&�6���8&�F��xXoV��E�)r���m�oo�ˊ���� 5��'� ��X��XXaۂ"�P���b�A�c�# y�urZo�~g$���ŵ|��W�E%����`nYesA@�x�{���D�@�y�J_���(�K>X����F[r����&�O�lɐ������~`.^�&}V�YI�V R�c���#��P
���> �\�C][@o�����$C�L�M����ߓ�ɞ�cTU�	��k\�+�EX�Qe�۹�pjA+gu�&�A{�.�<V�@.�Ψ�������%+t�ْ >;�%��e���\]�_�W##����A�$#��O�z.�#62���9@���
 U�:�+�07{�S��Ư^Ko8�/�=��s���*'8o�� "qL ���뛩�����}���G�!��KBL0� �ON�d��j�f�����1�(��u��!�1AF�{"=G}X��r@��}QJ�Wyܛ � A���:�ʀU�s3 w�ў,��7�@�M �!�J]���S���oI�� ^��S����:`.���խ�ۙ�}�y&WWS�� {��PO\V�=����*A������K̠n�9�C:v\#2p����MivOXST�x>m�vt\0���;%�ygN�G�%�z�aD�a<�_Ț(k��n��M��˿�8�t ��$�@V�z�����%��@������*Ҙs���~/�� p@��K�;p�����v�څ��Z���g/HH��}{ʵz�����r&���� �S4���f:������~���͛f)������vp�W A�S�ܼ�����u���}��w����
L���6���A���|�B�EK]?��V�j@��7��>�>h�)��w`́c�O^��*^Z»�-�u��F����ͩ��Z���#f���qUH��l�� �qN��:�$��6����F�?g������u�[�i��}@�uW�c��q�\����3�x���S��;ϟ1����1&d����,@�
a܃�@ָ�V�ֺ���������kڧ��t
��7��xwDU�)?K*BY!V�������nf������|����w�〾�� ���`�P���{ܓP��2z@�$'�9�9��^��J���}�$�G�������>�E(�lL{���F���~���l���(��ߕ!���sŢ�yl��-Wm׃�ꤕ=��+�`�Ā�Y�EK*�˝��#�z	�_[�����U�q��)-�ok9e
�V��گZ݈S�l������������@�Bʢ%h\	&���7�*c�Xd����1�/�VDK��ăe6�e}�"	b�ȼ6�K��Z��T`��Y�Ua]{7�ƞ���=���k��0O���Q���z�3�燪���Z׺ֵ���ZG�t�k]�Z�~P��h{�{��|�����]����bȠ��@�X��A�*��ن��Od�{��ڷ@TWi�9�� >Qԧ�	���L��{�{= ����������Ľ��UP1�֫�s^�����-�b*#X�V�;�1]��~�c�N�{�dЂ�N{2�/xaY 6��^7VQ]0,�=V���Ƭ�"� (L���W������n��],� |��'�K O�ހ+ UF���k����%����E�Ҳ@B����
W�-y@P����P�t�����ֳ1����'V�2�}<6k*}�_I�}�\f���NuE��\�,���h��@˙b������B7�Xo��8j	�^j�;�g ��=>����jRaU����6(����R9� ҄�[9UU%���s��kr�wbYV����ڛOo���T6ӛk	����O$�����F:���6S���r�lHRK�}�D��}hg�_�� w��@�Uz<�g�<&�?���4N�.�߂�y!��G�d� �"�uq�{��q��<y�@.�.�d�ʜ�j�&��U�P��\]S��bX��&���#ySYE.*K+�9A*�q/M��jJ�x:[�rI���y����Y1���,�Z�2�������k*��A�~�sV_^�&�cG�I4�hk�?WW�|,W ��������/�N���Z
0bʮ��OZ����iO����F޾y��+�70���sm�7�9�B�1?����N�����E��%��0� P�މ�����s�j�s=�x>������~��5�~`K��o��� �t��`TZ�	����׷�7TU��{>,�����#'"ӱ�3g��;��kF]�<KT�����k�����L1F�oC�_�s �/�O9>T��"��@R�{C=�9��:�]�]W|*.*�����`����DK/��������~��9�~�m9R��G�=�*d�/3/5�/b�}��}���vDm$�Œ�>���X�m(��O�Hj��i�u����1�⏿��J��{�x6.	�*���lE����`��?�^��T%X�����#ka��h���2[�H��򗿔��Ns��%sO@���c�� %�=�T�a��,�<��<���3˧(�[��d����B�.o$NߺqJ9���_�yU������t�"����fkY^�I���k�+c�����ɣc��O������ꑈy����k9==gU��b�9�P�J���@{��7z�zM�_�N�OoS�fy!(�`����6Vy�cj�Ֆ��?�)4���s����MqB��b�L��'��)�yM��}���?�W/^�>ݓ㣇��\���%mG����Tw^��H.4���u����ýC䓘�w�s�(���7��0&h�V";s�˳8&)�}���?�^����:6e8�a�fsYT�]z��F�vQ��y�K�O�{�s�͚�ȼݟbb�h���֠��+���Z�����-�q��>����jh�g� �\ܷ�n��kS|l��� �Q��{8�LK��������睲���L���P�̤Ƚ� ��LM�dTYe�X�1�K��e� �)^j�%LL-B��gY<M}wl��d�١H/���[�-�k �؈R��g��>�i��k]�Z׺��mҵ�u�k]�7o�x�=���n����'�YA��#���+YGs���y�K~>_4��>�N�|�*���c��g�\�\jQ�����^�
�>�h�����f�j�,6k�D�'�<~��� 4P��D�@Q��A��~��r�S�78�_�U�{�t�>�6[E����{-I�eIbǨs<#�i>dGV �
��@<�`��]��NwUWwWͬJZ��;�f��z�yD��<Oo�_��� �nv���UA�����!�YL�c�C �.�q�����w���-�����܀j��SVK[�+�8����l-`?+�yʧȲ>�{�G���d����{�F�v��F�`���).p��5Gn� �
 
H��~�V�B�K���=�X_��q�X�Y�	�gm�E;�]�G�N�ꨀ��Co�ՠL;-x��^k�O���ky|��Y���v �R_X
*H����ZX=���@^�}�;df����X;�M��Az������y�9u��9�B{����M�� Kj���2� Ć��A�٭%Zn�6wa�6��T���~�p�@�4�~D�;�K�U�U����尿{O~��}]o����Q���y�G�Ң���a� ��QX#����Odc�M@������@�oBR�	��9]�����լK����U����t�:�g��>�y! ���sm�[���!�;;R�C��g����=.��$ʥHZ��T�|�Ϗ~��!k���a���΁���T#��T���h;[����`�6�<7��h5�����O/�%a�ӳ�l����������C���=]o����2�tu��ܗz���i ���h���ݹ'O=�{�[ruq(G�ߑ
X�kN�\����X��nnqnolj�^��ɩR�0�_�}9&M���X�L��Y���������aU$rt�VǧG��@Ò��k��=��Y;������6К���{��[9?{/c}�|2$�hDDD೫�`�X�ƺ���Fv`�,���#f<��2"Ҁ0 �8����Ϲը��V[� `��L�g`J�X?�\�Ⱥ������W���9����c6�������3�ֱm�Zh���$dI��r��Nrn{}�����S�a/�:����tIz�p�>��������w ��oo��`8�-r��Z�PTU0�5y��LG�'�[G���/nH�֒���{�v�doW��R����K�&�#��|�H:Yв�2~Z$���m��j������Kwh�87�q���fCSy����}6��t���=\I2%ɖeU�Ba�y��s�p<PK�l�ʶ�=M�����O���s�X�H�O&�=
y~S\�p�zĵ��D�zM�8=�5k9�� TkkMN��f'��H�=}�����V���ّ��sr��j�t^���Ĭ �u����8��jo��c�_*<ȩ��
8���y�O �{K��I
\�	�zF,�f�D,��gZ*
��{#�U��yyzo����b��h?`��lY.1Al��?�N���K9x���>�Z�ʐ~��sᆄ ��m]wP��\���h�Pj�ZD.���z�P�^¢x/�w��ܿР�RY!w�~��^�z�]ui��kbHg�d� 	b�_�R�+
:���{4������S}��N�nInh_@U ���h"�36T��UA ��"�����2�恩?DF����e���� �����&�}�Vm�?�:~�m�������ݿ��,ɳ7���#c
�8���m�yN�8E�{�l�N�� ��d��) B�9i`�������f�vW��c��$���`���Zk%��;��S�h�Q�j��j��j�mE��ڪ�ڪ�ڟEX:w@, �:�Cdj���\&�T�Ź��')������x ��=�ax7�`� ��8���D%a�X����
��V��'}P�J�%�\)��݌ds{��*�ߛ��@�
h�����?2e�@��a�\Q?w��T�'!�th��Xm��f�BK	TԳ:��-W]���*�K� �.�C៿H�?z6�~(�F5����:�i�*>�x�toXu��FnL�#��K�'ᬎr��iN΄��0
bU��ф�*�y�ba�̷��2e�?�
�$�|l�;���c��R1<�}��j�Dz���b�X�@3���~��0M��ŐU��g�I�A�����m���U��
|:������"�|-Q�βM��p�$|ؗ��n�U��_��=�P\�#��������3>$t��{ѢR��"�Np���ί^_A5�G�Xs�U�A1&0`(��ʌJdv���dw�%'7g���ݾ'{;����)��٪��ى|����l���u~a����t-dsk�$A�є�\ � �Y2wdE�� �<\n4���#���a���z�)ǇG:�7T_��`sV-�k���}�|��6��n��lm�l�]Ʒ_�^.��������I�Y��t��9��Փ'�辡_=�D���_���[Z/�����׬UE�=�œ4d�=��ɇ����}	�L���ޑ����~bS7a-nmo���T�dH���6�`o�R��t$��<�/t�t{�����Z�A�`@q�Gxis{W��g���II߫٨���H�ɂU����	���m���7v����U���m�$aYs�}����C�1N}W����.��?��v[��<a���gR,F3�jE*�2�)T�����$�>��g���@�h�dR �u�	,3����j$�gs��5,�v����ܤ��Z�J�����[��B�>�,E�O�ڏ�<��O,d�V���#_��s���EZ+A����Va�5�9R���s�e{wG�t~���}���~����e,��+4g�s�Buɦ��i?�D?=<�÷���_�x�����zY���= �$�&��fs�2�t���\���S��u8A�[~��gP%|��:tN��ro����W���$x<��jS�aQ��x�}�Z2�^=��cD��d_+�d�ގ��U�����g_�P�@w\�7u��3��r}�gu?���ξ��/Z͊z��`L.�JM�"(^:�e��/~��w_���{���*�@^�O��*�Hbo�*�b���.��Mق�P���t.}��k9=��C*H��wTt`�C�[�?x������}�H����[���xAF�FkT�{�+���~�{���Φ<�����~>�z��z+�T]zA�L�b)�߯�X���MUפ~��}�E���c�2]�� @�'���5�YOZN��ԣ �u�%���Y've�u�K��6X��`G�S,WK��G���k�B�gq�ܶ2�Λl�Z�s-�_���o_K���L.�f��I�k��	��t�o��� &�x����x0��- ��{#���ׯ��#M'�UAQUս	`�d<�������\0�nAA4�y�NHf���;��B^p��i�@a5�iZ׵]�5ghE$Ӆ�oyog-���Z�{����'#��f��ϑ���/�M%A')�Y�Y�	Bϳȏ��T�M�K�f3�)��LY�pj���H��ewC.~�y�C~�w��1]BuG�ғ��Xi��$�����+��S@�{ژ�f�%J.��#�q@ځ�I�Xp��9rȄL���{���&ͬTQTT�=j��5 ����oX��+Лt�(eK�˪�ڪ�ڪ����j��j��j�'O����	_Hf�P �b�a	 �#(Ҥ�`q �x�G�>���8�x�˃�>��P���W?�peT¦aJP�?Hp�?Ӈ�Z�M0v0Wrc��� {o_֚u�/,^�zE y2��V���F����vKj���jCV���q͕�ɗ���B�=�#�,O|�J 2��N=rUEnK�h;$���+2�d�h*AA��x��0���G�"^�_1�c2��Y�m|;f�=A�Y��W3���%a 2��~	����f��AB~ �|����3���_Cf]�2B��T(2���A���8D1
L~
f��
��ea I]�0�"�/���{�O�eacnǀ��T�7�#7��#���:�	��:�ap܅��pb +�Qo���f�<~>�&�̉vI �~becn��y�Ώ0�YEŐV�⇷��V KC����~#��(
� ����d1�v�M ��kR�����h�	�3ǅUS�Y����?|��׀���}>3��+�Z �[�7����
A��v�Z�->�kDv�i�1��?p��yE>��Ǐ���9�Ϭ�b�R�rc|0�)m��V^��֊����g#�¦=zt�} ��W`���% ���w8Me�ą
+�77�ewwG�^�$O�h�>&�Ͷ��8��z�MZ����Q)%N]Q���wES�BI����.��y��!+�c=�T,��������vS���A�o�鲵-���J�
(.���R��m@����J�Vk�-�{��6�t�%�:s�ًD������^ �1�2����z��lߣ��ٸK"k�lp�+R,U��tL�mf	m�������H�"7]��_���&��M��Z�sܔ��=��ޓj��	H$��;���L�Z�㸑��}����ّ壪�NE��|��`�F�B�GK?y#x-��� �������=<����ics]�w]�(�5��Ȟ����g5�V���R)S�p�\/r��g����s��������$\�x�k�`�=���7���$ޗ>|,-]�����-X�D=֟�d@�2i(���l�ܓ�����m�{6#���(���u�<<�k��r���EK�<��EP8f�� �a3V,D\�r�>�9�#����H�����#u�{��[�Z�-kȀT��vS��`En�ao����c�����W�yBAߠ�!<�I|���^W��d�I=̽����� ���@�5�*��1���^+��zK�e[�Y�D:�Ǻ�<��c�{��\�p����)�t>�.-잁W5���wغKx�����XX��������̏�'��oe����~{f�i*��ߠ�k�E�q�����Bb�ާ�{{�e}�f
a�x�H���=SXΠT��=!�m���q������OC��g��{<�7�4���}�`Ω�?ۏ0OM0�H��x�`�ɘs��L1+b���� (���9�x�C��g�^q�Β�{����W�ep���P�2j~�{آ��p��R�C��NH�H~�(F���gy�� ����4W��
�?���������g��a��S�+�����]�K��I����3�5�2Sx��o1u�Z! P|���Y�a.3F�e���$�u��r�p/�{%�<ca�U���"��p��5�h6�j��ÒazN��j��j��jamE��ڪ�ڪ�ڟMk�k|Nb� J�����6�7�R���@_m6��Atn��Zu��0 <@_\���e�>�QT���rp��ԓ�`�g�L���&�{4I=������n�G+#�
�^�T��&�[mn�-�VJG�K̽ ���*v`	!�8�|�F��px�-�Ξʅaz�y �7:�S�{<�!C��Pј�ݴn�U�ȮX+�@h;,��0hj��1 p��R�ʇy������y�����y��J��T�?A����|�)�&rkG�ƀ����*��� �(���#$@����sa�T�Ib��Pw����=F8�$����.�0�2������\A�s�� 6KC��� 0�G�8*������l4�Bٞ���"b�T��*�
�x� � Ud0@%��92��p���	����9�s
�	?c�;*'sB$�z(�f,x��:����RZ��`$h
���r		���67X��ٜ�ÖF�r>�s]�޵#���`��g�&:�����d,�T5�Z�V$$��P����� ��@<�,�)�e�3�6A�C0��> >�\�.�r ��s���F�dT��X��F��ǣ�w�� ��V'(�1��,<�����P��� � �g��^־k�͈�:�+��ic�u 
,(8�? yX��Y[�jXd9j�ՠu�)���o�}P��{b�^��y����C�����A�Y�C��&��7�5U��c����4��|=�Ϭ�g�*��K�)�a�n���eÎ�fs�k ~�eۯ�����w��C�"��p��M�"�|�&}���H`�xB�����\�󋪺�a_(�:`�t���[,�-���ܵass�㱳�E�Js��5Ipm>�p�ٌj�R�쬤,��B����N�p�P���83���	l}u(�t]�:/��^�z�s�R�1{8��5�A�#���kܳP�.T�@I��_
��hkR:�XU���	m��բ����iK��9Ui�QyR 9E0�c�8��
�	�M��)����A�o���j�T �<�Hl�i���a&�.�F�!�v<������z>-ݓb=g�qe�\+�J��d����j7[�U@�֪s.��[��3�S4�A�=���@ҩ�WK����a;}-2C��L�5d!��1�y�΋0FN�T�V��$��Q���?�s���M�� ��ER��"w
{A92jM�sC^�ׄ�j�5ݓ�$������r��?�Z���r>JMinB��kqm�k	������F6`l&z�������I}b�e����x�5��;��E�����E�G
%^nMl;4";6�l�hfT���<�m�`����M�{	�<��'G}I������XkhS����s泅��,q��0a�׎�lby+�3^��ٔ�_��9��~���ǂ������=��[X�@S���i�����W���^�*�4Y*]q��e�k�c��jt��Տ�^ǋ�#���3�u�AjsѸ�[;'����!�����@�L���fc�;��Ƒ% #FLd���U�l?p��S�ޕ����n�GH���;�������%R�g��RSx���9aaPTJ�����F�21�+�D���8�!�;IBZ�</�e��|���.��E#�����g=���/@�d�ڍu�/�mq,��j��j���VȪ�ڪ�ڪ�ٴ0�d��"���C�8�/x8�4 `��!<��
6��d+h����xxÃ��Jӹ�t-�cD�m`�:�]1.��:��N`�Pqx�2��� 0
�����M�`9� Pp�?t�������J!,�v�oz=� ������	�N�̼��D!,: ȷ�ZT�A�O�������p��MY���2�n
�b�F�$< �]	!���������e�@��~�T�C��=����3=��7�2f 6�'�9�����U�Æ$uОovTq�,�^��N����V�'�ZCJ־f&K��O��RA�:� i��`���#!�^kKk}��� Z �0�P���AA�,�� ��CA��,8���6�|_,�`# q հZ�C�M��E�դ���=2B�`w�
Ox�Oa�����]�ln%$
h��gF4��anAqA5Sf�� ��n����rH��K����[X8��������
� :�U�Xa�#��1ϒ�݆���J�c9  aD�Mp�Pт�\���
`\���&A�}��޹~f����,�	�v^�����"�_A�:/H �(FR��@����z� P���;��

�`/PY�����φ��.* 8�	�5 p�Z�(,Ut�!I��z p�u�3�:E�� �Ho�o��֞���)3�w%b�3dRN&)O�V�K f6Щ��T.��lSQ���h�%��M�ʖH��Λt"W�k��Y7��R���w��zE����z��EGz�%��dH[���mH��3���\���,�@��t��\ � �TJ���Tu?}�����:�Kڿ�fEϧ ��E�`p�:6 J ��󑮴��� `>�_���R\�=�$�]#=6X���;]L��SZQn�k��B�/�����^9&��H}��j����{:�`#5�z1+�^�����u�� �9����KU��)�Oٽ�%{�:�{zΛ[R����Z#�е0��Y�5�!^;�5�$fH���2�>��1�[2�e�������Hǰ�>A~r'67y�1�l �؛t��4�H��7��@�(�dwgM���o�^c:�8�~��Ҝ�i }3fT*���K��kb�g�I��ҹV�^w@R��x2!��u����9��g$�jU�*�R�Ll�ҿ�i���]�>�+������:��5 �f��8XY���g����:�(f����q9׽�Q-Ɇ���KŪ�t?� �	��b�uXÅ"��纇@��*Eu�����-����9���%O��o����.�Ek�I�(ұ���C�ě�}�^����?Wz}��L'���y��C=�*͈k)������Ƙ$x#}��
&z.�@�v��F����M����Y� 2��N�<#�Ɇ}i5��cmc�b>#|J[+���ލ��i�{ĸ�`5~�k,.t �A�P		e`���hj,XL!�(�e���4l��d1T�����G$#��e�@v�p~^�<�\[�" T�����z������O�AS����}GhV�$��^����GK2g��N��T$�pߔa����\4�O-��ƴ��"U�!WPy�7�%�x���ոG���a�ԡBɬ��
z-I��y��c]�s�%���ްӳ4�}�@s����H��}_�o��H��qzÉ��av��G07Ø����`��Q��m���a���fn'�I�D`s�eT%9����6�����z��w��e�!%r7Hbǌ[�m����=���$��/'�W��#W&�,O�t�`�{=�"�_�L&�������Ǉ���U�?ZRm���)��U�_����v����˪�ڪ�ڪ�Ŵ�j��j��j�ӡLU�x��v;�'�����bŖ>����]�F2�郣� ��8�	�_�d<��P�1T�����X�4 ��o��7����E6wA��	2M|(���AOʥ�|���|��G��%�����]��5Nd������{.k�~ϩU�B�0���Y�!�p�JI���җU�É>g��>����Q��@�y!���O�U������L���Ȩ��\����c| B"*�$n��`�6WP�@�㣢���OnTq�&�Z��'�dFb�J�[d| �H���U�VN��� e�� n�(e����ݰ?�B%F$��c�3�Ul
�t��`݄6	���ȫ��r$�f� �C�V�A��p�B�Z�&�>t�� m��Yy{V����91�-���E�eZ��	_��_GR��)=������ 0���G�5���;x�[�.8�yf�&�K�S�
/�<�}�96N�@���Y� ���1�0���b �YX�je���$Q&��	 { u�_bs+*�ӎ�DRFT�f��b�r�x,�����,�dW�c����k�"Bu/��G�9-�P�M�A�!�υb	���'T9�� � z1OP5�s8*pn4�p��Df�Ȁ[#e�V3����UC!z$�ne�ϴ
r�=@I1�Nń���lAuIM�!��a=�m`3_�Y�R ʀ�GLс=A��w�&c�c�/
$0� M�)��Ĺpw��_F�m�
�:�����7# icd*Yk�a�I	������Ng��m���!d�F:f	� f�h2���U=֐���9��ַ���} ��	U�S<���+e2�&�c�`c���,l@��$�6�����qO&n�C�;UiLL�<�q�P�
@�w5�tpSdT����p��O ��(���4��!d����b���*:��� ��q���T�a�I{�E���>X�L��X�����@�V�1�:�k�b:�ZeS��ߓ����D�S�,-����&�h�r���Ԯg�+0�
 �'�ΰ���(
2�� R���1���#����\�������o#�*� ���u������8���j=����}���	��h ���	E\/�:5��Vy)��5���ε�|���s{�٦
�����9D�^oH&zPz짳!U3�A�B! �=J�0�i!��PZ��Jn84�$��bS�P%�.C-rYOܛe�O"��s%tװ4���n�l�4_:f�~
,��M��*��i��������2��L]���Ej+z�c���	xſ�½���0ۨԪ�����ײ�|"� ^f�-	ψ�Ľ���аԄ�d:K��^`� eŸmܥ�z��J���"�h<�ybv����b�kP��-s�Yy�9����q��.*��6�l�@�,�d��ٛ�S�8{.�dgn��D�(?f���e}���ٱ�[�'�˟���L�����K3�ݟ��dFr�9��
&qICS�x�?V�q�-�Ri���K�o��9���'��ֻ�fӛ���}>��$���ˑ��?���u�=��{5=�f�$5�d�Vm�Vm���ڊ Y�U[�U[�?�V��dlUii:�Ʃ4���l��Y������Z%k�A�xTwz]���|�<�v�t �.��YoNP�[�u����
���i{�a�
D�z�YJ�	�V����{��0������ �LY�8c�Ô�$��
V����4s  &��r8P�Q����,� �o<��|�? S��n���M�ϼV��{��~�?�In4�^�a���gN�
n s����<-�氣
��@����S�_��e4�g�e2��r��WY���@�r� ��%����mX����-��6�����)�|��E�,$`1P�Z�k@�@)��]8@%>�����@�6�2w%o�c`�T�;<�Cm�F�M�|�؞g������Z欆Hr���&�J�"��wAզ��P�ZE��9�
c�j�6f.�"���&-?f 7�)C�;�()�#��<�q	\д0�6{#Y0g��ڋj�(r4	�� cf�(슢� #����kaյ���-X��G_���#�����zł�l&���_���ޝ��������-�K���dKH=sղ��e�����Q�}��o�e�U�[e����(�ڬ^p����yR�K�? ����elȰ� t�,O,k6VXo��/ʬv��c`P&E�9Й1r�҄�3w|�1^X���B�c��6��E��%�8��!7�/�j��*�t_�u���8�f�����p-�h��l���ٟs�F��������%��E�{*@_g���|����@U`_X �c�G�P���܂���fS�#��u�� �m�͡z�-"5���$�w��nȃ�+�쎡�_+ːJ����E���`��(�j�B�F�L�l�`�<|>���7R �6(�����̦c��b��P&`J��!�;���R�u�fs�`���������Tf ���e��h%�,qQ�Pv����F�vDz�Z:ᚇ�)���lC�Lʱ,7:���2C���aT�!�ٰE1���������Z<��1�����k$q�L�@䗸��5�/�0B*A�[Hg�?�w��^>�~��l�E�C�9��`3&�9B���PP�Ĝۂ�	��vP�X���X�@ה$>��(.p�͙��=1�H@�F���y�a�)��dl��Vwe�7�b\Ӑ�3�ͮ��"�߮/���X�s�5؅&$-�Y\Z�T@�a�,!#.^�o�K���D�dF%#��̍YB�T @<�=�	�h�5$����	��S�����X���y2�An��ɉ�F��-��zi{u�����3WUZ���ǭ?M5�kn"����<�~�ǵ��H��%,ppvP W���]f܀j@Xd�tr��p*����M�Yx7��f �u?��	X*�@�@-�����y��NI�������#?��eU��g�6g|#&r�p٩�t��{�����b��P�f?��#�{τ�[.�]Rڃ���T�y,����Ȍ0qv��%��}K�����dy�����A����{րe��]N�)�<�3f֫ �'~tt��EU��/V6X��j��jimE��ڪ�ڪ�ڿ{��?c����5����3Sn�-xpO\�7m��`i� �* \{��iP"�$��xYŇ5���zPeU�3_\����P��������P�\+We��������`$��O ��3z^�A�*e�>���p\,��ힹ�k��O���ۀ :����	w����t��۷��p=���#�$
l���Uf��H:z̬�N2��J��ҹ˷�l<�`6���ၜ���lo�aȻ2� �M�X�N��ܸP��d���e��8� �̮���p<��X2�����=���d�0���IJ���h�y�X���к�� �$3�) UF���5	<���s070�V��c\8IJK�<���N�V���^�0u�9;+Zi xrO�W��{���j��]@��/pe�xb*"T/��l�ElW��;��s��T=��@�,�q�Bs
�-M���q�Q$	3���#!z��TSs�� ��u��/,��ђ	ǞYR�x17��q`�E6%@��Q$�i��IzK8�~��D��_�����SY%5��� ��yy��NA_�f3����KҨ��zx��8�{a�.̏�y E�sL�41�Պq���Ԕ��7�9I$����sV��Y����-&� �=K�ef�$*��kz�/�6��gv�?�/A"�~3��cL�����!��@��TJ���K�so4J��%T�t�NT젚o���� "���B�t{���OT�c��7�B�{E:&�ji�/�>c;�A;sk{�d:#���z�f��.C��lj�_N�dyKzN��`]{�T���*�U��s��Y��ku����9�����{�#YzC!*�3T-��J*�9`��iD�$4?���e�` 1&��-�|}_�|�W��ڇ��A}�9�}<z�� Q�3$e�<!����t}����҅���~@��`%lI�CI��K{+Z0y\���.(2�7+���]�Ҝ!�w$�|�/�`�U�L�ɰQ�����wrrtHr�����B���ʜ�B�:#�Nz ����7�s,����o�$��h"��@�����.����lf�)Y⬓�M�vW����K^,{ȩ���J����x�0R��kK('�"�{)��)�`�^t1�PI7���M;��.�k�ӄj(Bg���AU���x�k�t�Y���6�yLtࡊ��P�R��/&F~�~(I�.�'݃
.�|27�	�@�z�l�=��CRSx¶�Y��ЏP��_��:*���L�ȕ��TY�އ�\)����z�S���EѬ�0��ו����h�?I*�c��u�b�ܒ�� D����A�S���Z|Ʋ�����!I(A�����L�������:R��0�?uφ� ��TM�b�a��0R��bdI��#D�sg F@��S<�1��5G���	/�`����ę,�<(�C��N�����J]���F�Ȃ
@Zsqv1.^�:�N_���*ЎǬbM��Q�>�	q�	��ȝz��T��>;M���:�5��sS&Q��k��Q\!GD_]�q�=�W8٪�ڪ��_X[m쫶j��j�����j$~��O��z9�HMZ�`����t����'�^�e�8[���%���2� ��:�>lP���X@M����J��|<K�5�X�(��d�W��V��Z��h<��w�rxxL�>�k����ƞ��Z�����U�S�j��4oAPȩ��h���$x>㱫\-�w^���FZeu1�=f�	��d{gB ���L�����pF�:fesU�c:MH�@�Ͻ��<~��ո��Z(pss#�~�������!Ь����V*Re��<|�D��|%�'��+��I�*5	ÏۑV�k�޴�#����k_�/N��V�V�a噩;8'H$��z�P������P�����U��C1	�R��X2��X��Lb�3���(c|�9�"��@(�q�s�Hi���z�c_,;& 3��%V)������J@�m��"�#�6nsg��;���3�x�xԅ� ^HD`A%�п�u�x<0p+�֗V�b%�"��Yq
ذ P�]�v>���I�s#W�2X�PA0�%��Z�`Ap
 � l��"�k�s�F��b	�������bL��Ns��V|���64���h�"�@i��l�ǿ���R.�>��8�9��8\����~�
�a"���} �r�߳Z$Ӟ#���$�ܰb���t�� �m�t<!�;eMD���{%�v@$�h�4����A`}�Y\�\�pI�1������L.ί��#�"�W��1�����(��)�G��:��΋J�L����ə4ڛ6WRG�D� ����)������t:R�ڑRR=���؀u���=/.Y������}���+����e��,�%�������\_�ӆ��p@RY��i��2����'���FMf$f}qq��jHB���92>�]{�RY���\�\Ӣs� ����J�֖�m��u�δ�cl3�"�j1K9/_��W�_�O~��^�t�I�~��.r��T���&�ą���z,�ײ�� �[.�$�Ȁ=&S�?����@R������B��?�Zh2�s����!�c����#-'�N�F�Y�RZ�a�����=��������ʻw�x�{���ln�Ƚ��Ҫ�%Am�Q�}�3��(8x��@���4[59x���Q�E�- ��}cս^�<ߨ5H:�:���@��hu��
*un��}�3�H�N�Y���
�ı��:Tmا���aw	���@ϻ����/S=���L�*����F�>��\D�D@�++E^�ưW^��+b��©�; 3�0�qB5�٨ͨ2�M�Pf�u��+�
�0�}������m!���
�P-f�}������K���b�U�%����˛�2#��I���ܑ;�S@���;�&��`访!H���A�١���Pz��{M\}��K�1Z�Mͦ��L2w�av��N�w6���("��X6�x���/��m��ݐ�:�H�:�������n蓉�Bعe��_��l�Pt�D�9f
�e�:1�]۫;�������=��������;a�y�_gǒO#�9n���ȹ��x�}
��3�w�F�܁���X_�h��:}|���T� �ao����U��_�=�k��F���T>����V~�Z���v�Vm�Vm���o+d�Vm�Vm��,����d�0R�Vy�W�<�z�[uwt&?�Y�}g�⼏�!2����t�8��1r��9�Y�k����p`%�`q� j�ȁ_vK�F2����9�]a����ڱ�ׄ�t�e�<��W����Blj �{�f��e8&Q�����@����>����ߧ�	*F����{�w �~�L>��9?����,}V4Z��ӳ*M�������+p������6��P������_���?���+ҡ ��aP[K��9��]__����?/�|��$�G�b�9Y�*������ʼr�*0�_\�˃�]�������9%!p�@f`0�!dT�`<��>cX���)���q�}��	?<P�}�r�U~�q���3�(;ϋ8� &-�V0P@���7���@t����#�N�c��z�g��,�.@�����D�l
�����9��lJ�$����� ��������f�����[-ڟ�|6�Ju�y�j��ʨ�L��Vt�o�d�^�j	�>>��.������a���m��Ȣڽ���	���BI��*nx��&ȣ�����������\N�N�~�.�R��# �ulB��{n���G_�����7o����}�x�����zP�~D^����|V���]ɻ���\#A�Qj��e��K���� Bu&G�'rr|*;����M�s&q]ൾ�kz�$2�5C����Bz��ﵥ��o�N%Bŋ�%�`=���I����˰3��Z��߽��9T�0�C��Z���>^��D�?<�QIJ���۲ti���\���g9!	UWWWrqv*{K�%=_�̉S�A���z�N ��,�u_�;�ׯ��������7ZT�L=F+��D �u����2@nG:��#]`��|�f�'���p�V�Ϩb���)���ё<��<���%�G�3i�R�5��EItܮ�.x�T��!�@��K�y��ҹ�Ph���X��ܪ�ӹ)�t���8���ԗ/^��>�������*4_� ?36`;5J�7�1� �P�9�OOH��J5)W[گz��~N�1�YCR�}����������]ʓ�H�:?����]�K/���M�\A硯�_��ZuM���+��r��R	�>�X���N��ף�1��zMz��{�[�����Y��"�:ѓ�fvq�΍�}'G���)����F�l�p���]�Z��@���Ľ��ױ�rxx��+H�R�J�ʥ�zXdR�73]z>�uXZ�����}�~��Z\�������K)V+��ߑv�.���2n0Ϫ���3� =a�]��Szi�R�����K�Y�A�}U�pnj2�Ttr�	��0�I2$䌬��V�b䇞2̨RC�Db�W�rI��o���
$ p?�kD!.�>�9����1̙�""Nqh�Y�7���&ӊ���R$;�_�p�S?r>{�!fa�b�)*ㄪ5��˕ �1�'r�R�G���K8�\-�sf�{�+�d���3"�o�υř�f�+@��=Z��Z�9�dʜ�X���ֺ<z��s�-�ZQb�k�;�S4ε�2'�##�tf�P}$#�#\+0����q����BY�},��]�%>�O��-I��?jw�"YnW��'{玝�[��V��+�0�����c��Ѳ?Dy@��8(��S<#^h1"�9q�,�G
YS .\P��?klb�z1\�Na�f��Q�xs�[�+d�Vm�V�/���U[�U[�U��h�8)o���(���!%�PC����A��W�p����F�E$��:P Y Ó�>e>�H\�BAE�A�����Pd��?K(&�\8/a�`�\ч�JP� E�����x�m��F�0�@R���G�l��:�I8��cP�=�eޞ�[E�uy�U�h766d��6�T�_\\4*DD%�� �2*I�Kj�Bo�W�!e=�2U! �d�,X!�ȫ�o����U�'zl���������Y���"A�Vk�؟~�\�o�2��evq.�ۻ�\
��$� �\�0�|.E�  ��IDAT�7W&�e$�F#6�g��<cp5�`f3Y� �
,'̓VM)�� 4���B1s�]�Rb����9LiC�p6���O����,Y��.:�Ĕ�3x�-	����8�.+253�Ìy*��\���� �Ҷ&we�X���qoȳ@���5�O{-Gڥ���v�Xh��*�.�/��E ;���b�
J�n�to������ ����gT5�[Ҭ�d0����ϰ�J$�N����ȍ���/_ȿ�����Ï��^#0�N��C�MFOOD<�s�ίh4�5���G�b?����涬��7��B�<*�a#�������_\YD��݁�������Ky�ᇴ�|�q ��(����s��s��9<<����G��>��k� ���M���gg�q����*�'���=8�O~�[��_�dmcSb]���:)WK�{�I����	{.�9<8���������\�$(U�O��ǹ������_��� @�d2K��cY�R�IK��d�?7�(�/@(���^��B��T���٥|��72���䧿�zcM�`�k��g"��=��ҽ�j3��aP��`$o߼�{��������c� tρ�P9 �y����/^����\����3�u�� �,�#����o��woY=�h�}'�}���Wy����b)&��L�+����sy��')�rC�e؛����\����Ώ	���O�R�d>�o��N^�|N���^в�T��/^�V���.(P�a}�`w�}��\�����^���ﱜ��_~N�܇�D��Z:"�d�����<����� �����|����?��g���K:�1�	�Vd�_�ɳ￣�c�}��~���+y�ȣ��)�&�r�M& 9}�s�L��`8���vxx�φ���>�&��%��O�H���z�J�^�LH��|`���_ ���u�|�b�j�/^|/Ϟ=�ˋ+���~����_}�c7�_��B�<���fT�zX���X|��[�3��3d�������?����GR�6�O���P�Zr��J^�|��}�9˯�����?2�o�������fC�Q�����~���S��S���j���ot=l４�*Rno��u�%�1Bf�0C'�sv�}���39C���O�����,��Z���U^�`x#+H~h��ށ�ZگXk��Z����;��4áٛ��,D��o����Z8{I�.Js�b9~��. �z��@�����h����R�Wd�2O$q�Y��X��� �)���| �q~3]3��X���$�Q��ڱ�6]f�5�׌�{�Ֆ��lo����G=���������G�X>Sfj��=������)?&f%~�1C.'��l�,'-\�~l�i?���[_ݵ�rmI�,�0��"N�_�NYz�A��Y]��LS�f�w����vX��|S��nn���R^-i��c�b&� $�s�w�G 1�1��6���~/t�5f9�o�^�+���+ݶj��j��j�s��j��j��j���j���x��Al����8�Ŵ�C-ZFi^�3Z3�
���2����>�iy��r |X����s�� ����sqi��Q��M��7�FÉ�w/��� 4��[� �ա��Ys����`���&}��� ���m X�v[����a���;�>}����u�U���K�*��llΰ<I�X���jTd�F39���o�}'��O�<��ﮮ�Y���љ��w�R.I{� k��}]����ls�ժ�MA�þ�'�����\?Q�����[���;au:U4!���9��x�N�I��%�|�+�ǔYV%��W1-	6�5R����O��b>��s�g,��ѤfeeU�)���5Zƅ0X�w!�t}�l��i��Q푫�R��!�G���Xм���~�W��ʔ��~�3����L�Qi ��Y&SڀL��89	u,�	��ַhႹ��w����W�򅎵�����4O��V*�����WҨב��y�5U.�H|��}��9=�$yqtx*���o���;�����.|��Ul�:���g$��PEq{��k�:�_<Ie�������G��_���Ke0J:�3�����Z?SѨViYvptL� Z�\��J�Rӿ1���"�i�����~.n��/;�=}!��P~��D:�tn��^�Ft2�7�=vGW�7��_�0���~)�����V_X�s��L�w�r���z{S�O������*ǧ7����*�?�H
��lD*�r��J�>�Vߟ�ͤ٬���{� ���'A��A����j����N���_�1,���d*'�'2�d��d{g_66wHj-��ϣ�\��{z�3)Bi��H��o�_�X*��?[�-��B��A_�:m:H�1/��#��	����޽{�l�hm�l��u���ӧ��L�f�Yӷ���ō��?����d-�_��Ld�u7���ۯ������J�H�����u�B������z�R�פ�j�Ü�췟�w߁H8�/�P$񃹆�)V�T��e�ׄ�ܞ�gtteD��ohE`p����ɉ�����������A�Q�/�G�嫯����Z����v�r�ה�|BR�����FK�R(e��I&c]�G����ryӷL�97��Ώ)��t��_��	��h��x�2 ,s����Y(���<����k���O����C�y�������>_M���w��A�b���ߗF�-�Z�����{���?�`���Z����@�ZC�&��(,VHxԛMΥR�L�5�BϞOu
m�����+6�rA��]�Ծ�t]���2&>�J ��;�_���q�j
E/^������Ήz�.�>ib{�M�J��)	��~N����$�@�nn���W���1�50�oY �pwk��#ʰC����V��Ա-G���	���D���?���@N|�/������
 >��-ׂV��L[PU9��X`������*��
�������pc�U�n_L�>�Np$1<�`5Ց8��ު,�^�rAr%0?C�'qyJ~���Hl�$2�n��RTi�6nB��M�+�����l{�)s�>`�{G���9%$?t_�!�e:��\)��Ζ<~�@�? �\���/��)��[ۯ`[�H]�y�(%�j�B�1����ܗ���ލ��ۻ%���%D�ϗ�G�o��cB*��(F\F�����o���d�o��y�;���}�Q�k�X��qsH��[��ͬ<'��e�Y%b$R⛅r]LY�ZV\�b��(��B�;�����3:�^����`;� ��i[�U[�U[����"@Vm�Vm�V�Ϡ����^�=���ܗR�L�0���?[^�ϧ�J��VK�QׇUXǜ��
�AJ�����x	e'�S���d���
�e�x =^�e2F�猟Y���V0�t���^�ߑd�d���|�n>q���a!`u�j���fխ 6q� �Qe>�CsB��+}�e�kk���!���LN/N��+�Z�N @��#�g��a��� $T�'��J��S��~syC06bh��ՐGrzy����~*3���`�� e��D�;�Ql�����+����*����?����?���ꁇ��-���p<�R�B9T��x�o`�s~6X�# �{<ږ]49��,�>-e�	�݋qY�G�`O��!iE��,�d�^ ��C�EbG���r�#? �q�$P�5CH�������J%,ZN��@b�fOn�>h��g�V#�R�'T*♲}�j\��)�b��ѱ���<������BQ�D�*p���L�YB2&��QBKT�_\]�t>����yJ�����x`#�*������������RE�/2V p��g����������"��u�vn�ͫ���=ט��s�H��Z/u�We�Ք鸫ka��t��*�.Tb��h����/��)WNt��ֹP���	�¦������>����,�~�A�Z�9$���D������zÊ�vk]�����������\? 3ƕ�N�9�0窺/ ;�Ѭ���
�]:PO�����8��i��BW��3�S�͞�P���E��ѓ�7���������[9;���������v"��L
�Tk���#�T33���l*'��r~u)W�]2C=_X&��-�2ϲ�=|"��:�bl���@���������<2X��tޕ��c����j��S=�u���9;>�O�V�c��،�V�wz]���+=����o�������PN���J1�"H����@n�����#���cݗ>���=yx���َ�Gy���Ϳ|"_��u�P�T
�.\K����h�&��A�����������'/�?'���s������u_G>���5�כ��ڠ���ρ�����Ї����d��]&p������Z+�2j�k�pN`��䄹#؛��Ѫ��LYPe����=��u�o�����wo��o��-%`_�m���|���r}y.=�5|��#6oN�ȧ�~FT�X'��^�/:T7��[��7���t�0h(:�?� �m�G(�p}888�q+�u�\S 8�����Q�s|t*/^��O~�)�Th���x~N��^�@�/_��97�k�gg'�������{�T��ӑ��?�ݝ{R�u U


�7V+uۏ�	�%���=�+C$#u^"_�����KS����V`k��ȅi�|y�s6[Ǉgҽ��Z�5|ttB�*�j��^�
���c䏮X��^�w�����?�Z� |I�2���3i���H���M��r� ������O��g��鑮�¨�{ȍ���<~�����Oa�����20�/���x� t�{���ͯ�q��dS����������Vݟ��KR�)P>�Zd�*V�n��8$W��ey�����ʛW�%�o3��
$���),��#��=�NDK��:7��R�
)2�xȾ����e���'�ǉ;F��a*;l�H��ԊW�d���j�2r�П���eM>����辄��%�	�v/��H��T�9��B�A����,��c��e���rW�������/�@�V��o5?�#��KZ��*wsA@~�r'�CrK��*]�_��=ONf������z������9x�#��S� �O|��Kf�EՇ�T�`.1?Ɗ:|��{G�\��ws�-^�|�����*����kyck�,��j��j���VȪ�ڪ�ڪ�Y5T��]���y>�j�<s� �<}���P8;�p pU���F��i����h
"�V���@Z5����rE��i:aŧ�'����6,�4��#�{n^��ȂrZ�z9������3��θUgx ��ZkR�4�fzE�@�o������rU�mC���K��$!qx|$7�+�%��DH��0�n��BC!'�%�� �d1c�B{�%�<$q��H^�y��)+��7[%TC��@L� �������*�B�L�R�20�V)K�!�$}���C �,�{{<*ZR����k�
I&�+1����K�끩2fs����_�Ǔ!		 a��g����)�X��l1PM�y�@T��30%Qnk��#Y�l����Wf�ǪELST�BiAp�U݁�;�m�����i��(H-���1�ʒ[�- xf��d˫_s;�=��Mc�^�{�pa�p��xH�
VǦ�K�@�*)>ӽ����9ZgU*��y���p�=z�1`���3+`�k�R�q�����.Qa	���'gW��_�5I���Mft�� *;�}��]��m��Hն��kr~ѕ?~����ۑ��]�W6$j����w�������:��X�ñaJ���2��ȫy���U�����}��|��	�%=x�F#��Y�A"g��l�0H��hIP���\���9x�c`�h8�@����b�: [�OG�����c{Te�J{E�P�<>:�J�/È?�����/_���V��1��~�{���_j_��cڸ�q&�f��߾����:�kM�}�zEz�;��� �!P>�����&���=���3i�ڲ���*����F����^���kVC�*ýA*��
B�^�>��?�� }A�~�VgF�_|.O�~+=�r�-��
x��l�ʵ�g�;�kmٽk���} �a���[�)XX �
�"	6�C�������|F�@�X���瞁�������N`!�\��5��`��_�u$
����n6�������M\/�>�N��O	#_	s$!rA�z>�g֒���|�5��P��Wo^qU��lɽ{��:��1a�G���hA�8�]�8�t���˯�� ����������J�y��*@Q&P� �� P'�$����>�~wH*�@��r�!8ټ��kƺw�l��:[ )>oR���~�χ��n��� 5$��9ö�yu���.��є�� 	�� �Cl}��������:�999���x͛MQ���\ �T�9�,�˫��������:��ݡ�����B ���k���0�>4�(�S��p&�M��
�T�:�@P���$���*ͧ_#7������@7��Tz���|�<fu�u|�o?�5�GN�t�-"�W�nF�K6�/^�s䑇���_�o3��p ���g�~�����e�����������8� �Bݳ��1E.�NE���Jv�̡��.5 փ�����_$<G.~)d���R�yGTP���O��^Ӝ��	�U�S�_ ?fqd���ʃ� �.��Lu�BF����[��-u
�4M�,��/ŠD5�x2��H)�Ǒ��+�T]G����0���T�T�Z.I��2��RD�U)�>��D(T��<L##�}�������K���@$;�0����r"�OIϻ����^n��������2M�Db�������o�(�co%�91���#�&�����<� �/o��
����7m�,���[c���3+k�MpD�4�Ƥ���|ӧ��f0I�t�ZU]K.�[��[渟{_DD3����BvFFĻ�ﺟ�纔m�d��m��j�U}�]ѫ�R����2�x��⦡�
�X� �:�G'g�Lv�����Ï�ׯd[�e[�e[�,ʖ ٖmٖmٖDy�굥�����ĆQh�IJ��3"f�4�.�V�Y �A�������oI*���
F��,��=d5 ���к�ۑ����� �	0a�۔�[�Q��� 
!���  &g�3{#r�(�_�#=}*���<y���1�jx#�x���oo�e>�x�D�$�`�zz���`�h\�ϛ�=��x����G ��h��RW<Z�$�@�#�!~��P��o�F>��|��7��__2ҳ��:��M��-mϓ�'rz��Q�  !�����^n�����H>��3i��_�v��6�/grݿ��n=xJRQy�]�3J�prJx���p�18p��8GC�dz@A Ą,z1pm`�
eEb����7�A�M`<8�`N�g�_� 9̷��3Q-�Ճ��s��T�� ��X�58�o�ծ���
1��"!�s@ Ո�$z:ıR�钛TW��h�)�U�pxY+hwd* C(�j.�
c9d�:Ĵ�%d '�z�2g�tz��ҕ�~�F����h=ih_�sfp?`��tl7jM*j�t޾�z���HCV�7���ky���|��'�����/^2
�I7d6/t�/�8�Ӣ����/���F�>Q	��O��W�����O.����b,M��h��I�������9=&��D�D޽��1/��̰�ӦM_�X���]_�y�R�t�yN� � #��1�%��=�r�6F���vz��Mp{w��T��ي����W�_�Zי��_���y�攡988�z��W_�?�č�=�����M����r��4�pY�YY=�y����({����<=��gt���s� 	D�΅�ƵA� �t����o$'p�Ny��{��˯���4I�F� ��QR���ǈ�>�����	��~��KJ�(���B*/!h��q�����^�}�$��	3 ��������K���MѢ\VM�W&�ሾ@���r���x0!�O�b��	�)��.��^�7��s� <��.��@����:��$�Zz_$ʈ��x�sm˧?��*�sߚ�[h�����`+R��a|!������� >|�����ͥ���\�sB�~�� �Ga��0�s��|!���oI� Ol���?��C
�_ d�1����B����_���(��{�c^�G���ZC��ֵ���ϟ�s��tZ���%G�'��������0"Gv�l�K[�<dr!C��%���#����K�$ҿ2:{o��T������\���е�\���,�������u�;�rcnh3��d&��BJ����	�q��	�´<t�.�'�?�̙L�𙖖�#�f��W��\��\0�
>$���w\_�#IY@���~B&�1�oHg�T���d�Dד;�Ab]X�� �	E|v4�Ө<�y˽�@V"��P����Z~��_ʫ�W|6���)%�����y?��Ԡ��"3��D��x� ���Ea_^��A��?���z�{������
�*") A���{�~w��c\�֒[����U�9r	aP��cO9b����0�\!�[�b�t@�3�gq_͙I�YE���狅�J�;q�����9V�(���3��!��mȏ#IO��d'=9�=��}�$e�YƦ���]M�W��ŀ^/7�w	���t� ��2tҏ+#�l�o<9���]���vc� ����DG�e�����^�;�;"Ɯ��u|g��[��	��g��-㟣Mr͢^�sI	K	t�
�_�oP{��)+���RN���k���aEt{�R�k��5�����ISo�@����:����_�|���˶l˶l˶�ɗ-�-۲-۲-?����p�Cq���b="�1d�>+�N����q��a��ٕ���|Y����!� z��#;���C����+��䓏>�<$��_N� �I4��?�{�i�2�p*��u=@-v��4��롫���G}$?��O���#�Aj�@?
�< �����M:��~_,������s.�<d��#J;![�pQ�iM��Ș�$[9)&��G����A��{�C��U�ْ��C��g��<y���G���oh�2CeAo�TϠ�ld�n5����_���ۿ�Z�N�H[� ��������v���ǲ���&��)!�D�{�/�	��0�G�F����g��$X�!����Q6�i?�#�M�*ad�	����y�e{�uZ��������ba埊%?ߤ�~h2���y��٤=2�a�|���ץ^c�yT�H"4�1�#[})�k��! �n�$��^��X̐Q�&�1��0�Ɋ�����cR8 ���)HX����,9�c�*��b�I���##i�H��'�ƺ#99^��A]�־^��|wI	1q-m���H�R���ۻ>����Sfs ����^� di�7�r��-� Li�=�,(��X2L9F�cy����w�eF��W�Z�;�����ԙ�2(;�~�J����Q0���9��0��z�+�'��BI+�ċ�s�7 ����-� 
}P��J��Eiw�B$��e��9����;����d6%��Z��1��5 �!Y�ŗ_Q2c
�K���1H-DA/���K�EI��!����ݿ��-���36��V1�Ri��4I���/C�?Zȣ�=J�}���rs{O �$d�z;M����:�-K������`2�y�Mp�녶�Uໄ���w��\??�qVbN�꼗z�E$�{��|��ߒ����-�ᔀy�c,�9�L�\��ע��pi��zs��� �rH�@��|:�&Z/��`lb����ٗ_3�� 2r���M�X�aCH��y͌���cIj-��>�` ������B6"�A���> K#�.���ݻ������3�� �9	���}��ε?3�� ��]]wG�=`��_�5Bf"֐� mD	2�2:���C�����~٨_J��+/u<��Qp���v�yc���~�	�q�$�tG6�����O����C"@�c�F�����Z��c0���
A�!K%� LG:���)�͡~��_��hp7��8���� �0V��)�y��I�`_^�Q�BuK#u�>�K+�Yv1KX��7�u���K�%��@Z�$F��}#v~�����ԡ�1�KM �3��!���W�f����z(&�÷�ޠT�d�{�\�c2��ѫ��c@��2��{��;�6�k����+H�i�t?H=�歅�����p�����Չ��
{�G��I7�{0&���HM��|�s�3��u����*Ȳ�~����̲;�AU��'��j�,*_.+k�q3�v�]��j\~M��Ο�SF̠td�q y��뜞g3f��}M��v:;��	R����4}�$v�;S��IHg؀1G��Q0�;zf�A��F��1٫���Ϭ�6��7ɂA)����|E|�=;|�:ѱ��y��'R8¥b@ʍ:E���}�
��	=�e� �s�u1�#�G�_s�� �;H�$����@P��3�1��D߃�Z.����2��}�q�����K!}u�?�襆ZաVi��o	�mٖmٖ?��%@�e[�e[��_����7o�u HT����C�|:4����ς��1"�;��rF_\^QR'J�THh �|����0	�G���=J�\�}C�& ňD�\���x
i&����D^�#r�(�����8=;���]�s�@�;�
�O��e��b<���}I��8���#<
z�,(���N�E��� ͖�^������s�ϊ���̇��c����k�䓏hΊ�T��`^��#:o��I�ERo�R�:ߖq0�e��������4��w�=|YΧ�;�0�P�(�z� x��7\�����FȦ��	�5f�C�4;0@BJP���V� Ȓ�y� ��v,K�w;Cwo��� �"% >�i��p���TF�U !A�(�:���4t��9���I�2��Km��Y��C�cB��e�D��d-��>>��%ސ $#��N���r` �h�X#��p��Ͷ��	4�S���ҶCdiHD��&��7:�d/on���J�m� �����gZODڂ���B�ZjshemU@bK�h�� ����ݧ_ϻ�̰�3Ӳ��C�� ��ݣ��xwwOv�3��;���?�����A�	�ԅd��&:6=�4�յv�t0O�l��ܘ���cƗ��`�lu���e�3��oo鿃y%A�6�2g�
"�A�q *��l7(+���W���K�[ H �&�,��I�%���6��o�?���/���+�{�˂7�Ɇ����Ż�wD��fK�:�qA�g ��7����2�_fK���0 �אZX����՝��� ���R���}�iB�? �"o�L�4!����Wo�d��l�]���3��� � >c� �������к݌FR����R�hK���t���S?�B��l�x�I2��w��`���`m�����y�����$��{R����h]���G�Ƙ�d���ϖ$E��`�b\гEפ���K�����  uIÂ�\r�i9[9 7��e�����[��o)��h�L�9x� ���=2R���'1����F����=8��t��~�h���0$]&(�H����=�X�:����u/ҹ6��]I�+��#�@�fS�����1�?����k�/���A�� ���r;$����0�{tj�VK�GQ�1�k�Q�5��Mƒr�m�OC��D��¬s�L���u�׵�	����?��Hr<�͑�Q�}�v��������h{�η��̹W6��5�M�o��@��m�~B Ba��9`��qZV(I|dP%�9$��j�t>��1�15ҺL�+��D�G9`-�7���#]/J����s�/̝�x�{�@�/oh���*H��q[��6t��O3�I5ih����F����Yƌ#l2 ��_��x����b�b�i���Aꃌž���-/!���2k��j�����,X�0Y���ބ˭ʘ{?M�3���V�`�RW")�y�b�_����r���x�J#�oU���RD��X`��:���G��9d�2�T(�
�k?��Gr
%ݛ*tg�n�\�}~��&�pv�<�\'������2t�EX0�3g��I\��p��b ��@	�]�k�ˇ2X4`���l��a�i���=iQ��ڷ3=��x/$���}e�G�1V,��䰰��'Jbo��I�ڠ4�� {fY�4��e�lw���|6�=[�8L����Y�gC�K�xL��6����w�㣳S���~�u������d��-۲-��_�ȶl˶l˶�`ʂ!�ߐ��ז淑�� �0�GA���3
��`O���pa���H��϶�=   2�<���]=�Nͼ��G<rQ�(vr	�"9=�M��(�^"�ig#�Y�Lz3 �x�*K��`M6 .Ȗ��)m��`D�m��@�qD��AK=X�$������	�bB^%M�WJ;�
�: �L���H��<xpº<{��Q��~���z�=��8�(K��5eww��� p��ﾒ7o8?~�D��!͚�}�%>�OOd 2��;��.)+2f�������޾�'�d��u��#ka��Pz	_p+�X���u�s���L���T�Z�Cw�	f`TC@�g!�ᐍ��A����������V�	����+�CV��(}#H�D�?@��0�-�c���BOǮ ��M?ݢWM��)H������Oi(or9��������A�� ��p��B�D�@�`��$F�	��=n��K) <��~�\^<��<}����CڌR �_��RF���ߐ b�ʯ/.	������ ���ǆ`zN�����R��R�m��|������i����Wr5$���wD�O�4Gn�t.�A��������RG{AV,23���`4����I	i��5�V�C�x��N��uޡ<��������s�]3"pU�ޗ�Ȫ��;�Zr�ӌ� �ڒ��B��}�2�X���_~)q=�#�O�΍�����N���wZږ+)u>4��_#��H�P,����k�DZ +
$�R�Ϭ�kR�S�{9%�@�-t����HNO��mivV\�@&-˜�h�̴Ǹ�_�%��s]�ƔD9��\�1d� �����ԟ���g:� \#��@��	�>d#���Sk:<u������⾗���9D䘍Y��g큰W��c�u^_\�kf����:����3��l�L-�D%Wd������~@i�}�y��̪i_�u�̘y����f�f���������N��$0B�0��ǽ�IN ai������t�9s}��~i|>>}�����F���Ԙ]�(zmi�� $���*��?DF�-�d4Y��G߀��)4H��~_+�p��%MƠ#�j�ͥ5陳�l���Pۻ���!H���掑�w�I�,���g0��2{������K��P��A�9I�B�$,A��^o�2r�F�<!�#d�h� ����GA��XB�c��:;rx�@N�2��Z���+fA�XZ�%1�y=й�$i��ǟ0x����JD�(j����=� ���o�o�琥�rx�P~�ӿԽ��Ŀ����;��fJ�H)O�a�Ŋ�^S�OO�^�������<H��LP׵f:ɋW��d(��0&�)����]�����D�'�wZ�w�0 ���-K1�A���L��G}�����C�zb-�/ۆ�A��������#sj�m��Y�'yn�S$S��"!̇��|����ei�u�p�,��f�e���h�#ݳ��]��f �L	Q�����}��˔������?�؀�
�CI�yl �	Yi��6�@���o��g�4Y)>7P� �MA��"%�%��̈ߍ`S*�JUv��}`�/7�6�o�Y�2-
'e���,-���6����}��R���,�#@��:?</o�ٵ
'��^��Jd�ҁc%�i�l��C�k{��a�W�����k��ad�bl��:�a@�=���_���y�9�*vuD�e[�e[�e[��˖ ٖmٖmٖHq'R|2T��X
;�q�C��y���0�l_����2�X���f�8�"rw9_9s��ʠ�~tt������� ( t� ��s�^ϗR���B$YZ�h:6��0z�+��#���d��rUk{���^# ���+��7�����w���Z�	�0�^,gl�%��� �.�a�Z�>)8�!��.�Jki�@Z3��_��s,��-M�aj����}�j�[�%�^[�X��&� O2����5eX |��[����
)���^~��_��Ϟ��(nD�.f���g������g?�= ����}P��,#&�����96|����H�P�� Z�:�: �"/d�ͥ�&�{��x2�����4����d� �Q�����MX���-&�ma	��\�����=`v
 ^{o�zD2:C��i� �Jd��l1�}Yą�vQ� ᆜG�LhQ`1Rj=�u���?��
��H�y:�r��7������NhB]J�~�z��-"��+�������w{�/rN�R�G�nHrŉ4u�5[;:�����Z:�)RJ�^K�:F���. ����<i��9�:�S)�^H��c��2}%��x�;�X���V���n��pL���f��z��|	� �\�\�>�������!��%�T�ٖ=�! ܛ[�f4�7y���t�L?Ř�!�QI� �WI����5�Q셑�ɝ]��%�lY��ѱ�k�$d���b5�<����k��grrr첾�..��J��D��ə4:M�PO��X'�ȼ�IlĶB?Q�M�w�����K�&���@(�u�Qӟ&��Dq��Q?�I"�qF�r7�J���8''�%����<:�ܠ��`ܗ�>@G�1i��/�"�LB�Voj?�d>�Qj
~9�l�P"[@�'��(Ơ(}rTc� ���F�������(��?�Γ�݃$C\_�V.��N�IP}6�3'pWC���:M�5� ��3��7�|�w`=��q:�'��})��o�XÞ�L#�Q�����#�,���~=>ޗ�?}Dr�?�������sX˚�:�dZ`,"�ۑ��=��	�ký��+�W�H��	���sȦ����e��fS]cQ�l6�g_}�����s�c����5u��d|/H,Im��t�kOS�;0���� #�r�+<x��c�F�c^!��2�FNNNtO��X�^2[�}uIJ����/�"����y�3�F�S���X�]G���t�/&��$ A�@�$'��~":� e�̔ј�(Ȁ�^so�GRRs����K ��<ҧ����y��	咀'O�'�Jv?A,b}F}�Z��ԏ'̬�j[!��� E6N��#m�X�����39>��d
��p���k$/���QG>�ъ�,���͛7��BFͱ�-����;�27&�ߨ�ݽ�Y���{ +�r4>E(U��罁�&�YfrF @�	��k#+�{���eC:��X�����8r7�Hd�F��z����ؽ"�Z��K9.:�3_��O�ZMHT!��M�"�̐X?'x/r�Ğ�H=v��X8���~i�
.6��@�f��6�y�q�ȅ���R����~�f�l~���L���z�k*���S���HPe�ؽ��g,��}]Y:��ƙ�s5�!)���f��O �j�S���e�$�,K�2K��*�����sS�Z*�2�M����x��r��R3�k�~�A�l[�e[�e[���v1ߖmٖmٖL��&�\��i�~��@���,_�@N��� sT�As 30�mʋ�/�I�Hj�.7s���F3����.�3y{yNSd M8!�cow�,�{ ��QS�i'! Q�$Gf�f���ȎL�L?����ECK2!8��:��{���Q����&S����H��Ј����@��� "P �d��^�2��G��z6K��%躔��dS`X����{��k���0��ve� `ܜ`:�&x,͟��&���L�NoOz^���o m}�'<! z�d��+o./u�Mi5��<mH���/V�]��|+�}�哨�vպ��M�0��:�2�쫛��jEpn��Vq@�0��γBZA���04^�C#[D�����D!�X����	 41FЗ �P���gk�+�zDI� � �S8�
#�,d����`D�3��<���a�
z�d��"F���-��#�~X{�𰯿��駟���W�g3�����DL����G@�|�
5�?���r�2O�����౎�l�q��0�Ϸ:A� ���S�ӕ�h"W:����Hc_|�|g�	�<���GO�ުT���x:� Q:N�N����ˁ�W�O�-���xF�D����a���^�wm�����v��Ӫ�k���4�6�)�����V�Hq��:KᏨtd�$����oQ�&���HRH6s޶�}���Z��8��vFXԗǵ�����Pr��R9˙����G�ۥ����A٦���O,N�T���O��v�8�����3��"���I�=⍍�I�A
�x_w�C�;�� �}�L�D�t���/���[9�T�<=;;��n�d4���}#r�΀�I�wp(��Rf%���gs��0��7��O���̮����v�3�c0�ӧ�1��cY�{��3 ������s�����1�o�9���₠����=m�=�靶1���^��������� hku�r7���x��	�;;}ȵ�|�6L����c�i0�5�j_a��� .��'�����?�ᄀ6Iΰ����e�a��� >��p��l��T>�u>H$���=�:��Ȕc�s���px����|񝎻{�?w䯞|�z�x���Y7�SԵ�F:Ϯޝ�ip|�ȉ� �  ����>5�)��3в��ڝ��y t?�iC4�c�w����C�X���q��˸qNcDB����~O���R� Л�>h_<Gd����&u�'X'�A�����hX�DG������ 3���e0�>��{@�(���%2�Y���AYLm/���;�6�hl5����0|���<���.}iu�x� �� ��o��恬��������A�ttbk1�!V���+	���
�G\eKXkЦ�� غ�3%��a�1�q�[ a�~a?d����=�0�H\������Q�)F���(��
8�w@�2����̒�*xX�aJ�����Fal�ݑy��Y6`1�DV���;H:W���|�9ty���6����.IȆ�q#`p���'���Gw�=J���k&�k��5I�'ù��������x�������\�>��5��y�yo��2V����<�x�	&�.!��̰�pCn+�딖�ʊ�#R"k�y�,�땹όɌ���<���6�,;�ƣ�^qc����ɑb-F��;��7]`�΃4I��eiQH������۲-۲-���-[d[�e[�e[���D��\0�K�z�Iz��M��r 1��� �f�����qJ������&�5� �0@X� 5H�IG�&% ��h��NK�É�9<8���%�'�������7��t�������^����6?
L�a����e������ЀzH���v<�߽�_������2Y�)s����6�, 1�)����@F����;�v�~w/��#�a�
��҃5�L����}uww��2�}ٮ7e�����o�{Bz
��|�un��>����D��<��?'`�$@[I�&�s1=f 0˖U*#�#�y������q�$�6Z��y���F^�����ӧYt2f����:��W���w�P v`���a����ݎ���: ,�  �<E��*�'���� ӓ�n�o�+�e��8�4��̃/8�e��E�����l�dԾ�����$�I�$N�
`���9M E�Z�	��M����Y�#N�RKCJ�A�:��+�t�e�XǢi�C��i��(`�s�Āĥ^{�\������Ϝ3o/.`�v�hMSl�WDtG�p��`?�J(��������к͗���� �O �1��@F� xa����	`�����|��2� !@_Ț����;����G��y��)>�i��57���L��?^P���[y��G������O ��X�g|ThtU����Ϥլ��� ����OD���ǵ(��$�F���#�. =���ɓ�������uF��F���rZ��/�n�H2��+^��q��0ɹ�\�����y`B� =���rrrD��1�XD�2*6N��"	ߍ��?:�{�{��y>#�ٰ��z������k��-����� #��sdrm �@2�O�zA�	�M���K �>|D���7��Jp'�* H�j��~0�zb���G��a\�y�%�צ/�̟F�2P>8�'`�z�(%d�	>�<��jn���\��cy�c�^G�2��g+���ik��>�x�z�����vG�"^��i� |���墚I��ZN�I�Ɛ4{��a����|�@B�H�8d��K����r��3�}`oo�sc�Xe�m��Q��G�A2 >�o�U��}����y=Q&(1?
���,<k�8`��hҵK�����/IW�2��m���n(��G�͇����O�֩��;]x\Y�3_���s�'I�҈�CmC ��^��f���mw8�w�{������n�ѡ��-��>�HWYzy����5���<t�}���8<>������<�$���i����HB$�Vfﾯ�r���:�X�*�����G;ִ>{�{���� az��(-�e����}6_f$��X��#}N+���:����8_.�C�R����?d��H�F�9"&��1<P��W�#�d��1�,��n_ ኽ:tٟ��#�hi�ux�D|���	A���?���Nv��w1�`��}���um��� ��ׁ=�������oxb�9�$HBqbi�vǖq��}��T��{����?C~Tk�y{��@FW@b!4�Б3A��ݗ\,
mK#7J�t5q8��2���8ϐ¸z^E�'B?FfoB)������ɓ�����I`��h�\�j�}�l\�� *��[�0�\_���4���Ї�e>g�7;�d���M�n�2���Z/L`b�l	�mٖmٖ?��%@�e[�e[��S�v"��i��i�� ��Q|�G�!��dDǞ���A|��A*�w7̀�
">�lIi� y�؈	D["*�&�Bst���!��!�լ�)op���j_�>�1^N�>���"�c��A,z�|��[�?d����x���G}I�H��񓇔� ��m���`=�-?MX_D�"|o�H�N��3=��_>{&�W�z���c8��x���6�"�W��7x	>��'����'�w ���є�rNM�@RF� J�ً�N�ކN�nD���)	l�k�=��4��IS�����/��o�����(�l$a�����E`d,����h�LFN��H@�����Ɋ)e�P 5(���_�/����x�A:��i^s�:A�M��IW�/";�2LN&�D��`�����X��7F�罖:�W��  ��T�(�/+�0��l��0��+�B�/�c�\A;÷��>��Ci�����'�
0�"����!�{�y:��!���1����x�{a2ZާŃ��S���R.@>��)�Ѭ8��v����3�r'��鳟L){�����e�1���*��������r&��	�fm�(k��0�4_U���ѡ�I��m��CV��(yUT�7�绛ʾ`�vv��6���"�����?<� 8�d�%��"ˢ�ĎA���@�_�(v]d�0:������@yJ��N
����ƖE	;4����G@f� ��>|��5ځc87�"DO�ǅ�E|<�^�!�I�T$2�V��,A� ہ��1Yi����F�ϧ.Y@�H��O�(��8�D�w>�^n��m�3 � ��<�5�f����ˣ�Ai�=��{A,�lGP��#|�-k�| ��Q�)���~;�د�W\��d�z��Ǹ��yѡ$QD ղZn�rS��c�9�qِZ���E�V��A���d\K���e��n}&8���̳n��\)��~����=�1��2_0��A獞]�b�A��}��`�ᚈ��5��cm�-��"�m�؃$��_��jԅ�w��F�ӣ�f�(��?w����U6ޟ�g*��Y,; �J/��y9!�.62��#_�$�ʜ���?�h�e�Ś���=�獰�� "g�1�$��O(�g>S+���DسO����|��t$/��f�4�w�ʙ��"H��K�g^�sJI�`�A�B
1rf�\�\����7�����9
�r�2Rm^%�e+��s13	P�,zϐ��6wJh��"�ږ2�?tY����*��׳r�t�<8�X�������K�GQ�L^n�.S�p�a�$1�������u��3+(��<�h�^9&��2$
���$.[��JV��?ȌZ�9��"��(pl�ʑ�:�*���!���Q:�r�	n�D	�7��e�؝�/��[z�z����7J)R]߽��������	j����y����e�'�YU�_�ú�
��
G��YCr%	LfT� �K��]��g]�:x��m����V��ؕmٖmٖm��)[d[�e[�e[���R�,C���@��y�J�U`Q{��%T�����!� �̇���#�����؋@ҲE	�� n&q�R&Ĥ�Q��%��?2	�Ш7)��Gx���n�g�r��K�r����u0�Z���5��U�?"x�����������5��݃Cy���<zt��!A3����:I���;����14�?����'�ӟ��t�m����?�_�I���w4��g3g.
 Q��V�z�D8��a]vቲ��?Dݿ}�J��!#CqG$e�Q��k���r��*�$�S	"��DJ��̃������!��A I ���{MRx!suy%��Ԉ�Zݙ���`H	��� J���+�6��`� �a;"(��7b9G���%(?�높�u�h W��Ogc�}��7��er�	=���iOg���L^�9��a���D�yz�hO�5@�4@0t�X�̏��ڗ$E,�y.5d��1��!@�D�"�$�~/2K0o ��g	�� �9�ظFX�>
�k�s 5&�e pD92꼇R�x�,c+rƣ!#��0d.�ѩu	�2k��b��{"I�  Z�����ە���o	��bb��&��l# x<A��NK��`�][]C%��ɪ�7���2N�QvlY��u��,Xn�����f0Mǵa&�Ho��ݞ<~���L����i�n뚋��2Z�� ��,3�����)Cq�E�yn�cA.�zRJg<��,��1�F/�|��.K)b�x��0��J	ۂ uVʲ4�$#FK�Y}ր��1�� �ЯF��8F����!APʑ��~��Ό(/|V@H�d_Aڏ@kQ��yAi�[�ё�z�d@�(E�Z�����t���O��`�Q:��ι�1/����(c�^T��澓k���z�"�1�����;�q�1���/��a\z��I�A���� �5���{H���z>bl{B Л�=���bƨj����Z�h���g�Ŋ}�H���𿑭II��U����L���[�{,R���@��Հt�e�'"�O��9��#�t%��쬈	�C�k�:n�m�]1g�� w�w��u�L�1�9�	�[;��IX�}c'y���'�����3x^A{r]��	��)������+�����rUVcӈ������C�A@df*�yI2��(���e�=2�@0��3��D��Ip���f&�e�H�z����X�� 
�D�)�;���Pך�LGc����j,)�����3��Y�s!��HF��{��2�ٿˏL:%����gda.���A�9o��K�8����n��bc�cu������ ���,���%��Z�kG)N0���?,��n��5��Y��Xe6d��~Vw��y/�^���82�_��IlD�_�����!g�J)����ԛf둵��&�Y�p	
�=������u�	���q1n�@>�����2����T����L��ɶl˶l˶�ɗ-�-۲-۲-?���&�E֮ T  �Ңoq���47�����L �@�H�S$��b��%L�'(�8�`�: ���D�Y���CaY�  ���<�0:��О�I/ �,�(}Hx��2D"�O����N7�u�ot���)eP`����+�r���﫫w4�}��'���ݿ��J	 ��A9��ܿ��K�����I�?Hr��ەZS���&�h�u��+J����� �2*#`�B��L��(8,B�rb�݀����ڙ��M�}��P>&��<=9&�Y8�%wr��g��؁�!��Hy~Ν><���
� !as�F},��R��T�y�L�"C8sӐ~)�AB��a�~e.|�c#�{Q,;��u���u�^��g3%ġ3�/�qz�@�ɮ���@�����r� `3y��#��L�3��"���u�iS` �v��8 �{������H,:�����<#@�XTQोZ]��C�5R�l��'Re��� 0����E>�Pf�A���"B�k#]gj�Y6J�ڋ�_n�� �0�B}���uMj̀�Ȣ�C[OVg���d%ɣ|j�yE(�3�A3L�����}��L��B�v�w!Z�?.���Ϙ���D�7�["U4:%i�u�oJ��#�Ĥ<�l�9D-�N $K��3�xz��>ul���Z�1�e�������i~�xP�����G��\'��=Q'�Ŋ�.�b���J;99�1��<YY�Lvu�\��{7 s��L��Z��v?%�08�����+�~~-y]�9��|V�e�������� ������4|�M�����Ĉ���{�~-�;��G`v.(<�-S��������ڿ�V�­o9�p^N�ʮ�Y���}��P#پ�z�ht߶�.H�FͤxB#(���!��eQ�A��l�7^Z�@�͖�����`��.�����_����p�%=&bf �}~^z)+�Zgu�h$�'�<����:?���-�R��멿����ʒII�3�)��|�ZZV��EX��z���=O�ttD���'B"�&f��z  ����|�t!2��s���z����r���#g^�Bf֙5
�{%V�9�
y5��k�Y]��92>\��f�F!�jm�ڇ�Gx��t_�#�g�{r 2Z���8�2s��(�Ӂg��d���"&Ryln?�x�Tl �����@R�X�o�3�(��zEv�3?�Qx�A6�;�7���������SKO�xb��s&QUr��N���#ߤ�3�.aVݞٸ�����"v�~�QR-�DNV�ef��f���6-���P��ϨM����%<�g����f�l˶l˶���-�-۲-۲-?�R���Y3�f��y���@��
 �F#������m��wdf$$��\�R8Q��� �+id�:]�!�c17�X'���w�߂4UN3jDz�I��LU�N�A*@�A�gE���'|2�3��Jj��a*LR[( XF���4d6��,��ǧ���#�j]�傇q�~�����������_�~E3�f�agH�l.i�
Ck������_�mwz]9=;#	5sZ���|� h���".��$��铣cz9 ��_�oC����ɘ�pD�?|(����\o0�з �"�WS1�3��rL�!H̴�;Z��� @����ج�"���H�Gϳ
$���fĳ1��Y% ������F��Vf$���(چ6œ���#�)|���r���i���}Y�T���U&9����a�� �F�#%hj)#1�
�ei�K�Ѻ�H��+���Z�>:"�u\���= ��"��܋�Z5���^eT��{@j�����93]��i�^OL�j��`�뒲3$:��E���[��U����`)�Ĉ����V�	7H7E&s�f�	"���L�yK MѮ�&Y��>��
��i�X�ɢ¡�f��I���=3} 3�� ��b]�n��� ���Q��a})�o��<H�5|�^������S����̿(�-��x@G�%и�V�8-�u��sJ��X�bןF�Nf�$��2dFT��g	�s#�8����s}_d���$��sh2[T�`&N{?c�ATF.=���k#f�d��3G�|�O��U�K���Ȍ��9�����:�3��擁˲ѯ�0�g&�䲧�����摓�C}q��*�j>�l���1��tB��$��JJ�d����?OJ�0A�-��X�IPlj�\�kQ�,#FA��ݚ5�pP�����ɒ;�	G��s��ڞ-2�z@_���1�*�k���$C�C��U��բ�-�4���e��L�ǜ7���smֆ��#t��LAˊ˙Mjr�=6��1��*;}�6,�g�M�kל���� v�8Ĥ���3����0�w���h[��;?d;���2q ��u�l����FΘ��ґ�fܾ���f����c9�"�<D�/+J��|����1#8^�pWl*g0
�����M�s�4�}�WΓ��XגTL��:�W�37�"%�?�2��e���t�c?���\��N�s�[�@�9ncC���y�[����Hv��Y!X����&��}�2L3+�Z!�L	��ֿ��,�?S8]3q�����oOB��Qzr�����®���{�rّ�T0`��*��[����zd�#b��{G,Q鈒u�|����"T++*b����2�H�3g�VZ_"C҂
>;%i�������e[�e[��^�ȶl˶l˶�`
�c��h4ɈýOz^�ͼ.�E/��A�:��e(�z���d2]��1�K�ECi޽	n��4K�f���m��ݵ���3���^oG���ҁYj���ע��G�ȅ�E��ق�K�8�K�L�v@�vX�A�Ȭ_�\./.��V�-���7wwr2J��`ی�C��~'�v]����?��Z�F`���?�gϾ��W�Z꽍e>�K]��t�9|f�I�����ֺ���<�N���[m�A$�VSH�h��QNh��+g'��W����?��������/�?���[��L�c$��"w��^��oH���%X���F��	i~ƀ�ȉ���;�d���>�$t���ƒQ��Ң<���$t���L�HV ?�u�ђ�#��	5�Q�#�%{>TJ�g��H�?�Z�4�� �܁ �-��oD�.�9��)Ae�)����(����{� [	@@[H�h����0�z>�'>��G`ALY�����` YKh�l���t،��R@�>ձ�8P9	���k ���ݤm�=�������ߔz�����U��TV2�!!Ṓ��;K\�� �cf kJ�Y%��� �R�3?9'�:1Z{UIF���j�%N*�׵�!pRza�~|��R�b�2������ĕ4����s��.��+	TA�޲K\�k#�?jk_z��/)��y��V�'c#ˮۘ0&sh�,����dQ��%�Hf�} $q��_Rb@�� ���՚�Wn�7r�G��L� xWT޿�G��)�,�*�å+rl�����>v�q>����Y1ޏ%pD]eB��Q���ˊyRʺ�$ߦ��ʲ�Ϗ��@W�w�̪�����!3��e���L�����ȯ9 ��'����� �	I��V7�ⷐg��+֝�Yh�؏3�?�H��D ۃb�,*�1i|J�1���8�1�%�ӭS��֢���9��YK��$����[�����Z��#"�K9=�$G�ȵ�2���d`�V��Q���
b� ���b]c�@`�ݺ�\�<z���!�"��~�o��z����t�x��L�6��&�R�W�O�5�C�eV��Uɶ�\��e!�~��B�۩��е��e����"��P������@�}���K�ݯ#o�IB#��i�֐ �\Wε���ܯ���9k�5v���>j1���
oaViE���	�k$�"�\[`���Ԟ,e-Y��5.s2x½E�,��I�Y�_��t���~W�,�<� ��eFʙ�Y�AP�y�.��?'%�y!��A��d}'���I�6��qQ�MU��{�'8�d{�G�����2���bY:���tb�H�������.|&�g�,Vi��N�A�������U8���ev9M�J�������1ʇ&5[k�Qۗ���l˶l˶l˟~� ۲-۲-��^`����Ɍg+d!���N�����`�g��0+��uf0t����A��A0���Ǽ\Y1d��@�L�{>�,�\vvJ;����6�����T'2����kY,'<���^K\�z� ���$����9�x�X����F���� U��t��]�R���w��Hv�=MP���%n&�ڭ�Z�����5���f-�˫;��#��~�4�sF3�j����=z,�ގ#z. b�����^�XK"F�7��Pg\��Ç���������Hj ΁~��L�� ��d8rF��yy�*�V�� �D;.�M�QB�/�#drJg��eF�'1�H،���I�X��Rl��Qҟ4�-L���b� ǆ̇y|���)>b�Lͽ�/^�����޸uS� ����D�g}����n�J�;@�����k�7k���I��b{�Z *R���;YDL#Q� 0�Q���`���)33��9&WTĆV;Ƣ�Ѧ�Z��6�2�>sg-Q2b��F1
V(M��8��xԗ�oB-x��x� q +I�8y��DDvd2Щߔ)B{Û�Cz���Y+�e�G�Ӭt�'.� 0O"|�J�8�� z����Eb����.��sD�4�,��$���"'%%�8`ĺ$�kq�L����Lb�"a��L�˙��b�^C��I؄�U���;*�֨m�Sz����U�f淂)�8Y1�̀��rc�+(=��x�B�x�,w�ԙ[�}�9�Tց��t4�W�u �<�齕:Z�6IS�7�&� �-������~wK��C]�> ���Hg��u��g�` PopNѧc9����R��x���'�⊝��ld�����d��I �o�kU�UV��;��P��i��D�Ɓy�A(��!F2z�����s7�ٜa�Zf�� �9�A�F����@:�c� ��ٕ6R�y��w7����1(����G��u����[���/��b��@���~�K/�P~Ȳ�2��e�R�F�쫢���g��Iȭ�����<��c�pn�)�m2^:�����&�W�2f��B��"�u#��������>GFH�'���I�F�ω��B��{��Ч��[�&�(��Lx����)V�g��i֥�{�|:� ����� Gf���=U�x�o]L���!���m��6٦��,�:���{w2�Z���sy��|�������������9Am��`�������ah<<3�u��/�D$�i�?3�Ϙ����'��!Kq�W�����t�ۑy?.gE�]Sdؐ-�=�c�qǀ���$"K�����ifb��NQi$VY&|�T�
Y����y�����f���#�&�_l����φ6�[zBヲIZX:��ߋ�Y���{pqc��G���1��K�6ZϜ0���:YA��� ~�dv1$o��y
>h��0G&�Y`n��&/g���ܫmߴ (<C"ӻS�}�0��Zõ���(~[�e[�e[�˖ ٖmٖmٖD��L�z�)]=����XT0�(}$�lDq�T�%�V��w7�=l�h̒��z���r?�٪�%��R���H_���(|���J��4٘f��سg_�8����(U�U�S'p5�N	f �ʜ������	�0p�4�X��u��@�}�VnooxG6"��4�� q��_��<���5ypv$�V� d�����Vo�o��:5��O�=����b��������#� �y�z�{r��!��w�������?��`���� D�#���1#[��3��@H�JS=��s���t�w}�������X�ӱ����"��d��(�VV�<#Z�Ny1�* [���
jAG+1�4�}7VF� bW�bg|}9��b?���,����P�ƴ���7Q3�����a1؞AV�D��3�]K^����
G4;q�^���+�����֌��󹌴ǁ��J�����	�!拌�"�m>�L�����)"�K��!I�"�Gә��q��_I͸>p�<��Hmo%�aS�0ɩ4�k	�:M��am�9�Y�ʪ0� �/~ޛ������
�ab�}��/|"�͛% ��� @�����o3�=���_rT���ݹ�V\C4��k�w���ё䵌@"�~�ZJ{�g�i��M�+D�.��0g�A��h�l�k��vhj�v�69�ȹ���1�S�1�"�8�K�M���Ʀ�'HL�D�#�?3 ������K�pD�]'��Ff`�@8�,�e6]���c&^���ȅ	�I�y_��ɠI�M�͟��l��X���h�ׯ^ʵ��$6�D÷�w2�t�z$g���w��E��xm/���]���޲�A�b���� ��~��?�۵��0�o� �z��ݠOp���r=F���5 ��R�����G��������Z����G�����ƚ)#�͸�M y�����~2�Xo��fJ����ȖhDd[`- iP��0�S]��>cmAf
^E&i�5��ai���wr{w�y��4Y_d�\^^�ջ����c�@������:�����\���;8:������n�v��z�ڇ$t<��c��10�H�LF�k�k�5�el�1��=��~�@;�"���r^T9�9��!{��J�ݑ��]K\��1��� B �l�3��~}��8�u9%i����'��D��޾��ɺ�g��۾���"���v#\('X�������іC��������~>��l�r�~ǣ)���ǡ����������\X��C�04���ޏq��	�疷�^���;#yr� �Tc|�* ���~��y���\�wL﵎��(
gs�J�V�%+�Z1g�
3CH�$�k�%��:�/1�Y�.����i����bx���ʧ9o&��9��*1cN���1G\�|���V�:1w�/%�(�f䥼G����:"�<0
'M���V�~�3���ߝ�,�u�t�62?J�g��z�ILrJab�� ����2Ng�`l�����Gb����\���]2|?���0�',�rM�l�ܤ���<Cbϲg������85����սl˶l˶l˟~� ۲-۲-��(��3$F���{x���8�n:[�0C0=7��} 0���8���Ĳ\�w��j`3�0-! �d�/��l[���۝31ޞ������3;��p<�7oY��O� ��ݽFj����ܗ�����Y6��	X�z{�i!�Ì�����G�ɇ��w����x�~�D OFZ��b O?�^��nGp�|�ݷrquIɅT�cП�@�Rn�"�kM�W��q*@q�:H�D���[��: �u�����T�����c <���S����/��k�GC�h����̘�:%X����
�~͋�x���tʿ�M'���R�'�R4�ۨ��<�/�K��e�"�ѥڦ �v�hx�����@���`d8"�M���q�C/ޓ��.�̝�
RS�:��ĄW��X��Or�4` a���T����!UCc��J�������7��Nz���a�?H��W!2�\�7��5���z�;��mT�5������.n����D�|��ɓ'O���o^�B��$�?rn�@��@�}��0��x��d�똧�<BV>ߧ�������;5���1��TYQ�d��깿�;p=\��iW����N1	�U%?U:� 3lϫ�V���<]��u�j׵� �3�̌�74�uF_]#0�@z ��8?70E�J�����
�h�ι��#�?>�O?�T>��#��l��_���L���+F��!I��_1*�����,ࡃ�e �5z&%�{d���n�����tz�(k��C&82��X�J'YF�am���F5�51��>��[o6��m|}����}������c������t�rL�mh��deH��H6�wf�>���ؽx������� �1^�߼���yA�����>d�	�/d�����Y�u}�����ŵ�"�͓W� ������u��\��ջw̪!��ߏ끐����|�?<��ip�8���I����pRB�%�?�"��#3��� ڱ�u>��r?0@.v�hCO`.a=F{OS��Gg\�I�$�UW҃�m
�" �\�u}!8_7�*�c�3o_�!)���#���2��_��^?���<�k���������G�W��8��?�����3d�0SkugX�  8�T ������5<�K�H��. y�˔2O/�)2!Z����ǀ�#���6?�6�x].rC����/�np$�$x/�3-�O��sRsX�����.#��*��U�u�W�p�^���e�$̘A&�`<���Q@V� Bf�f�D�^�4�2f�8�v�ޓl��$�F��>�E�M��o^���g���q}Ef�9'�T��y���FK���J�ɀY��3�O��$A��*7��ґ	X#���#�1|��_!�T �uzx��`����A��L�׭V��vw���t̉Dfe�n]�!'���1�#�jU���)�`���R�qx��aj 	�t��u=��8�g�)���F|�ڮ��1Q�2�V��ͳ���)��9�]�����{
���We[lfY�̑`��J7��	
��'=6���f��%�6����K[uۼ�'@|ֆ#.X_��ߏ�8tuG6h�d���»1�?����:�(�}���ZI߭�a�+I@Jpjߠߒ�t�0�	~��G���O�l<�1<K��@�-۲-۲->eK�l˶l˶l��,'#	��>��Y�5�c�q���h:}p�\�^(��g����aK�=�����KJ���bDid2IFP�c\��t6% ��`GT%����!Z��� ���8(����Nh����<R [�AE�pC����R����n�� � �@�l�hO�w�M��/,��o��f�������~�B���U���j��U��6 \y='���v	�@ӹFc0s�A��Cv������k2��
��F��Ӡt������;� z���5��"k� �>�2�t�-	�*xp8]��;(���mmmF��&i7Ud9u��������":uM3�<�X��:��@���ܔ�Ba�gi&�)��Rj�X��@╋�fF	e��ע��lM���d�Ō�K���m�X����%H+}�QO�{�rf��� ���w ����;��r,_������i��Ҭ���O	Ƽ���/����h�
 ���e���;�1 Qǳ�Jn�-�	�n�ڼ7�Q�� uz�f���C���V��2!�c��+3In6]����}v	�{6[p�i��'k����1��2�|���K�)����!u���}�@�@Ѳ,B��� u�������8@ѹ�m���qrrD�y�k�~�{��`����P�n����j}Cἢa��t��t�����7��o~�+γQ߈�ץ�X/j����{�?�уc��Hש&����	6��<A�Y{I9�V���a^2^�=��,k�d�(����̘3�3|v<��`!��F�H��ވ�F�>���|��g$|A�dL��üAD5|�9gkh�������}����햮�t���͵�?��'%��߽��8X��?�Y75]g6O� �&����D��k����m�e��Fa�D�t{��X�}!c�J�aFMiq���"�າ�|��g�ߣ�X�X�G䐘I����˗>�'�>o"�u/W~�'��m�����ud�v���6�ò��?{�lI���PG��E��RYY�h F��8|�'�ь34�cF���W$f0��tW�JU���{�>�����qnV|Ew�ٍDf�{DĎ-"ܗ�sL�����C�~XC߾}/�'�T�L�x��T��ڼ|��YP���/!C��{Z�����J`�
�9�9HQ�o�Y*WW����}�cü��L���
�3"[rZ�bxg̵;�)fm}C�,�=�VQ.��>�ܱf�KZ���7�PeUvArN�Wc�<�%�>@��Z5{���ZϨB?������ǉS|��	z�]˔��'[�ǈu���|�5 �٠��.�V`��ɗ�2�W@�2(�&�+Z�1�D߻p�L�����2���S������&̴�+�s|%����\�Ԗ7�*~#K���L3�i�� ��%	dSǂ�h�p���bښִ�¶�k[�Z�c�~�g��ԾF��6��p�WD$���:���δe��2�G�
8�Q&f�T5w�����u��L���f��\�߫�+��#f-W�5�uu�Tn�9�qm�D�Ff#� w��Ȁ��^�4���d�j��]W`����?wv�Fb���^������R�6z�;��	Qi�4�^�ʒ+���]�y�0���+'<�k6Xp��
ȕ�H������<(�qMq���$pǐ9���]̑��x�5�ճL�M�ٛ�f����ȣu[�u[�u�]okd��m��m�~���ѱ��ҁ���-Vh������ek�Ǌ�:��ҾM�߬HY5
U �:(X�e rA0��`���ax��̗�M�\.�Fjʪ���ְ��؇���!��.fN��
�	�{]3�V�G���#�'�`�3V���#�&o�dkD+)wI���Y@x_�߿+�o� ��*�Y�:��VovMɠ��A�/l�҂�� ���lP��4��F㩞π ��ֶܼyKn��Z�C����o:�64`4LX��)��?�9+ӯ�����?�D�����]�w-�Pb���7����]	���\���fj�65�8�Mfhl7�8�nf}����w�a��% ��{��)UO@��'{��Y��U��2+���|����Ԃ>��7	�p]fK��hd9#ec���xz�#�������(�ށB�[��3�_:>�8�p���P�S���99:�]GD�-a� �	� �+�O8�!@-�o^cz�;U�K˛ ����C@7�Xl�04P�<�˪p�b� ���F�UEiY+��$�|� 搟����r~{¨t/�sY����hP];T c�{]��*�� �~rt��{Xp�	����cP1ȷ�]��ڒݝ�������w���߸)��tN鿡�1++���@m�����5L����LǗ���\^��B�/�꯽�����thwve>���{y���^�&�'z��˽(�������r���{X���
��A{�iA{a�,�M��l_"ڙ���-�����j�nm�4s�-��\-��{Д���)�avx ��'�x���tZ1+��c���Pgl6d�\/@�����u�6R�W��@��1���R*���J�	����+��,�=����T��rF�rA+�5�kX=�MN���|p �)��5�:�H2�߄��{@yT͟����K��-�!9W"��m��ʦ��;{{�&�q��^��r4b	Y@(. ~bt�@~���[���k*d0P�1��,|�=P�؇�k��3(����ǎ�l�tJ0�fu�uNǈtr�=u^�A޺ςT��}��d<�?#Vl�t���a)�#���aO��̌�[;��v_zr8F�xa�D�xe�� �p�W_��F��<������k��e� (���!�<��``���V��k�9@˸�ް���a�F�Q��b�yB~FMGa�x��m<ț���!_F�(-���,�~�e2N_4���8N��e+A��Q�ӹ_�p�-=F�W.-�*��:{���B%��z�P�X: z����N������J�qX_wǘ�(7T:W�	8(I����il��̙tnv��P�*.�#��b4\)x�����`%Yb�[��[$��?�Bd��"i9r:l�^����Y\ܫ8N�!��p������cn��
����?5̈8b�O��fЇ������{&��f�`D��j��#��H�e��XjO���+wp�;�bu>�D��?�:�����f�����Ȯ�_S�D?�=�z��`/���w�(`h�z�����њb+�K�\;zϝ�K�}Y�u[�u[�ߏ�&@�m��m����~��)t;9>&��=�86�a5dQ�̲��V�:/儠��<[�}ho��,���B��𼎪͹�g��
N�N�,̫ހZ<+AŁ����]��ݑ[���������\&s�6Y5!��6s(��%Œ�(�~�DԖ� �m4�"I�}�q��E�-*�H�A��}װG����AAصܾ}[�kG��	�͍]*VFWS0 ^�m<��Z��9i3gn���˭�=�{��ܺs��0����&���*8���g���}/�Œ�~��˟I�Y!�'����3��'f�`X>��Ϊ�BC��cE�'�* U���!I�� H��` ���C�i���VR�(��UZ��-����H�"3 �c�)x��հ�)��0���>&֑e��w�|)Y��]`K��*4�0 qEmc��0P��cAu9��޻�*U��^�)�
if��jsL �b�0�XWE� `8�H@����iC���71"*���\�z�`�$7�SDp<�<׋���>��ͅ��l�9��@�o�m��{���"��K*�a]�� >͙�������1�f��B׈VuP�������e�	*��nyNȡyWA��x`7�` ��hJ�v�W\p]���Ңn��. И' �gwoO�`n�P=z$�}��ܺ�c;�z�+ڐ�B�ύE���Vg�υm��[�}!?|_~����k�{�ڲ �l��U�$&��綄RE�.p67�'��2�5�20t9[��&�uI��V*3�3�iT%" aSL��u:�9�!�/�>z��D����l�m3k1��}��4%\3c^����{��x��Cy�������� ma$uB�	����\�1_J���Ք�{ �|p��+�1�\����x�=#}P��DV
ܸ-�n��4ȋ"̥Uǜ� ��1�T�1ˍ؀B²:0>s�`h3C�����*(ܨ�K\��YA�"���u�@�q��]y���3l	�_���N4��:�
=q���`ww���>��ӖlIv��
CƊY��8.���{ó3�Q�X��dc�����ʶ��
4��Б�P[L����T���?7͒|uf!��X.�کbی#���a���1ǐ���w�x2U��8+�ͽF�|t*����y��گpdUa�9�|世��Z	�#�!��ɹ���� VJ>�>@l�"��NTS�:����D/J���v�3���0�:��p@ܵ��@�;
�W�*؆��T"@�\&�1�X�������Ĕ��]�E��f �#�[A����B�o�ƑO��������a��,������B���Ò��kn�>�sZY��Cӹ�.��P�����A�
y������|-�
l���w�E��q���}�k�t~*l���/�+5}~�Uu�l�rG�A~���}�~ދ\S|�x�*��W��������5�@�ý�}_w�$p��W?�q���y�JMkZ�[�s�{,�<pʪGB�]?	2	i:�k�+��&�5�j#K�4���'�ރ�]�����U�����[�Um�����\��]�G��m�x8U��:�<@T�J�X�n�n�n��mM��ۺ�ۺ��oE{���v�G��0�I�������t*V.Z���t9e�*��|52�]_��,Tֺ���ְ��pP�����Pƪ���-����̸}�<�{Wn�3�|�P֙>\��s�̪P��!\Z<IE@ 	��+��c����> ���gmأ�:ܩQ-:����@����ܿ}Kv��Y�Y��b{g�v ��;���vy{��U��.��==��L@ ��߾}Wnޢz$�/؂1�5�
W��;i����[���`������ w�����9��ƪ�+�
w��"�&�"��^�#-����m��=x`�܂�^�=9;?�墐>H�8&����ź�Xd@�n|>H��W��
x �H	:$��	�����(�� ��p؅'0������Gdջq�,�,D �3 
¾��o󨄬�ҪΙ���f%Y�8�9�UL���y�h)����� Y�@����  �T^���� s��{��,"A�����=؛�f�".=Z)e�����h��!������g�]��ʅ��oZ�ؤ ��:�q&�����W��B�����	j �>�q��5 �
��CP�1#�"X8[,Y	�9@����1Ɗ#ȒX߃���C��[w�Ƚ�IK��"u�Ǒ�Xw�̥��O�k�-�0���y�Pnߺ!��ݓ�/��x��4�.i�W� Oz$e� 3�K��Vբʆ����:�7���y�� ^��V;l2��t�00�:��c6.п;{$�oݺ-��?����Jn��?D�u�4�6�� k+�e��"�
�lel�CY7��aO��z2�M�rM�5�t,�x�N�������*ItGN�o8�Y��}�!�P5P������7�� �������p�YU�*���0�j���J�$6�4�!ʹ;7������GTZ��߯KX��q��8�d����B��O>��?�L>���u�-�p�Y�r)9�C� ���J�g�Xmu9���!Ǟf�D�G��2Y�U�ͣ�
@Ȕ��B������=0�s˖sfn wg�����e1���rA�l��WE�8��|X���3*2(=
躛a^���|f�d��,4/m��z�"��u�F�0�Á� M- ;��*KIP��[� g���E�3��-�ՂZ3�kn)�K�k8r��\m
�(n���Vhj'\ �贿�9�l������c��p�s�
)CeK�{��B�)��rI�,���]S��=Fg���b�ѽ��b~#����c\��n�"���ba�T+�?j�:���)�5 6�:r��3�D�ah�&�U����������+=����­U A���{u�}�:������
ܧ�T`}S�������f]��A��I���*'���=��"f�����E�k��=��<e`��n�d�S=�������7�$�_k�0�s>� t�}^Ea�e�B̛͚��.��2�+`(��4K0�"��ь���p�J'qL�$�/2;�:f��{b3���q��[)x������ڲK��z�|"��#F��}*����yY�?:+o�e�Va'Y �n�n�mM��ۺ�ۺ��oM�qk_�ޟ6�m�=�Z{��KT)�B�z�"x UdyQ���P@1 T��0�(�f@�:҇w������A��ҭ�^�Ue$
Z�۱t�a����'����la������*�T��j�� t���]������r�;*�G�<�A��\����C����`dw%��x��8X-��7m�q���C|�@Wy����$�*缴\�(N����N ��p���Q��A�m�l�j	@�!h���	Xmk�>,���] ��/���USUk���`/�CڙT�7�eq�c<�������{�Y,����p���+��FӖ mQ�<��U��V;����]��"x��$)r��&S�^�B�{�����$�����$0�JH�kS AI�x�Hea�$����9NT�A�
��M^�Xtt����(,P�^�G�k��U��O\8��F� 16 H�߼Y��|j�
d���6�z��2eVM�}?�����l"\��HW�#L"ڥ�Fǎ ��p�G����ׯ	��� hG�M�ksg��$K��@Y4T�� �a��(��'2�L�Y �1�}���w�\_� s9 )��	eB��-�u0�zl�V�~�C�9l�"���������Z(>:�^�Ѷ؟0N���6��VK���D����=�꫾ܽs�U���װ��+<��s��q�(x �0�1_A�VG%,�"]�1��{:_���P�a\�i�j�V��O�s�I$�q��>��#������ȝ���N��A|�$�df��22,vv$)-w,T��>�rLϯ; !S1 .*n�1C����wߓ8H��B (g<��� ��T�oN� J$d�`N �����
 �'CG����rpM$���>�ҹ�L�/�ʠl�f[�Q����*w�5�]l��c����;8���X=�B>��3�{���X��x�b Y���|ʜ����#{)��p�i�W�Ŭ�~�}�׹�6��c�wo_����Sy���Lu��^����?�8�R�{a+D�:��6��j�s���ט�b�5��p���.y�X뗹��з���kN?�U�N�L��9�f	���Aa�Ό�!��v�Z�-�3��<㺀}�#�s�<1w@~�N���S��f���e��@\�	�2]N�D�[ۑ���4pģ�\�eeaAѦB0�*0{���N�^�̹�cmO�R�Ŝ��:*��ܨ#*;�e!SX���C�ʗ�̌�@���C��qjGN�S�>1�ڈ�a�ZЁl�ܻBQEj�^Zbc��U�\P�"��P��}F��E�� �ɘ�NMؒBק̑S>P�J)g��3��֐�?��:�0�]1���sS��E��*��T�6jS(����p��a��v�پ�s-j�o��8��SU�oA^9Xe���˫#�$iH�Fm�S?��~���*��F�!��|o��}^���Wo�cY$�xA���
��ru~�V;$+de#�K$d\�:sY��*@B�G�w�|nt�Zx,�mv��b����#[3��Vp��A�y:�K�;O�t��W纭ۺ�ۺ��5�n�n�n��-��Ə�1ъ��E5-+�Qe�j3���U:� t��_������c�ӥ�?Z@�$$A`b�s�����C�?��Y���
�nW�ܹ/;ۻ��Y����&,rV�Fm�U �T��,�!����߁�u +�2��1"�`��9lп��A��p�i�֬¤E��]����'/S��ry]қ����߈VO�bխ9�k�;���|n�r` se^�,�D�kmd������u�=����3�,���6805Id�� �EDU�x2a�Ơ�T���y��9�V�+����L���${��B�z�&)�
��B���q��k*v:m����[{ L�̘��в3�I͋�{���[�����(X���3G���{Q�!j�	�#qA� fhu[�@�x0��^�8����& ��/0n�фpd�a��޽��ގ���ئ�ǯ}k��k���udE�YM��D�����ܾ{K������_�,t���`ktC_��u���*�i?�*8YQ�}�mwH( L�℡� G\X�*4}���	6Ř��7���3�ܫ�+�M;=糓S9==�~;o��[>	��7� �f�wf�7��`�����g��;�e_��`���@MRW���9�E�٪���N���XG�#	�0'bk��.&Y��P�w��-����$����ْ�6��H�b)��M��P�-���IZ����l<���X���a�����������b}���r����1������/�x��� �6W�Y"H�Z��\�� �@�f��y	����M�`�֥������;���쉜���'|�*��%�ȫ<��].+6C�3_�%JC�!��-3B_?ϧ�lo!�믵@��G�yD}��~V��M�=�ں�w@�g��*����P��qowO��O�D>�H=�R�H���c�"U6q�x#�����=fӱ�g��޼y#���W��fٱ��;w�ȭ�m"w�F�:<h��m^��=���3y����5#vAP-�%	 q�-�9����H2�+����m�'#�K�|�.�!�Tym�%foaN�(��)KbV���ƪ�
����YA!h��2��9�i����p�qe����EI�*(�]W�sS�E��X�yE�[�s�`��T��ܛm*�4���ǵ��b�z��?�Q�t���?�;�^���7�7�r�=1o�^��a����MY���!�ܻa�����H4�\*w�&]�_,��H�ky#�L�^`y;��"c�z��/�뇭�c]WtM�������ϸ?�-�y~��*��J�h�:���_]AG�T�F8���q�W̠(*�ϡ�/�g�o#�-z����I�U�>��'�S��NE�Ռ�,��{���		��5$:�*+������4�����g���oC�XN��?D��7�����B3����]p8:��@�l��=I����a��e|�kǓ5�g�;a�g�II�c�]�ا�����5��~�9��*�djX6�[�����,���b?����O`	�����>{�㫳�?�?��x)�n�n��;��Ⱥ�ۺ�ۺ�V���-q�8rx�Pnސ��-����#?Z#(YVK�P^��h����Ī+C�M����*>`��r�L�VXV���nԓ{��c��s�O����`�9, p{|r&yHw D<(f`A������K �`�`a�˫�̗���FG��V���S�"����rxpC:�.��UlB�����s�f��� ��W>�����U�[@�&�������K=�'ap1 ����8"�C����өl&C����f����B..���A@��� u�Xp��M��L�N�J�L�4�럩�nHLy?n\������t1����	�Ҋv$�(01`�3�Y.��Q�Zìc Z�y�A~�g�T+aԌ�*(���?5��ZՠZ�-<5�Y���x\�ڻ\0X�@
 mȊ@^L�� ��1s:-�c�\�u�u��<|�P��M*0�77�<����N��9{���5[��f������L�r����?C��1^m����:>$`��9�?�N�u�E�7��Y�_8?��$��#������/w��g���S�[�O��q	�D�������:�g�Tv=p������B���cgK�	VAx=�Z�AM�T�! ����:{�.#�?���H&��ss���2_���&�@2�iT�TDxs]�u��A<`N�㯜��}]��>���&�?�Vl�&4R"�۲�ӗ� ��h,?�yOn�8�[7�Ȱ�xS� �b��8��� ှ�y�6-���!�%	,�0�|&�l>�}~�@Y�H,����=����Җ�K�T����_�y��p΀i�.t�����}��Ã��4���ax��/rrj�Y�C7-�?|�H���k�i�+�^�H8�t���C���AΊ��� KGB�_�U�C���:����Z��3;-S�U�0Η��bH;�ej��k���6s���R�d���$�pgX�a�F��~����>�\��O���W��n��1����|����d$/_�(O�� o_��zt��#�|�<{�\..�dS���B�\(oݑ�����ߡl�۴��Z�����/߲n���P?|����� m�}#�
k%�֦:ְ�"T����[;,�c �/z]�4��&(�@rdX�]>��u���+��q=]a0U1�ī%؈��>p<�xdE���Se�z0f��pK�U�����\�̞���e�\ۻ�6N�̺)�p�uՐ�S$�����fY�_�߾�>�^;��b�CG� ��d��p��e
��������;��Ȉ�e��"�rĈ�̌� �`;�s�):���;��^�ϑ;t�/�gu�G��d(D(��d6���������wnr]Y���ʫ��ieWO�b����*��^'y�G�U�����+����{��]Z��-�@B(�	�4o�a�ƹ�Q����Etދ�� _���sz�5Ք�ڌ��%�K�u��S�"S8nbw��R�jr�V�X�H�d�>���o�T.��n�;���W5o	j�:�F���h�Gc	�	��[��	MY�U yb�Of�5dG����|���?��F�T�ٕյ<���)wq�*���n�.-z_��h����.-�����b9}���{��O�~����KY�u[�u[����&@�m��m���mnn������U�V�H�*T��S�\lf�J�M%0��72Fu�<���$B�����J��.r���ʱ��5��x�d� <��PD�b�"��L^�}'�߽�bs/�>T�_\�r�0J:����@f Z rX��֞��J��ˀ S��&�1��DB cc�Ūl ��X@E[�OkZ3�RH_xT	"��4��~o�s�M�X�G�y�D��t� a# ^�{�yo8`^@�v+����JV����QYh�y��\-�A*۱�U&ղ��"����Ω*XL�ڱT����4-3�I�� ����dz��>ע*` .��i5@jkg[�NNd���������Tz�^� ��xG��@��� @f
à��#V0�!�௓e����Ui�]����氉�@�J�)Υu�{I��B�E:�?��I0ѺJ��Cs�������|��ݿ/������G�� �Ŭtݽ��a�g(o�~e��KU���c��M 7�aV/����`z�� �1Ga0�oc��BHC!��oi�簨� ���;�>�#������@X9^ORu�f΃�^�i�T�s�\��*m�������9� j�f�ѐ&Q`�P3ܸ}���t��{��ŵ�{<�4ݒ��&�
��ePaT�a�pM�:uvr.OxB���riڼ`q�n��j��	ʗ��>���}e�ε�,B�E�Q�c���o�����;͸���: �}��Ya*�� ��Fd�e[B�f�c���_X����1'�ʬ�`�F�$��$�"oc�4��6=B��D�5����2�<�ӓ�rv~$�AOj�+�x,�߿���+gSR} ��N�-�oݓ���,_��H�0�&6r���t�u�~������	�I��(�ߘ� �F3S""�Z�	�:��P�����B��'u����Ht&'�yu�Ŝ��/}�?��"@wP��{ZL��oT������f�ߔG_|)��?�����H*���E����ry>���y�ꅼ{�ZFW�2]P���>��m|~,���9׵y.	:�{k�N�/����uo&�|ʰ����`K]Jc���z|�L!s=�c~���,o޾���/UC̹�T�����.��t4�*���L�4LR=�6G@͡��e��6�
��2�CT�iQf!�!sA w�m1G��j$����:��F+��2��=s������ q�F�؆�! Z�<Jw������p�'[�[r�����k*QY��8���2�;�}��t�DK�$� ��9 O�=2e�MtF�Hr�K䑠p��B�je�*��l�q6�wI�R'#	���}��*���|����@�-������TA>l���cS�E�q���#o*h�vk������-$�P�0/�����*b�v7y��9>����{�Y���%		wʙ��a�,�1������NK����O\h��yf�'�6I�^�B�RsUs@0�����̖�f�
ؖ�4P��pF�y�V��%�µӵ��ne��0tc+�:���B~V�Cݻ���u��
����&�X�x`O��cuX5��@��4��������%(d*GB8�Fc`l���$>%j�Cm͔՗��4q���7Xa�GR��Ĥ!?�<@�ڼ��wԴ���'�k�%(JH�5��A��SN�㜌�2�F��q��yӁ�9m����m6]pkݰ�ɱ�s��Ǻ&���`�˻n�n�n��mM��ۺ�ۺ��?yc5�{8;8
�V�����x`ă+*�	�&1+���W1���N���j�<eE)��]���G�폏n �C#��ES��G2tUe�V�H�����(C�7����j5۴�)X���T����;!���* ~z&1}őU����$Np:4�v c���]�q�Lku��Y��>�e:1����J�*�nw��� �`�3��� YM�<f8���Cs��
�Jx�.����{�O���@���gވ#r �Bq��8�JD�� �C[%�vI�.0�� � � +�Ɠ�̖)	�E8bg%���vR����C�)��-��L@&\'�#R�7��K��C�D�] $\��VB�?�[��<����<c�H�"$��L��3��ayt�0w�ڗ�M�?ȍ[7������Q`�{�״�A�u�@nص��� �jGT ����<�pr; m`��
��T.ڿ��t�]�.��YnY"�ɱ�S�T� '�\��b5p���F��� �Nnv�F�`%j�2tb�ץ�K�>F��LҎ�5�X�SES��F�����oK[��$#g��/:�~h���u��������5	+~63	�
���o���)_��Wrr|*�n��(��©�
��6��#�0�C=�Ϟ��Ǐ�˟���}p_�޽��̩�*	�u�}�[�"ւګ&G	�� A:�>�P�A�{G0UR;łB��fe����������`�����B�-t���\��.?��������N޾y!�HL�������l�͋T����+>'յ�*�u]����D�T������?�T�� �#/�I�j��/��n�׿��\�q�XE���_p}�ˏ9!�ןʮ���u���u`/�X����q��P$�Hu{�ӫ����J���'}]۪ҭr�o��(����ܾ/�}�P��?�g<g���$>@��X����ŏ������׿��o�Ж�ۆ:hKn߸);���w]رG �(���]��12�^��:���[��_ʧ�`����.�F�O>�<��'$OG���m? �r��ͭ]��ș�\M]�{�24L]g
����r)�oJ��*L�O��b]`й4�,�z��'���!��ܩ*l}�b��}J�,�FSyr�ӵ�DX���ޞ���|l�*som�}+��r��^�7o�H^u�!ǿo\�*˜�Z՝C��V��;��\��cu���(<e�˩"'9�~"��^�?�>@>�u�Pr�QJoe%$7�ru���Y^�r*]��{����OՈ�����{��q�,d4^���ӊI
������X���S���7H[(@F�+wf{t���e���<���u�^Ar�V�yӟpS#=�|�`�U�����m�W�!�#�k^`�T2��f(<��5Ԃb�N܎Yp��vw>H��N�IDƞV-�����2t≟�q׫�fc� x�X�Ko#�����9z�*�	.V�"��N�uU7�5�����V2�9��q���
J� ɭ�� ?�c-���u} IҢ���,�˲Z%��檅�X�b� 
ȷ�F��[�'�������<˳��2	:�EZ�I���n<���'��߼�u[�u[�u��hkd��m��m�~�Z�/d41� vOx�j1G���rF0���J��I�(oc���s}ؙL'T. �(*{��`k�GO�e>�}P^T�n���U:F��G���7�xV�������[�9��I��+����N���C�U}w	��v/�(��<k���YI��ϩY��j�h�����_�Zf�9���X�+�_��"���ę���H&WR���nK��tP%� �圡�(
�DV�
yX�0d!٥�B��
	
��;_I���Ջ�?��v�����(�I.\��XH��׿��.������'�� ?}P�H��DW`�ej�S ��>/��-B#8~��K�j�1,t�h@P [I������U��cZy��{��,�:�H
��Ed�ѿA�H�R�I�M����\�&�VfFfUr�DR'f_��,��Ko�b�r4"h����g(`Ԑx8�q�|�d��6���	`�9��e�D���ٜ�h���L)Ё�J�B���D�/�bR����,���^P�:����� `o�KP+��w���)UU���e�J�Ñ1��rU�u�-9j���ōٛĴ��ն���2�����L���<�\�ܑ��ߓѕ��S�e�����t�jk�)3"�<;�7o_���/���{�<Cf�!�;{(-<6R	ʎV��e`�+�Ɔ�B{�ϩ�����Q��0-~�p�_P4ŭ�J(���	��}fs!g5=�¨���:cM�����y�������{�Hە��!�b'ֆ�h��ڌV5 䨀±���NN�/����t=;�������!�s2�od������7yl	�&]0vz�~��� Y�P���3S� r#	����<��Ul�W �@�1�ǃ� �]�n�U1&O�;#��� nwɓ���>l���zMzá|�%���|��Wrxx�斫�G�T o޼��������O���5ggǴ>�nS���ͩ]����Z�R�g!�X�@�,����f�t�j���?~@�I��/��;�e �*AÂ��yQ�����9B�e�p�{�� �M,!��L/ؤ�:`Y���4ƞi6����ք�7����o���F��
I�1O�̅�E��d�5���9�ɱ�)�a�-#�x�5�p����eM�}�n)�L"�����Nm����E�G��&��/��c�aźC��ݙ�wAhkc���d��z�-���L����[���s�����"TYd���2��j`W��%��Ef�[i�/0�����JU�óe&���_,2]'�����|��l��pc�}6J�x2rj#��xb��D bʲ9f^������VVR��;*?�z �2Ȓ�}S#���B�
��(v�D����\�C���N�E!�S,�*���LG�G��T�,��v����F�T1� S~T�B��&I
�lU7�>gc�� ��S;��5�q���ȏ��"�)h�Fj#S�\�z��L?j����x�^�jO������ӿ�ڍ=][c��rW�n.wE볚w�����I��+��.�kU:~&�$lO��N�?_���x������?��'�n�n�n�7mM��ۺ�ۺ��oe��8�"�$G*�B�x��'2lh� �   �@x��C��r5�[5$~�� ��#е�%X
� �`��u��]�wY5���d��F&=��j�U��*Z	��Q �F��;{EE���8x����6�����$�a	�qa� 
���c8�|�Ϡ��bި?�>�g�+Z��~v�����^�yF�坻��=��͢���V	�y���c�X�!	V�ִcY�
9?=�'O����	@x{r~.�>zH�΍��5*�C�8��.h��ED��KV��f�����l*��l-�{yu�
x(@�RZ���Dy�t��q�o�d�Ci�*b��w�\_T�v+��` bQ���6M�˭k��[es��x�@�����r���Y�<U�j��l"MȶW��P���r�\�+��؃�ڼM���酼=zC�,\[dX�u��>����\ކ�%Ǐ�=���� ����{���P�������1	�v�\�X��wd��A�scn0����^g�:b$&*hq�x6�e�CL̓=r��ye��$E/HNF�
��g>�������)G ��������PT c��c��\���Q��{ˌy��秲������x�T������oK��Z0v�Z]T��Ɛ�/��@=s5�����Ǐ��O?�_�����\v���q�1�D
	EY���L�% + �N�3��9������1������L޽yC���k{v~��{����>��`�D�!(a�3�5��rD[�����)[�@��r��TWQ}a������H��	��������2]�,)��Lnm��ѓׯ_˳���o�2�{��a���Vb%H�Ȭpb���z�k�c��Z��b�,	�҅��\'���9.������ �S;x;��r+��ʅ���B���_<�/����F��������w�|+�~�k�F��1υ�NK��e]`통-�`}G4O�
R�[)���a��U��?�w���x~_>��3�u�.Չ�V�s�,u������S~Ω�,���Rk��I67+ ���_�۰��n8�k7�����	VgP9����8i��ڇj�2�UCPDZ�8��M���⺐d1b{M���8*�U�� (���M	Ԓݞ�ֵY��< !9>�iӪ��$4+>���s�C��0�dks?a�X�M����ٸ\�XV�$��������Aځ�J�+>���W����h�Y~�~4y�.4���/>��~�>0���,��ͅ~���ܼuC��}+#�.��z�%}��6���s��۔�݁���4�V�l>Ki�+EO�Je6V����U�{������0���PLq)N���Bڢ��D�ƁX�)>-�+4P�p��)P��.���m�c��j(1;}]��Z4u�_����gx����PS�>]�0^�u��N	QzHm��8�kJ���?ha��p'(A����7@�����:�r`�t�S|�5����~VW��đ��?���nB�����5zz�6�;�OУ���na�W>w{$v�kE,��I����=�����yxq�A����.����~��y[�Ņ�ۺ�ۺ���U[ �n�n��O�P��:P�j:������e�@�8�����.��_te�NYA��w��lX`��p��~(�E*�� @��YI�$]>��a��>x�ŉP������ؾ 3��MSt�~�а�@�=dNՑ8�﨩F'�Y.A�^Y���#YY����ٲP���B8�����b!��	�7dZ���щ��������_�d��a�S���|gI�`2f%&W��j|�'@��l���.b��kV��U}�@:�0s�j����;����������WT\������/l�x�����KO�U���A��(���v����Be%ȱ%H��%=�$7��wbG�0����خ:�+A<B���!St��V՚+����ٳ��� ��a���N�B7��a��2/t�y bk����x�����bS=ԑ�k��b�T�paF���ŕ���@�x<e��T���&����@��@�IF�5?���?���?� ������܃��9x�����=�#@E>����?ߍq���u��ؒ�~�hd�:��vh�@�m��8O ���w� !�d��6vs�ӐaS������)$|�8,V0Op�����!� s�P��pk���}�Pb�� ؈�����Ⱥ ����%�{����%y:�7�7�H�@ 7��/� k��ӖA2�u�*��Wr~vJE	������Ν;����\�S��t<�*���gF��1����e ��c�y��z}y�����kZ�"{ww�k���1) �oߴ�{*��|���<뚎���T��jt����=����PǪ^����s�.�s�9a3#DW���N�S���R\d�|��2�� �G_���x�6r����蓏�:��Iι��ĺ��(�]�)�^�y�����)��zla�UAU�;S)�����τPo�>O�y�1��<�k06�j 8	]�������]�|nR�C�E��.��N�O�[=��뿑��~�۴��{,� Bg�c_6�[\�l��6��Kf�,�C%�I��{�c����o��{~��|�������XY��tx�'}t�$ͫW/��;2�5�Z�
��ȩ���~�DqB�<�ʭۺΐdh^3^.C`t��Y����b����� �^�nG�o���X��1���r�#@*qk��v{;�R�mP�.���Ŋ��-L<���@a��C2
i�'ej�����#p���h��	�5�8���h�w �C�#�E �i��"Mj��5*�	�AX߈����"��a��bD��Zd|����� GWf�6v��������=m�`�S(�:�!���?Cq ��h"�Ou]l����!��}��	�j��Q���P��$3�f���`e$%���|����twrX�2G~X�F.�
hl|9�������|Otn�b��e󥤙���/�`�d�Bƣ��$�u�e�9�؈��V|^wh$�0ri|��ґ�o�R��Ҫ$)|��Vʑkc̫iQ�|��/�J��#vU�'3	�xՇ��S�x��� t��v�N\�Gt�sV!�u���p�cM���ӵ�V�DvS��f���:���<M��Q�}�O��"�M�°Z�����~�����[N������Ⱥ�ۺ�ۺ�^�5�n�n�n����Ɔ��B��@���@�V�,(�{�	r5��
X>�B)��"�)}��QP�(���> #� ~i���� �4[&��OTe�a�p��@�>����w�*�|�)ӊ�@\<���
���R �n�
wJ4�􌜅P���� ��ϭ������eSM��?�E��W�����s�R]2[,̟;�����f݅c�t�f��N-XV����؁C*5���/�����Y. ,r�p��6'��l{r���,���s+��a��� U�Ul�<z��ga#@��v�D@ l'v�9ɏJ2VH®	�}!)e`Y����I ��E�����8l��
�(��'@�:r��" �VPE��'�k��c�0�s�yI�c����`��QJ!�ɔ`	ZUY�-C���P�b���$�������~��|��|��7���[� �A�̧� ���� 9@p�l��0�'r	PM�k�D=��Ax�:N  �E�cD.	���9Aj�[)y ,P��P[VCI J�w�����^C�[�ˡ�\�����\Ƴ	���,��?���޽$� �?~��m�;4X�A9�j��iF/~� 	t/�������Ű��^��dD�����6���� z@�xsor5��Ǯ�as{ ;z�� 9�-ؾ̥�����j�O8gә)�2>LTɪv䒔�d�YU>�O	�b��;�����������[��}�F�={&'GG$- ��{oy<�*�K��|�*s�C�~|�L!\ԑ�o:_R�i'6~bLb,!s�׵�{ڥ��b� ĝN'T��eN�x�;�	�ͧS�K}��Ζ�݀k�\�bI@�;��$XY��_O�|��<1�?}�u��}�DIT׶�w�O��,I�xK�a4q����Po���1+4�ޙ隌<S��n�71ң(-7���u���q5AVo�3�&wv�m�8��L���5�@�O��|��w�7�����7P�hc��z�����r�s������{!��=�/(ꨘ/3�B�|������7M�{�f��e �@���q�8R#��(�ݿ�%����N!a$+}�Ä�G��mM��U�`�Ə��iTU�B{s9D�ړs��IY�:9�.K֍�b#�▩V�T�Ϲg2 ��^����}$��KX�1��`��}LdVT���1	cg�r�H�2�I_P�sC�S��=�u�F��1�A������*��Rb���ER�}�,���(đ4���
k�b�v�����*���}|{{�� ^Р@�h!j9B���'�k7YO���>��k����ŕlnm����E���F��w�_p��tZ��N��X�ű�(�(2�6�^׷���E �a�Wͽ��C.��1�����v�3�,�;r�"m*@F:g���H̚�*(]����k�����6f�M�n�5nS�jS>��r��:9��Y��ɜgM�s>�Yh�棐è�L�cF$4�Q`!�Ŭ���#(W�����	�ڑ�D��{���Y�E��q?�ɏ-�J(�xo�V���2�hƵ�9b���ZI��ާQ4��`���]�����.�o�����N�m��m������	�u[�u[�u��i��h�����k>���9��`���e��l��d1�*��㑳��d2���+p���*o2������-���lS�� ��~�*��	on�đm�Cj���ͷ<�T�����eN���$@j�,1������*�~/*������B�6sZ	���e 3y��X���@�A{I��/��X��*�R�����k�}���H�Á��(7�P��	B�$}�<;=g3��͝-���!�������L��dgs�ծxB͊��&�p�nHch$�#���*U �,,���/���Ȕ(��!���T	0�H0 ��~��X�[���2��U�BT}���A D���(a%� ��+ �ȩ]|����E�פC�-O
�'�{q$I��&x����+�mlp��LkI-�;���yM`7�������_��_�  T��YXH���tu�K�0���n�y�j���
VAImǳ�'��f6�)��K�����LG�P^��W���~ �0�
�O �*(A�E�d%7�3�y���EV*g	�j\=��:�@�k�ߍ�c���c�����o���GO����\��Y�$O�@VW��g1;�z(1B &�~��J�&���<�}�g9��!7`ЃT͟1�D��"we{�k��uܷ�{���ɕ��X��.2/,D[�ją��V4�떦-9�8�g�����,�pO/������~�Z��G��i�jGX��� 5����/~�����!"��t�,����G=�B9�[��Pцم�EE��J���A���e9�������l�d+r�QLp�rYL�l�Ff���7�>::9��q̵���	��: F���s=4��HV��>���P)i�Ϫvm��yX���0%$D��j��
�s����t)qB�R���e�$N��p��Y�.���� -���lO����������o����T����o�m�� �0�r��N��jS�������ޡ����%Xϕ�o��'����Sy��H���1s�&2����;y��ɢ2K@n�*0t�!+�� 䠵,���[Q���=��U�B�)�����Sp����-��*��i����& ۬�b�P��̭��Ÿo@&Wh*�VOK31%�Ol7�1��PҶ�p�J��N����F�FfER��^oS^6cD<
=|2��j���J`��péCZ�C��U�^�Y0f�����(f�j JZ��,��$��"gv�����ޮ���R��}�+�]^\r=��tl�}���լ-�W�/ڛ��^J�������o��ct9�=$��AcFǒ� �r�rj3]r��=G�?�Ҝ��8���U������L���g���f�93�0�����9>A��\^��^���ކD��D9#������w��fF�q:vc-�\ֆA5H,��k+����?UY�J�}���5�Y5��D���N2&��E呟+�;���[il�[pY�G�~��W"玱���s������"���[,rB>��������F�T؉�MD�S+���@���GK�GݧR}36�S]W_��>��y�ǲn�n�n��mM��ۺ�ۺ��?y;�p��D�2����n`�u[��G�� R]�F��i�r����$�`�fc0�L%y��<�|�XK%�ٙ�� ��
�`��Ä�MA�8���L�����X`^I������8����fwR.o@Va���ȌT�)|����s�98g x5���Z
��fC� h���E��?��_�J����Grz~&��J���@n<<B�)2>Ҝ '����ȣ:0���2���*�PY��Vn޹%�����dam�pzT�Nk�R��ޖAH �Ν�MO�=���� P�(0?m\3x�3�YId8YF��lG�KM�=�2$�5µ��t-�a���rʊ�>�BGt�U�gJ滘�#w �K�v�'�Lڜ]<g�-\*�B�U�Vg�R_��*<�T��-��Jl�P�`,PU+�4�x�ji� qae�T�&>g G���Cz����}��@x'2�^�1�� AU�۲��*�� q��+[PB�N�Ĝ�$�EYW��=������� �:�U 2��������QwS6�6��	8��^�y�r<�XE�Pd�0�b.r��+O��u�P����8'���[y�����{��GV���]=�.�-X���YP	�๚'�e���|@:���q�1?P���=_YPseA�EN2�>�I�:*�QO˳k!�h�P8��df.��%?��Q�〵�1P��LѶ��d2�l��r~v"7�9��y����r~rn�ΕZ�#���a��@x0m|���E���)8XS��*�i�BK��D.��������yH���������58�ߖD� Cס:�u{��~�]�.�L�ҵ��e�zz,W�WT�����:����C^���ޒӳcZ�!�ȭ[�	�����5�zlI���3s#�m-L��ş�%��f�t-��W�k�/0wz�.צ�Y^q1�¬�2*?L��kV8 p(a˔Eic�a��q�u�;�Jo4�p[1���9�]D�,(B`)6���_��.3\�H�ܽ�@>�l���GG���o���cGD
�PMF��4�7�x=�����>a>��w�7C�	\�GCS2�tE�2X6]:�D�[K;$�ml����zk:(�0w�^pI�䪿�J�pᚔ�v�0hE�_ʲ� ��H�e�������W����kp��iE����)�d����g��EB}� ?��������,�����S�`l�.P�r�\^Xe�Mˑ��:��?�~�Qd��j��(���Yy��"J�� 9![1����=��i.�9_�~ۢ���*��dԹ��1��͡s���g��|A
��2�k��� P��&c���+6z��>�=�Fi�^��r��h��ǘ�L=�kd��ABw>C�N��`IC�4Z�����B���.,�jw+�p��Wíc�}�Q��N��'��{x(VNϯ�N���g2�ړ���.4F,P�Z�@�E
���ŎEtL��	r{1Ȯ�������*\I#��q��pM��f$H�p����3;Q|73��گ�5؇����k�#�|�N
ȏ�X�y_A�,¿[���G�ӌ�Rn$����Nܧ����>k�:��L�iԙ~�k}�K������__ʺ�ۺ�ۺ�^�5�n�n�n�U�?c�C5Qgr��=V�M�cV�V�g�XҊ(n%:X��ɃAG�k�-`yc�A�J��� %��VkZǘ5@�@�( J�a��hw3��h6��8Ҍ�N���CJ��r4��� ��a�����9�6P�[)�ق���7��a},'''rqn���م�H��W?������>I�����rd��Ak�����z��s}/��\�j�L�P�\x
Vv;�P�ڷ�9��E��\����/���7�-g�G㙴�]H�t���ײ��-}�NuQʳ��9�V�*ԝ�A �P��o�d��`/�%�0d�\ �@F,�S�:-��y�k��N7�e���7g|���P��D�IJ�>� ���]m���A�	Q6!� E��pA�L%ȥǋ�zT� �����9�Zh7�=��iu8V���7s�� @ �u�y���"L�ƅ*���>�"
@��n�n��l�,�ڲ����`@����B676I"g"�m�Y�`�C�C{"��b�I,�aW����Cfv���P����.��Ǐ�ʯ��F��/e2��b�0ȕ�qc_>��z�g�)̑�����(�2
��pKe$T�I��3z� �@�������^�-y��������'\P���wdg�)��)�α6@�^_*W�*w4rP��Xh���� ��ܟ@���bn�^��CM*p���;`e�n[ן�����{+[��ch84U��{��������~�����}������[����m��b��kK��^{Tx�=*V��NAe1]I�}���~1 ,[NBN�B���)������%���O�#��Vn-S��]��Lb��X2�*����
���bgW6tmf^B����)}�oȣ�&7o�����;�����m��7oܒcX����Z����;Z�a{���.3�6�Hn���LG�Ü )��[�n�թ�i���G���uHXx[�:�I�@F�5l}*�a�q�1?���F��	]o�q�X�r!�kt��)�>�g4�˒��yY7��X}�3HT �� �k��=	j!k���\� �S]����h�׫K�f�seK�ۃ���;��g�>��,�u�k�J��KI-�V	����Z��YPi={����$Ee�� H�bkssK�Q_�TaJ��r��h#�Q��[
�b1� pD�3&�W.���#�m6��k��2�6
*���������q�Y��=2�!��P�aA�O���UΈ��@��+���ȫ�ͦ��=���m��>�0m�|&�#|��i@
c����\�
?� �� �+b��̦"���"�eI��v^b����po*���zġ�dT�Y��j]��WH$7��~c�708QMV�v� �q�]=�������������P࡟�@��8��	t���Us��2��I���
�yJ��;;;Tc��9"6�e
(�Ј*�`��-2�t]����H¾	�h��j�3e����D�=k4��2�.��6MA��	k6�?H(�����X�����L��;�}p�9BY��yK���`�
�z4�D@�7��⸫��13�#M|He
����m�!��kvW��.����x���#X�����Ì#kLi:��O�ԡ��k�iN��c"7�d�uDE\���ʽ��}�}�ձ�����ESb�3������c�`�y���l����\ƚ��#��X��z��雳���������A�m��m������	�u[�u[�u�'oۇw���S��%�{t>����pU��J�� "_0�óQ� �(�J�� ��𑟥�-�v �� C@��BCC�x�������4
��w��r0��7���-����g�<;#��Mz. ֪�恲�q߻wO>��y�� h�$��J���!Ũh5�!�w��仸���O���������!Xy@2�NM�1G�����v�
T�C�AkT?F�<���囷ry9&�����LΎ�d2Ӈ�t!��9����}���-�(�ә\�k� �s�h�0�W�2 �$.��h����.���� ��qDp`"h��#�աe*Q;�흡,��G�%��o�����)A�����#7hC"�-i����`*wY�[8˓�t��Uu�� ��=����ٰ��0��*��Y�x0�W�VNuP:��W��0⌟������;+�8����7kr%;�ľر�\�~oU�ZHv���p�e�"�~�H&�Gc&3�gF���"���V�5�L$v �>��DdV�6��.#q��Y7	D�8K����z�[:��?�;�.�o���f�f�Se�J�z��
��$����|��sy�����d�?�	�v&''g��c����fO_���#9�;�R�՛W2�[�	�jS�y��.
L�nSƀ8�py� �>��#�������@����+�g��ງ<��L�pX�^�P����gKY ;
��*�4Ŭ�n��Z:�� Z�W}V����<��`Ӽav2�/}���8��Q�7uiӲ�4�^�����	����:r�����#y�ч����<m�����9!��g��L.t] i'-� ^��@bS׿a�/����:�����۷r~�����j>#87-��䉍͒c����!Bc-]$���E�*Pi/�E~�6PȿX��5���g]��^W�Y�k���V"��L�R�����|��G���:�>�݇�erq����>�>�q��� �~l�X�-��
(3��`	gJ���_�����f1���!�  ��[�yi�iJ5�k�׳ߑ����%�U�{�( y��]YG%8� rh
SjюΗ:�˰��z��UE;L�We��e����_ΰ�I)�����V�2����)���}�������3y�ه�wp���^�;��	�%����H��9̡��ݝ�,:�����ͺ׎ofT�`]����iLj�l�+N0�Kgue������8�\� M�#̡�J{o��-Y^�T��i�{�P���|]��Z ե�n�BF�E�rm-�[?w"�gG���}��Qhy(���<�^�i�ek9�
+������Pl����ᥬ��)82�Px����𠠊�~-(B�� �r�9kGGh.�c*�B�F�u�� ��,,�I��e�����ހ*US�a����F�q�%��4A��.�w�e"���w9��ϑ�k��[X�֛B��/8v����]poe�B)v �j�r=�S�B�Ge�ϐ���T��� �=��G=~
X���L��W��0ذ0nI|��Vق�9��{DZ!���z��fo��c&�=8!��~����}�����~'>?�Reb9/f����pDmV�h��Ⱦ  %Ȋ�7X�7[P�.[(�xw�����*�u>�-Y�y�-�AՉ}V�r����6rגΫ��)I�j�Q���o6�4�򣫯�3@W�kO��3@x~���8�b����o�ڲ�T�a^���U��o�˿ʮ�'+��eP.d۶m۶m���ۖ ٶm۶m۶E�'�1�w'��Y�є�<�z ��*� �0�V�$��$�j=��<%(���^?fE�r9�mx�Z�!��2�����sK��������#�Ԗx�����q��`�؟J:^`L�r�_d��nmq 7*����������1`�͛wru}�� �j�J���i1X�� �^�|%߾z����<5��PąR' �[�0� �(����K� �/�͒J?��*J���zL%�П��ܬ\�@�(�\7�G�nErd��9����A�{@�>�$:x-�� 	 �V�%�>�#O^ڙ>S/�K�'�&-7rf��;��^ �8��m��	���`���Qe�2+�B?'6�&�U���z�*�K��"4����ܕ�63A��@GE7�T8��3@�@?0�����_y��̜϶#5�~���?��b*Ox�[��W�U��1�$��÷��b�f��������������)cc�BZK�P	�����t��������Sy��39���p�s� zL���{/�K�N�6T"���ѓG�}wr,߼x�� K�N�oy#�J`������|�,��@���G������^>������?(U��~�7de2����Ti:��΀���H~��{�*'jZ�-@./�i��q��`z(i��*��o��H���h#��-'PpMG3��즔������/t,�z��c<p4��$ �W?�6*�u��zzo��s�'��7�o��J���Q�R��}}���(PO���pu5�kO޽cv��a�5�	�<��k�k��@���eE�8���s���y��7�iB5v�7H`Nu�:��hz��D�{�R��C��;�&�v���T�ot-Iײ3J��c@�h%����3���l�`�O?���������A���2���B�:�	�~b\��n�F�uV�]�\Λ:���	QU5�Y^�HL���s���$��T�,7YNO"���~r/KiQ���Uc��{�l*}�b�4��²�c�d�68N��{K����'��f#��z�| ��ڏ7S(zTn��y��LW��_"�=�1��շr�������.������0�� 50��Ɋ�����>��Őo$NH��X��%h�Fz���`��H${fS�q^��NA&CG2+�>�9+��oTjxV� [?����J�	)�i�Ըxv��}�9Ř叅� �iUF�;�J����:dw+ ݨ�ѯ���PT�V7�/b]w|�@U$y�S�~���L-�� �@;'طpn����M�B��FY���!��Y�q!��f��B�Qش��̒rC�OUN�K#�n�� ��YH�@I��ʭ1+0��3���,�ܠt}�k�J;����\�i��(\p9a��C��+մ�+��~���Y.Ge�R��b������a��a_9��S���
�fU(�@��W�~�d���&a� �
�*dx��i6���K���/���?�'�D���-�@ �dp� 	��0R���"Z`y�}��?U�fI�y�Iy�`��*NÓ�f���hY"Vx����~E|xdl=x��g-Z0qR2wsH,c�2KB�?
/!�Rx-�?�s��2���� �s7�A>Jp/����l�DG����ssTYd���:7K(A������O��l۶m۶m۟M� ۶m۶m���lG`q�O��xp)
�)]E��J���x8h	�|�����8��{��N��uw����`+�܃��@g|�X�ѫ~F�Y��*�a�@�{�^�U<^��x�HT���4�T@#c!��f�J��\{� ��̎'"�tqq!���#x Ge��pH��:@M� ��	&������A���#i�;��r���!Өt������w�^/\�t��w	�����Rư�X/��#2I�K`OD�����{�@�;����Ih!��S��2�RB?|�G�"� �~l%.��߽� � $���v��!-cr�X ��� h!�¦R` ��I| ���Q]b����k��g$*|���j�BYs�N��kң`�n�B���G�Ђ�(��icU� i]��ۊ�
�7���r�S,����|��\�8�J�r.r^_X���ځ̚/W�~�υ��>�O�K���kyp�t�AaT� ��0��b=7�/s����v`XE Fm��1 b�cyF�<MRf-����Y����������?���'O�<c54H
�.�`���,��.�>U+���5U:X
U�} �7�Zu���s�kJ�
}�n�)�^K:�D�ӱ�-��m9e�_8"?���q�1<b] ptOܓ��>�Z�&��h<��>y�1d�|��\���R�\���C���.7cV:Ӈ�̈́���'��Bh$�Ђk�s���B�`#I��kH>��T6TD�] �1����#-2�������x@5�x4"��̖N��tu��||����[��5k@����Cf�$�on&\��������GٻwH@�ͫ���������ӳ��"�����x�<���ю��ݏ\P}gʄ���A�^`J3Z��	�Ǧ���Z�Wf{�̎�J�R3"ˈ�YZn����W��fwE�ҳ�]��F���e��Ś �����Z@�e�������R�g�g3�#fA��ztwz�w����|$��HƗ7��7_��_�AN޾Ĩ���-�J=?��؏h��1�&TC�a�g簹��]��;��E_��Q�85 ~���5@0�'9�h�����g� �E�����ʧ��V�-�,�� -�2�,no�?c�A�^s���*�.yΖ�
HT�y��ʝSb�qC�s�"K��)-�QN���3�6wT�*.��k���H��T%��b�~_�uƈEP-��ľZ�;2G���/t;�.[��|�X|����v�F�T�_�r���@��.n�����@р�߅�3[�t�x$��'�捯���xj��)�h�:�B��o�|w���X���\&��k��`�\��	��P@���ą>�����Ƨ#A������.�Q}2*��(�ػ^��Qp�y�k<���)��e�O.�/�����p#���9B��N,G��x*`�[��B�Y�X4�E���i	W�j��0?�y��s��^�Ш���C�:�����-|�S~N�a#�O0U6H�^#NYR���
$�N��������w�%m];zo�O����i��O����c]id!-q�}����_�]q��m���FƘ�A��o���Jٶm۶m۶?��%@�m۶m۶�GӺ�C9=9��{������t�JX2,׀,x��P+�O���Kmx�[�f|(Lי\_��tm��$I�!���*?��6w5 �T���|g�#3�2_��G���"M}�EaA%IF%��BgOa���,��&@�, �;����\�~�=��M،<|���4Vi뗅;������{IK&pX��{��dH���	�gS�����>�Ho0�VҤ���zĠy�p	;"z��t��f��^�,�@����`m@�' mTj2/�4�Tx�egg����K@��6;�Hl��Ĉ��j������W��]ɐ��.H���� S;Y���<&��+T�F5F%�O�#���gi���-^i \���MW� )�V��
�"c�J�a�̾�ܦ���.4�n�j ���~��}#���k���A��og}c�XB%*w�*V:~����������&�u*"�z������f�U%��La�q��'Ϟʧ�~ʯgϞ2Oa>�r\�
��q���w�Ͽ���;9�$dŨ��|-��1�\g̉ÃC�1S ���@�=�tI��*�;��@��O~�3�����{���a�3�j����w��o���}C`d�0����gox�1e���x"�xl���G~)V�kI՞)�t�B���y������|��7�콺��l�P���32��< H��/��TT�ĺ^tН�|�(NH�N�o&�:������G}��}��|�_��?�g��5�=8������~�+��@������L'3��f�����ǟ�X��~�s{�1� �WPiV��MA�a�����ە��{��gr��'O�<���F����N޾}�k�ej�FײHg6@Rj���°�qGQS���C�Yf�rX��ţ��� ��l���}���_��W��Ζk��Ǐ��������GE�|5�k�����������!��9J ���O�'��^ȍ�w�1�|4mֈ+ �:�P)1���.��,� �";�c�6���o����φ�ƒk�@T��O���YC�\
g�_!�� �h�D��:�������]��U��c�W=|B���tb�������ٚ��������'O�P��W:�������/>׹|.��{��ĈU����$�L#��{f`�Pf�9�;U9���Z�W�B�I2v��Y��~*�H�����&��2�#�pn ��c�|-Ǜ+��<���\nɄv� yd�T��^V���?3���FT��YX����cV�%�)��z2�:���#j������Ǩ(@���c2�� Ip�h8�@����T.�[:�,�co�g��9��%�T7)�_��V�����9b|{��G&�LֽFF� EQ�W_~%�G���nZX�;ο�ti�} ���`�a1A��yG<�V�$a�������Q�QR!��N��Ƿҹ�4ڧ�Zm�+��w6�e�{�˛ I"o�&1E�J ��H�����X��ӂ���8	-+(�#*E���]�(�B���)��l,2��4�'Tu1[�:��X�0ȯ��=�(����3�o���p�5���
?�?5w�Q�.��TM���������Kq�].?�&���r�:�3d�u�|u/k�r�U�!���1~��32{��3��%z��3�X����#K�r ۶m۶m�mK�l۶m۶mۏ�x���33��������b�-*�����ܝVC�
�@���f� ��\e=ש̰j[�ME1��\@n鈌�*ͤ!7�1�����e>[�g�JFT�Tʔ
̾� �"M^��LU��N[���c�	%�p�,��S���d|0�*�3�� ���w��0�� ��DV,� ~M�f'���|dA4"��uV &PE���1 ��,~�c P�n��7a6H
}}�tS���	�܂��-�p�MN  GV.d�LaH�����@ϭɼ�ãCi������R�4����f�A{'<I��������66���Ҿ�� ����ø @�Y��
�2��Gp1�J�8���T# ̬�Ys��ݗ������4��D@˥���  ��IDAT�1���KaP��3�w�U
�b썑gss3��a��	R��]�zC�Xw�:/�k�n;�]����<��׷��H:o��:>=����J���s9�8ujSV��MoX��~տ=8<�Mf�&����S(-P�j�����_8�ޟ��
����1�������߾�����V>��o���X��hPj!/g?�^�'}�1��"BjA���P��`�O���1w�2�����?�O~�tۉ����_���w2zy%Ȝ��$�Y�!OgL�wP�s��������莌�m� ��[�#�� (A��=ׇ�=g%5�ʯ��\^�&����>�b��b6���=*��������˯e���� G����CM�{y���X��y�,k��$�uMh�����=������{O���k� ~������7_��.d<�d�?�%��[��v�<w����� �������SD����9�3�	֭a�G���S�>/����I����:����dL2s�Vo@�ҷ,���X?88�qPyt}}ey>���e9!ˡؘ��f瑏�c��ܬ��9�J�Ru���*�?'�j{WT�A~Ua.�>e
��0�FYK�:�6��̝r�+�J�4�|�x��>�z��' ��F�J�>�|m螶�5+��!Q��օ��.V�c�C�b�ǜ�5c~k��ڴ�>��+Ϋ=T��`���L��/rX�yn������s�I�1��F6E�0n��qp��H��p�2�	+�������?ޛ]��?����=��l�}�X��P��
��,�@p�^W�,�ns�2˱2����#1�{�����j�$��B'Fv~�R�?שF��������w�bJ���I3�(�H�\W�*X��e���!Ab�k��w݁,w�B�a�E��Y�a�}����2�/̮ꁎ#����T~���h�;�uZ�:ą�����\�06���t{��6�,��{uX�Nf�j6)yLxZ�Q%�� ���
8����@ؠ�!d0OZ�yq��b��1�����W��[�pEn$R��85f���<�̱��n�;�L�����!��y�g����ʈ���~#�t�U��?Rix��Ϊ�U�zt������������� �D�_��J1�,X|�<�|�o�����W^[?J� �y��޲��M�}��n�o�7�4����c^��&-�CK����3�AG�m۶m۶�ϻm	�m۶m۶m�Q�{����?p�>>�}e,��� �� dJ*|VW���n��b��_1 ��Q�jv	z�Ŧ���}�}7�!ˤ�o̖`�v�r@F!녅�n��s�1 A�@�f���f��ig΃Ю�=4�+.��@o}\�ͯ���s<��F����ث�6��;�΄�N� b�դ!R�G$=z�E�Ey�� ��G�9��B�����Ċ��H��Ӣ��`/%�w�pH`.i��_�
��R$z7r=_��
[>��A��z�9�E�j�H]���u�K ƭW���Z"c@=@����\�LJ�#�A�|�d*fA;��ڬ�% h�쒒���@�������2_h����5.JË$+�(��[)z�CePB0~V���
F4o��5�d����^�]��1�,���Z��T8`���Y���C0�|�Cn��%	����ڃb�(l� �F���?�/��\���L���o�8Au{������`�6�
K� ���AO<zB����N۔Ԉ�,@X�(@�t��*v��<���ȋo������}rrʼ��x��݌����{8g]:	!�  LA*�8��	��LY�x�X@�H�<ztO�{��^�\>�|�k�O�Tg��� gs퇹�;��_3�g%��{m�z����|�1Ċnd���z �c����HZFl�;@��h4���S�^P9޿G��OJ�rvyE["��.G�$G��g��!�~.�~%G��.��	B�h4ͮc��8�UV[ъ��$pоE_��+�������U���?��8�����/�z�6(f���bB|���:�����w�q	K<��;@��n�,��B��'|8�}t�P�E�c D1�GH��5 b	����}(�@4��)�ܢ4�D�A X�b�`}G�L����G�5�����V:�.�W�ah�
���Fh�H���Iڂ؂��ٳg$��F��!�A��p؟��N*�Թ��/߽=���	�&�T�S(�: v0��>Xg�<ts�#Xm�)㊢R�xTf�~N")r�ȝ�`� ��j!ض���7��#�Y��'����<��k!�)����
�;p�,,�3Fv���>�Lr3v���u�Q�Ʒ���+2�ES�Ǖ��(|�{@���+��#T����>�Su8L��<��T��s�YY���Ɯ�Ȋ)h��Uc.��p�JP�R�Q܎=q��DH����FN7������L'�x?�9���g�՗��X�/�h��>�u�~��<}��0��r�ȅ�6���ў���������P�b�.� ��1U]�I�&�2!��ϩg��Ƒ����:��%�u�~��e]�P��cu��GR��9F<�rc5�v��^��@N�eK��~�M�
���Ա�1"ճ���6>�����Vŝ�"5*�@H6�RR��q�+�-U8{*�XjJ�BR�,�J�g�,`�*�5cC�[:��3+;��=m�rN|���R�m�"L�����ys���j�\O,R=�^2�ִ�ˏ)h�9���b��m۶m��Ѷȶm۶m۶��7 ��i���7,lv�>D��*�� �)�Obu�e]}
� �' f?X�����<}x��꙲��@R����(��,���	�TP�	d�J+�n��]�'�
�5xC��3T�qϊ�"X�T'AeyTJms�_�Û� �:˝�,)�$4
g3P5�~d9��������Lk�yT����WPg0w 0Щ"�h��[��:�H��]�DD�$�V�J��h�%I��lv	�
�|�9��aA啰K-�E�d�6�#xTLp��
QT�����p�������=�wt(�'Wry6v�()��}z�G�Ƈ�+V���4C5nA���̩X���:V#fs��9O� �X誻�m��{TaX��©��bHo�Jl6�E�@��4���\�M`ՕP�N݃k
�
Z����J`m#�v ���4��pL�b��UH� V�gm�iD����A�. 6u^����?�?�U�z�5�� +o&#i��,hY�7�����C�����
�n���������Y5��Z� ,ֹ~zz!��w/����������Y��9Ԃ��(I6�gK��F(�f����ʫ��2�߳Ŝ��������#�ږ�w�����\n�$����Ia˧�æ]����,�VK��[������Q����}���bx��k�qx���\'�����oetsik����Z}�w�g\�|��]�{��������WǛ͗��	1M��N��Dk�ӣ"����������b���x��x.oߝȻ�M�$�@��Z��	x�a����Ҿ>>��\�@k乔��7u��drc��.�L�bB.��>?��9|��O���L��S)�oR#T 2��4��ˆ*�5�q��Z(������������+�]	��=D~C=�$JH"���� �}�q�l(� ��SF	1��y�I[<��)ڭ��u�p!�4Zr��sD(�!9V	��,�o77�:�#iw�T;�`���q]x`����m���1�e*o�ɣ����7���ZQ@+�7G��Lh9I`��/�
�7�B���?�k@u�^{@u���=���X���+�y`L@�F;-�nP���rq-K* /t\��W05�)jHc���@~`�~��"�1��0�~�dJ0o8�3#�p�5�X#�צ$H�D����N�SE��f{M����{vE���Va���9e��p����dVLY�j�zD�B+0�%���u�y bV�̫��P��36���dde�%�9,�pr��P��7��K�#]�pͱ� �[fK��dO>z���|���.2�R��}��ձh�_�K�������vwv�]�T��\�����R
"�cO���eq�D\��j;�����=�;��j�
�c��9��"��l����z�ql�.PulH5��4�I��ܫ��(���3�J0�����@N{�A�#E,(���+]0K��j-�XR���(�Cz��L����P��8�
����]�+���~�cE,q�!���=�����p�U��O��CJ�{�����W�\]}9,�pbʮ����!�bF��g.'��,\炊�f�O�*����e�h[�f|�����m۶m۶�9�-�m۶m۶m?���_x��ݘՇ���]ؑ ���|~#I#b����F�0�.7rrvA�z��I�7`%@f � PXe�Ͷ/Q�b���,-d�ZK���JP:X�,�����07]|��K���Ocin����?yw*��혂�|���A(���� 	�:ZfO��~��0�~b�_�탘⣮v Y��Ag-ey�*02=����̲$H:F��C��)��Η�c������i�8�"lt1&hQ��x܄z �"��BA�}���y�����<���a��*��|�`�B�႕����+霞������u �?��>Ȯ���\_Ld�R�-H;&� >[��pG��\��pl��_-�f]"F.Y�U�b,2�l����}�p*k�+mD�
��'��[�m�c�2$����m�XԷO@LE	?UӅ��y*a/b�-��r<�Q��-NBZVX\+IIܒ�hL�4 ��#�l�T:�O� )r�"���*������@��\���_~.g�g�]���8���%���5m~R���i�w/���9�Lj�j.	�Gz��Eu�gb���r���~Y6�_~�;�?���(���gj�;���1�"�0d��\L�� ٳ�c9;��R�0���w�/:���F��/�
ף���s9?=�?}�\ǳ/o_�ɤ���B-l�:������pLAi3|�Pצ>C�E�[U�>|��ؠ�Hs��oݶ�;ڪ5��O���|�՗����ߩp@�@�2����z=oO��weW�	��Z�������_H�ky<��!��t2g�@��5�M`9�L��LU��R&3}�����;��_�Z�u�m=f�No-�7W������==�ղ��H� 4���9�Md�!I�q8dFG��r�59�O����y��__�ljv|h��<�_��_�?��?ș�n��}�澂��]K��Z�)lm҅�d��[�f����}��辮7�4ZA����Ejj?��ձ
�2}�`�B��s!��Ƙ紗[���׿o�B{�r9�qcb ��9���b̮�)my
��Ú1_Ϲf�ϰf��)6n-�*�^��|��}M�~:����/Tz �����$����<&P_,I� aݤ�{3��߿�����_��ピ��sc��1�"$��u5׵k�r��ޭ��ud&)l�tϠz�J
1��Z��Xi9�qT��$��Ț��؅���7�unDX�0>�g���1���g�u��%��)(��W� �S�|������:ֈ	Z�|�͠lL�X :���,ZA�뤑	>m� ~�n/3m���ĕ}�\`��ޏ�1
��6�W��]��B��i�	0DqT�u�)�䠒��(��10c�S 8k/|H���s��!�~Ĺ�
T�/�VU��2�����اG�,�+9>>�^�+��=~.������<�H�k�d�3Ժ�Юm9�t�*�ݒ{������fAZ�7�oѡ�@�=����z_t0��3P�?�a��d���y	���3,*X�r�/R�?PXS��D�zp��^˭*,��m�~9�N��kK&77�i$,'@���AZ��1��x�s��b�wP�r/�x==�
U<J�u< ��z�ǵZq�3�D\�LEn�E[}SYV���Zx�J�\�c�����������'��[�N��ʏ��j�jg�F*�8�3�j���Ү~��A��W��.��uR:F���9�]��>�5H?ߑ~A���a�}3�Y�(���59~Û��^Wf�lV�/_,g�m۶m۶mmK�l۶m۶mۏ�!������gS��ãRo�!P�0^�{�zN�v��}��8��˛��r~~I��Ԓ~̰"H��Z/]Ш�3��6�xwy��+	$L�SZDD��@E��`F�q�e�5c}�G�3,gP��J} e}���|��7�B�7�T�jD�� EJ��L,������@�qB�T@�����Q6�8?lT�P�@FT��H��5<�H�����wlPPyާi��a
_� X�̳��6�LY���W_�۷o	l?�w������ɱ�@N���h�������1+�U����Ya�/X�,ׅ|��7r1:���| O�`w��*�Ws���5M҈���eG���5�b&22(^ �E�����%��;���}]%-�	��d�J*Y�����k��R��� ;�ǔ$ �J `yv���ԪAs��Z��2���}���2S2#�6k3M76ϐ�0�����$ ��xd#s�A�S��j����@r������.�Z���VS�����#�(��j(�B����X��&�&���]k��[�Ā2��)2p#H?k���8]QQ�������K�ͦ2H��_.R�[1��T���\����|*�Ō�8�q1F�TU�h�O�4� (P��㇖}��A��1��O~�sy��}��o?��~�;��H���(��Y�V�~�/ �*�����Kl�)�1<�	���E�7�r������K9>y�kӔ�A���s]\���7�F@�V�}����eZ�����H�J��h3��k��6uP�����w/���$\B�����..lm����b��Z��F�{�� @���s�� =3��lV.ϦR�a���E�Pr��M����<!�y�cc6[�G27ߡ�������h�s��IZ:�u킊*�l���Oa��J��=�6�t�0y߅M[FAJ+�׮R>���]%��b�8�2w�w�<����>�+�<1��<��v���Ǿ�k%#U z��[�ǳ�D�-a�7ƣ�� j����N�ǰᵓ=]�Bƣ)����C�I��>��˰J�:��*�����=��,�����YsY�D��*���ʳ�e y��j9#��>������e��6��Ȉ#�2�0k'����(*nC�9낊B��l����DALu�ܠr�gP��Y������{鲥E�,,��5�]�3
,�"��+���
�,_��%���1C,��sW9	(; a������-���N�J��L�!����*����_yα��A�S�s}u#o���]�1V@�.t��u�$� ��2Ȭ�<�[tN�V,4��}xp��zO&��lntL���{1��(p/SRyB*��eʱF1}
�N����¸��5���{7恙U]�' �V��0wp��}܃Vn���P�Pys�����ȢiV��Aq\�}�'r[��G��G$FHc�{�W�w�~��,���b7&$ȰG�9�����?��2����6*�	[}��-ɫTξ�w3s%ֿ�~��W�@���ۑ���۴yO�	82'��G��-|���k�K ��b�C��+1-V� q*���
�E۶m۶m���նȶm۶m۶����
��U��1� k�r,�s �l��r$��<�K�����?X�@X.W�)-��D��$0`_6�����6|�2!I����`<���;0�=��r3����5���X���?�B5���w߽�*�t���Y5�j7����ق�WT} ������U��~|p_:�����M�<T�SU��$��= �����������6^ �a��sD?�F
`?�X��6��f�oC����W��R�0츙�1x�>��-H�o��Z������^��]�t,�AK�={*�]Z�\�����J��Z����H|f�X��H��u_X\�fz�77x����ΐ���' 8`��J�i� ��&��h��	R�jW_��oah�G�t�X@F� ��E{�¼��];��J��we��=��L�
�(k^���v�YXki��r�k/�Jp\3��˴έ��p<�kh%-V��tT �6rk��ۂjD� T�h�x�p���-*1h#�ci�ѳ��m%����8E��H:ƚ	�(C��TG7�K�����F��1DɆ��z��j�Ũ�NY9���p��X�{�-�6X�`�9��
�;zLk�P�I��hc+��Rň�f�u����iޯRƠ���tzÿ�x��q�j���0�d��+=����
���c`
��ye9 ���+��u���Ⱦ��H������t~u)���o��� -jnm�*c-)/2Yl��KC9�L��kG�X�f� צ
fT��`��Y.����:�0M&�+�sS������zJu�o`,v&�)�|���Z��a�����H��a���Ri��I9Bz"�Ѻd���������pg���M�)�նJ�,F�m��1ՂX���X����~���ׅ��}�~���"k��IXN��[0�3�1���ɴ6�� ഩ 
��_a< PY9 ��� ��ґ%�k:�Y���E4��|s3���1�1̑��5�P�
,�:��^��f�Y0/f���� �{�]��2������S7�2�Li��7��e���m�y�r+� 0����*�A�����Mʵ�l�ڢ
�ܫ����6��:[�vbP���֚�&�E�vp}��.�>�eAn���7ԙ�zqN�g�Cʼ�*a$K�wQ�hD�����w�]帘��mMiD�=H~�f�f >�!rg�)�u��s͞��?��bdRn9 �1dVf���#��%�U�D{-o]�/�t��v��1�y,�>�$�����:�? �c��GG�2�ձ�0,�g�o�vF�ȨY��XKuM�}H�j��\�z�フcO�*�
�u,�@o���+�A�5�,�G1Hv��������3S^�p�AU�\a�-X�@�1O-�����t���SgEa��=S5�=�-�|�HT9n
����O7�6�$�� Av��:*��ys�TR���YD�w������&+2�R|��	sG�k����Þ�:~�?
sw�!	E���֟�:�����]��z�J������>󎕗�H�Y&�_	M,_��[�.Lx��w�������^�k����R�۽�m۶m۶m.mK�l۶m۶mۏ�u[=Y��x���*�B	�ȼ}�2b�% rT���	��QɻX��{U*��X�a�4�����C�+�r�
�K}����2 U �F�2ݰ��h�	�T�m��\��k�򫥼y���(-�5PUU�ڀP�� fe	�?T}`�k���;��5I�b����j|~>e���
���>�X:�i�~!#e����ѵ��#J<삀�3�u<���
�D���Z�/�	Z�K �,H`#ш#ٿ�K������J��H���1{؛$D�a%b�*�%���S4s~zE���y�{{ڧ����|�ͷrvv����0�<����Y?�2X�WUȬ��c=V�*�Y�!3DSU�뗌2���Tٸ1��T�*	:�X�g�_��A��u���JY�ԃ�)�|��R%�޸����!�cU��z	�}m3o���?<�c�Pj:�����ְ �r�G˞UgY���@F�����k��un�fK�������a�~��"ژ48��^��l!������)��Hwۖ� xFa�����8�ш�$5u�	Xe�'8?���,!���1U*�j��r*ѹ���;ؑݝ=]N�ރ��/$�L�Rdk^���vv���L�N��.;;;\��	�x��- �8�;.��7y�K���C6�¸E��
��8v����PE�M��A�À}���?�#�%�C=�2az�ҟ�]�����\?g�}�5pI	~^���=��}���d�#�^�aA�@&������ s4�{g��a��^���_�� A�޻��6�m�Uu��³S�a[��څFp:�+�g��	@]]�7�F:�����3P�,��J�����Ø��l�wXosp��@�@�j�༌�/K�;���P� *��+'�[�j�'s��V����l���9;>c%}����:ᚆ�w��;�=��7I�P�Lo���xj�M���Ln.��Du?:�L-\v{������MB*�@Z`$�Y���R�)fa�� (R`���:c�9-��N�e5�Qr���H굻R��U���^�,��j+�o��{ �L�1�5��޷ ?�4g�)�3��R����op���K˯�֦���U��f�4��k�5c�y~Uu=���=��j-�=���v�8�����w��i���wD>n����>�3��n��x�.���$q�
ʤ�
���w]��3r` �@J��}��hM�5Ub=�%�54`��KL���}z�����[i7�:�r���x�0o�ny��{`�It|�_�\�{ʃ�q�&��`'��z��EA�S�w��^�q�����6d�r��Z����2c>����gߩC�:)�̪H�������;*�A}ҹT��d.	Q����o�X�VRvm��\��n^�%V�w%(�fƩF�
I��e}�a*N9bR��<�����G�����:��T ��aH^&T➤�S��_3�S�3e��.q���QҔ�~fS�Sq'�uo0ܥ*������ٶm۶m۶���%@�m۶m۶�GՖ����M�f��6,x�gvG^P}�\Tz΢@_�y a�i��f{N���������\�i��@����n�:<>Ͳr�^Oߧ�������9��-��G��+J���OAR�[>&p��S ۩d�]��Z�~v��h�/^�|Y�ٜ v��g+��R��U�B�dU쉼~m���ޔ��F�Y�]��A� ,`Y�N�
@"a����@4������8R���S[>M%P��_F������H��vn曅��{#����@@}:]H�� _��4%x(Ƅ����W���5n����^N ���<&����+�I��wLb d�B3�*O� FV���}��'��_�T�A�9U��.��B� 	F���ɪ*�e���: 	�(����J�h��,�`���B�}� �},V)�
�b&�
x�#]��+I�/�(}Z�����	���|5_�T����\�ǒ`7���$�-�0�p�)mل�c�X	2|���e��0_�6��j�^9F`6 �r>�9���oX_e.��Ȩ������-z Ęc�13|���s�e�L=���z��[��L���� ���F=}�@{H���J�b"���� <@HX�x�F�/�w�o�K�PkTX�Zx<ƕ�l���H� �q#����Dd�:7�7bD,֛�6~�&�F�p.b=	"	d�`�'�F�{f�D$�`��Ǉa���݋���[��>���u��I���k5�(`��yqI{2�y0X��EȘ�;�<�s櫹���H��I�~�P��,=�mPl5Fځ$������
(C�8��a��֙���Ζ2�̘QTJO.��i���u�c��@�˚�~���Ąq�G�}�GeΊ��>��bfm�Xo`��e��{��*��R���	��KMj�����T� �yk��־��@�y.̗23�X׀A�1K��� .="�\�0�&�������+�����ܾ���.S�}X/�.a�6I���0���^@g^M�`��q�:R
 1�z�v�lA���c!�ިm�`Gi}滰i��	Lc,FL�. �9竆�w����Ƀ�V~܊A0>�ā�?�+A���i"��a���8E�1HnT��z<#�z`��Ɓ�f��G}���4���N���zqP��;�����*�I`c\��rD�o\NUM
O0y	A~���ٙ�I�����p�;XgQk�"���_`��5�t`�}�xR��N��"��LJ��ߗã���:?;���������O����85kB���Ǐ���B���j<$�8HN���	\�K�y!f���)jp�b?����
$giUF�1�K�ȶB1�7�rƢ��
6�WVk��a�߻�?lzo���(��QJʔ{�G�AO�	�C��0D��Y�/L��2=���F(s*��6�����
9���!��d�m���M��9�BP��^�kI�.	���޲�c�ig�œ��V�����,+�����QR��}��q�>��P��>������8��d��)�������۶m۶m���жȶm۶m۶�(�Bx��[@�9*�����
�TZQ"�V� JQ�`�-%=�Q��a�o�}�L��6 F6)zªj��Y�2'�p�V;� v��|�� ]��aS�{�����G�bx6_�j�d��U�FZ�/�/ U�1X��Y�l�`K�#k\U��7��ʓ�����5���x�&�#hxA�
�55�P} dӧFTV�a����b��j�獞��JS�& r��P�U�f�p*p�ͰC�) �tmT��i�j�e��O�ۓn�E۫����Ïޓ�b&��-KV �±�9[T��Ah� 찖y��T��  �형H����c9<ܗ?|�y���?22����9�0b�J�*�v� T7���		�U�&$����g��V�\�yE
�(c5<_o��a�!�6��z�?`��{�m��Z� �*�ླ
k���k@�g%��j�$y��PUĞw�%�Ϸ�����/�P~�	���j$��XN������r���<�f�)	*��w����s������W'����==9�bǴ��g
/gG�L�Ām������,�pP-Tj�WIU��'T4������6HF��f���38���Fn�Y��~6%�b��
��й���P��lj
���`4 (,#g#N�a>��v�|퓞ܻw��@�j0��,��3�va��"��)�NףK�� |���b�c)�"��92W��s��k��	�a���	�"��*�+�9��ܲrp� ��b^�����ȗ_���7o��.��Ti�\+�J�4���ɹ^@��s�awbJ�W��vc��a�}XYV����#�$Z�� �$jԹ!˹�} @�T�0�;^�Pe�]i�� �5T��N���T��J�%��D{5��G��9U"�_��׵y��]��,�]cf�0$;�h"TI�ԫ�aq*$�@�=S�NMP)����o��\56$���jB����@�;C��<�`꘬V6Qm�Y>
�n,�3*����zD3�yv�F��3�j�s����S �q/=��?���P���o�2��T��>��̓>,6��&�ʩ��Y�����ڊ !���s����s��X�����	"y�s�ǉ������Ì̙p
=�	X�V�|����ϧ��1�H*c^�Qѿ_Yequ7�"+��������8F#lA�c��7��֑5�\��Ү1�����zM���~nFbj�;`w��S��B��VT>K��( �������ڬ�i�Y��
rs��#�v̹~��s��������1HeC�z@H5�ی��N����>���!\B�Ak��x���u��ߡ�ōS*J��S�x�������4;<f�xH�
�A뫝��6�ql�ߜs��Z$ϫ��� |Yo9�t/a�TI)��z���O�"�]���2!���q��cc���8;����r�s�W���*"�}�\2��NAR���^d�{.�c����5��oGt���y �Ἲ��u�o/wL�Yj}����H��Kw.��`�n�Ǽ�h�s���5�ڶm۶m�Kk[d۶m۶m���[;n�ja�"���C>��D��^d`�|:#�P��Y؈�2�uêo�I��C�Y�j���=���
���pA�@���z<���)�~m� U�yzH�.���D���3Z|@�Ѳ�r*��:�_ f  �!U��2���C`*>��|G� ���(A�UwAi�����=�#�B��t��Q3�̸����fM�`v��ʆ�[8��i�|ڝ6�TH|x�#�L%���I~��f#�^(�������\�]��Ź$1�N�`��g���Wr~y#��)��ʔ�A2Lԗ�Y9��_��G�YΗ��=}Jв9@E~����"3����2.�u�9�z�g!-��!8��k�Q�g�-��A��Xp�����������=V'�ߐl�[3Y `y�e��l�,VYo$��8i�M�d 	> 6����b����D�n����N^�CJ��"�2�ӓ3�<��wo�2�|��Y=�<?]�N@,��*�=��*d6�p�`<��k�w@�@�׫�H��Z�n:�pn���� �
��_�HfSد�e2�H�5d�XX��*gB�e �?���C*H�G��z�c�5������i���Z�(�rS�\�|y K�v����L���A��F�a#��w|�|��'�]���}�3}|�b�x1ruN���8�
^�����$�p�>��U�;c�s�9A�UN.&�Z0����8qθ���5�|�8�� @�<}$'�oXM�е9%�ײ��e�?���9��[w7N�ês�[x����kGG�v���x��;7X#�J�GG�!��jt)߼x����YM��X�(��In�����n�6Ii
Ԭ��WM7��L�q�Ƞ;�V�C�l8�uD�/S�ᬖ�&FT�x�ۉĞU*Ӗѷ�	kI3*͂:��v��1��m/��F>3p����$"�'�Q�:�d��w�[�.C�7�w���P)�o���=�P��P�
��#���ISS��k��o��䝼}��s��,t�L�3ڞ���^�����	�/�n��<Js�h\�>_2̨�̭�2
���J����(t���en�4�ȁ�"uVu: �`�2X�;!́�����DχVc,l�&8`߾��?'�q'���L�%Ȁu����B�[q�0˃�µ\�2*�6��δ;��Ya�P �Bg)&w�Ұ�\5(��g�4k,(��5����5��Z���OۼԩB��0+���T��aqK�����F��K��p�+3S��$��T�G
�Q�Cf��S�PB=�s��[��Z�Nrp8�A ���$��9�3d�h?��6ֆ��r{d%�H���_�-j�2͘�"Ft�F��2ү�~�[^���q���P��"��0���[J�,�%S�8����LZk���*-�Od��i�w�\�IX�G?�{�b������G�WA�����`J?u��ZY9e�tܛ0Ĕ�Pc���&E�+$��C}���S| �$��!�Ĵ���3,�����8	�+E*.������E�$(�5UP@�P\i���go۶m۶m�_N� ۶m۶m����r?+=}������
���yB�}g�"x�L>T�@�.T������T��l��l�76��vU k(%/j�j f��)-P��C�z4T|��ż����k�
���
Y�7�`��b=_R}�<������§C���4��#�gz.���~�v�S [�~3�72H�A[�g�)�P"K[Fl����81��dFK!���p�󼺼�|1��U�E�u�Z��T�q-��;����J��a��r��� ϑߑ7��J�?^.�f m/�@�=:�w�2_�d1�
���;�6��t��U������^,�mx,-��]�t:::��~B�� M�sl�
u�I�_)��㪚G�׹�hMw�۴8�M�bn�~�k\=d��9w 	�����µ���ت�^y���<��ބ�	�,o����OB�y�c<�:W
� k  �M�`1Z�a�]�i{���J#��9���N�r�����PQ�3$ճ���.�Mh9'5i�s�5��3s ����P����aT�g�p���Y�eg �Ǐ�T����Z��d�3���X�O����ȁ�8? �~Pg��;-�1�d����,�o[D˚���[f�-�c�{�DD�2�b��S�"�M��`����H>��C����J��PڍAT���̮-]�H���C����9�K��tA2o���X��b���6��Jp�� � ���!X���� �� %1^�y���9o�ۨd��H~�������)����LV����Q�tr||@� ],�e�������ɐUޏ�:~��O���=�z��W��im���tW�mS_s|�"@��/��u|�[��g��˯���[��#�K���Y:����
�����)�Ic�g��F�z����[]�}��d��XF�E��P˅��= �	_��Vyna	��e_���m-�i[h!�/��z��F��t-Ag���� [�� )۷��&�H����ѣ��ӟ|��m�c|@�N�gj��D �H|����~C����it��
��2�AĜ���2��C��!l˴������`Y���/�-�K�*#_k��/Y��cC�2��{�8��&�:ӊ.�C}����������ZX�:6`Wf���V���Kn39PuW~Ob�"D�F�q��3�J����(�.@ܲ�,�p$-���YI��W?����/,Q� i���%t����9�K�l5��s�Y_sO �
�(fJ���z-��+�fXEv��|����OX���w��(p�R��$�q/W)�Ж�\���1Oօ#�M��59�<7�7�����=%mQS�����>��=����^���e.�׫���:�)��@ ?l=����,��$si�I�T��ު��>0t6Q�)khQX��CD���}7����^ǟ�|����qR���ܽ��`M�#"(�Й��C�$��|-����s���@_�N���M���l�
�夑����י�UBU
����)%�S��T=w;d]3�����;�u3����9P��'A�B5���Awb��ymh���d˶m۶m۶�y�-�m۶m۶m�����r|1.z{���\]x��C-�_��X־���RX������mN�uT�/��
�Z�������lഘ��4�}P2��2P1���B�a��
?���ֈ��>p��2 q��9A��i���M1� ����UCpN,t|e^� �P-�,�U�������7��6�U>Z��Ϝ�z���o]��|��-zAЬ.���9`���T��X5%ؘ�=>��MGx������j��8@T"�>�4�����Gd��UUi���j"ޞ/o޾�4_��GG��$ч�F�!}�\���9�P��8��Ӕv��}�� ƹ$x�Y�{��J���!pU���~��{�#3� B�}��l���s�<^��$K��KXUZZFBH]e
 ����
 �,��VT�X ��|��E�IN˞傕��#���+��%�h:� }E���y3w�3�|4 � ?`��s��Jpz��n6H2�{���_�����P����҆#	�A;"�Ԙ���~G��������޿����_��d� ? ~.�K�0��`������ux��#��������ϙ�BB"˨Z��ۺ�|�����cn�9��>}*'���_��js�����7;�5��aa�Km�1Ꜿ������?���C'��� � �*$�ևR�՚���qL�kPL�����-��
��F��@��'�r�ޡ<zp$�V�9<�����sU@M��"\ �Ǻ�\^�cfR톊�B纇s�E@S�u����0I��6A�L?����G�˃H `@G�i"�?�Ō��)"��������q9�_������j��lf;��T�t�ܗk�g�1
�����o_����AZ�5 �Y�D����OB�MAoW�������X^��N<�=y*�?���b��+/޼�x�k4�Z$z��D@��y2P���G')H쫫���KYN���}��1��Fܶ�k]�`�;?�5�jm������c�����)��!�n�(��I��4�<*�x0�,'�$؈����b�^���s%��V�J� �⊠1���ގ^�Ta�@��+�uU����|ʲ�`u�BcqS�a�PϹ�����B�c�}6x]��>��f�7�m�|��y3յ*S���>S�PA	��¸��L&c��=�ʦ�?��?~$������a�+��v� ��s~�\ؐD���� R�[{A�Nb����~��l�7�íu��]U^��$d�z��ܑHZ��И3�H���H�8�����r�����(*����Q�C��pM�{��$K�&�}�J�:}��s�.��$0hv����#�����v͈ոثGէuw�J�p��Ȫ3�^.���a�XO�S������;����9����DY�@Pd)�`�ٌ$��0�n�Ҹ�U�~��*���{tTD�*np]mlCC~��	?���V�q[\#��
�vMhU
����o�?��Ь�^K�ļ�?�/If����<��~n5��O���]
�|���0�D�������V\XKu,ռ���sO
�jcUـ��id}	��O����S��dv�����54jB��}j�.C&�f���N=�e`��\KX,�0��3�%էq��e~G���6P���\P�Y���=2F����Gljɔ1���{���8h���8�.���.���n��J~4$_\��^��'�/�L����_Yuޡ�`:��?����;��o}���?ZO���o}�[������u�gI�p��Q�p����'ȃ���������f���r���dV�d(� ͪ�
pj�D��j,09T����n��F#���h��>�Sː�@��g8Qw@�#�U��@�ZDi�Y[K置6
z�o�s7�7�]��)��% �X߬��F��W6=����~�5d�%?7 >�v�! 
��d<��  :*�[����4|p�Ox�7�; ��j��Z�,��&�%��A��n���	f��	��?���-��g_s ��:L�=C�R0账�ze ���o/�ɣ�� 6���ˢ�>�T^������<��T��q��ۋf�8��e�1A����f�4�yh�#�p�@�VU�����uR�" 7�׍d�,h�7��rZ ��7�jk@^��J��>3��4mda�Q�� ��� �T%a�<�O>�H�={&G''$ dhQr�*!�-��G%�tx$����{��ଡ଼_�����2O<�pF�u3�I3VvC�����ɟp}���rz����� �kw�n!D�v-��c�૵=}D����T��6p1Þ
>PP��J�!;�j��	���?����s�sשJ � �*~�6 c;���*|�.��Oju��g��UHC`��s
̫��N ��g>�q�%�PF5���vdM)c?g�&C����xz�ߛ��o�؏����ҕ]E$��A��Z��Y���8��v)���|�[���$CV[%,��W��׼��VG��+�I�a�x�743z2{�|�V��B��p<�ֈk@}� Z}���Ih_� y���<�油�swq'��;y{�R���y��9����.��0X;��H���Ə��H�m�\�ӵ�h(r���];��d�ך#�y��|���<���K�}5����g�Pp͝q����T��t�Gk��h���ri��-T��	�����g?���ǲ\,���ڟ�5�}��+X? �A��� s>r��D�SUJ뺐u���zA��[���{�<��K��}��{�o��:y�D���N��ч{̕�����������(w�Ԝ��vĶP��{��2bR�8R@^��i�X�}B`�&���Sx���t!�j�Y�F:; `��-6O����Έ�	^��P��H�����iv�s�Ǡ쬷�.�
�M��>ȰϹ*YPm��@�
!^�[��2�s�\����mUB�&b���ֺ�z^�Z'b�q���Ɓ���@��?�����/-W��l�`�T"��}���Qm���ű�������Z"n�.�f0fB=�N�Y��u�G�)m4�^����@�'�8�c;�]LF�*���T����qw�u=n4���z��޺��1���ڊ~�k�Z3ǫ����������X���NRCVUn0�VWQ�ݖ��Z�h��l� �0��k?���M�		�Tw�m�S�"�]%�ak�3����o�ь��F$x�n 8�ͫ�-�ޣ����;�hL)�IۨnJm���):5}���o}�[����n=ҷ���o}��o�C������x4�-W�b&�I� Z<�!�[��+Y-f��w#C�k��^_���%+�aoT���   K�B����7�����86�=X��ߦmh!��v�z!��S��z<: x/vT�w^Ψ�D5&*�X��տu�@,$��<���.-	�3!��LѰ�D@M+���4���jeS��cW+�_iU>��3��د�D�-�hQ9��d��5 �I��))]Q�@5&��=m_������bfE�Ң���F�`|�ݝ,�s�몔��?���c�=�<<�|�)	������ۻ��|Ԧ�1���l�����������_�g�X�͒88$�=�'c9<~ _|�~�auj�Y]�@t�'*)�z�� Q��-��[)`����	U� 튦P�q�/5��A/��)��s�Qk��瑟��xg�UY�m5p^����ݡ"����x��C�m�;�}�����OH@`\��Ud� ����*��4��{�(e4��mme2�� ����j�A�.J��]�`�?��'Ġ x���l�[�VG���Z�iea�S�@�sN������ϥ~p,L���<��e�/����)����Z��pB�Ǧ����X Y�=~#�� �������M�F�-�e�v=��%���/?�c��kD��TZ���\�{Ik���񃦂�j��E��y�zAP,uC��\�r)�5��|���r0���#��-���?���Cߧ��b!�M������|��=@�J-�p�T|XnwP����}5]e�S��_
����=~ތ���% 2/ ��FZ��ȏ��p�IDF�m5%���f�%Ѩ�����`m�.e��v��_�Ϙ�q8�f�����_IAU��O�;�Y3��6t h�k�p\r?fr�����-!(6 $�bo���<��n��s���{���1��e\�k���D1�L�8�&"���E�RG���H��1B�%��P�\���o���~�3*+~��k1@��<_�5�b�
��H����o�%��*PϬ`�UWf��,d\�9�g${]���3.�5�k"��~�����:��?��s_u��*L�K�bG��Ȗs���q�~�(. Q�=��P"����u"Y��:ͯ�S�O���b����j���#( �kWk*=��:�P�I%?�����1
eO�����d\W�$cc_A�)��\�@�`��)�B�3b9j#A�Z����x���p/��X��h�شj�� ��Z��~}BX�x8K�G�S$E����Pc	~��Ԧ�f��{��	ҩ>�=2�Vf�5�+䄠�$�c:��w��X�x*b˕P�	L�-FTr�E'�i�
�GjE X@p�v��Z�T`�kkH��I�Ꝡ���x���~�mA��D�*�.'
���z2eY�5E<�=�h�I�DH�)CH
���ɱ���[�'�;_�3ЪY8�q�}I;�Б-�էq[�>� i�y�(a#f-՚�?;ܛ�fK��Z�$HY���Mv+�*�ml��<��ءz'����2o����@P�=��P�������/ξ�{��ַ���{�z�o}�[��������Ͽ�w��=;:=�\-���	w~xtt��ɣ������lv��o gx�l���էշ�VF�\�z�|T���MV�������h�X��h�z�E�����y�q)Ô�¦J�-�=� � ,�.� �QV�Di����f8�=����-�`��><G�';ڇ�Yg��X��nW:���Ш��T�}5�"��j�# M���׃0�t�Ҥ�.�ᲅf+J� R�4$92"��jѦU "iv�bn�-q鐀�4���������M��{�?��?��?)_�R�v<?m  q~��pTPg�;I�S�l�U���<�>��d�$ȋ�����\^��1��A�l�V�Jݝ G
��C�
Tm�gjY�bi$�� �r�{�GT/K5�>Zd���ȏ�~�s�������	�O8���C#1��cE��KT$cL�̇�<zt*O�>�gϞ�b i��P���T��y0H� ���;Y,oe4Ѱj�(s�9s�j�Ձ� �G~�MFj��m]�����[*���P��	 , u�M�� �g7����ky��V�TG6< ����|�~����Z��#��h�����O8oJ��/~F����VٛSQ�z׸�~ ���r�_c�h'�4 Ѿ����2��3�����&��)�+?��7�>H(ߑ�(j)V���}�S���ne�į6RE)��ֳi��L�z��G��?�g�\�nfru~.��+�yd�T�j�`!�HUe�?+����,�ЗP��F�1o)��֤���u����l�P�Me2�@L��E@T��5�B��T��k��v���bv��՜k)*�g���5�s��U�ߜ����^NU�2_n䛯��_}C�û�Z6���u�(���z�Pd��y-C�?ί~���qN�!��)���RV�B�ÜU�P�=y$��$'.��e{s㏱����|�}5�\���#$��Li �n�}l��\�:[g�dJ ݱ���3!G$d�h�*�a�5���3�r��Ҝ��
BGilU��;3�\3x0va9���!�ݟ��������^1����!m�@dɀ�օ�����mL!����׋�4����9�k��x�>���<|�����ٸR��^��H�yJ�h�*^'T P�fa�+z�en
�ws�kdkxx�Y�u����*����@U=��G��|���$�T�b;^���?V�8ռ^�]�ݯ�ڋ"	�D6���G9�6��t�4[�py�t*T�1�=���ĺF3�$�w����Ǽ��T-���b�W8�&S��u4�G��#�n@8���b�M5��1�凢���R��Y�4H�s~�RU`*�a�S4� �+�Y�� �H��}+��"q29�yA���F������9Cb�CX��@+5�E%�����2�}�V������T��v�~1��h�l�k�m�������.����\X���8l7���$�$�t�ܿ&�3ڰ�a��=����Ѿs�z2�Qط�U�i�<
NLǬ��14�����ַ���o��n=ҷ���o}�N��d|��/��������s��urt|8��� �Q�*�,I�(�����0�e���񆕍�K����Wk= � .W(Po� ��!� i@" P�����zۅ
���I4&0���z�6�T�d�jm"}�>�V��ߋmM��ةu��w�	�9!�û�V�i>���w|"�z(0��X,�*�%������4�ǀ~�{�d�]s� ,�5��0; ��T��^�,>�VT�c_c�w'f)��$���a6�l6�\_����ʐO>�PF��`��0��7od�\Jլ�p�m#4٩��V���D��Va �6Wk�tI淓�(� ��>}Jk����s��A�0�/�g���2�*v?��c�l�<ҟ+�ҏ�-@ z��;5�1g������|���!
�(��6ZM����|�5���V��P�V_�j����QwA���bd���`@ld� @%9Í�{�7<��棌��o���i����m�)�d,���`e��+��O��~n�d4$����+�c�8����dz4efK�g]�E���ٽ�^��7/_ȋ��a�����V9M ��V��Rs<�����6e�*� ��耠����~X���a+�:+���I�b<c�`a����L�<y�Ks+~��_���F�-��*Y1�rMA%0�x�������,��`��w(*ѱ��;>g~���t��]�K�����XL���)3�4����6A��>�Bf�]�>�p�j�lq��'��;�hf��� �9���$`D����P6��т�777$�p��< 9D���?#���O'D�@2<y�\>z�\V�k?��2�}+�W#�X�	�y6:~m�xE����ܯ���;�e:�Z�����5m�����H�~�O�}ǃ1�� �����FnJ���!At�{&C58���-f$�%d�\�\���CyxzDB��O������	��ȣ���4���nX	.�@�~݋���sc�G��ÑYd�y���`�����ŕ�|���!��p�5���	ֶgI��� ���z�"����V�m��G~?�����\�����S΍��S�����h�����23b�j���3y����.���J6���Ï��@���Ǭ�3,0�@ƀ��������>�7�$u���s���B	\=�&l�0Y� �8�97F�!�#�ub�N#��`ե98�0�t=u�ω�Zg"D�3��o�5'���q��Ñ����į��FQ���Д*����"�,Oi�u�VR��I`� �5:�i�Y��L��k<��1v0���V	�$�y������[�4�nV|]H��]�������g�d(�X�?�c}�I�:u,�6h����!����6�f�e;P����,�R��u6kz�� �����ɲ@�ڈ;U$W���w���U�3E��ӂ\�1��N d�q�jC�IS4a��_p���N�l4�K�f�P���-ڍ����o��Q���ua��F�����J`E4-3e�}�����o���.����(0Z�"-����k{ [v��]�Dg���}}ǲ�}6�P�ҙ��Z�5O�UZ�������ַ���o��� }�[��ַ�D+�f>��כ����z���õ`9���.�"&ṗ_�@� *q�#T�Ne�=�/�|�b��b��pE��@��S�a�q��@iB��yc�⨢EP)�܏PE�J�T��DujJ��Z���o?@�x��~̢
$Lx(W4�fxx�D	6�hYn��=�����TX�j5C�*Iq<8f�^����3m�@�-�QA"T,4��kV5:��1 �)6����a�G`BbZO�f�v� �P��5��Պ�M���@�q+�Ն��~��TiŇ�|��L�{�˕�X.iC�>ß�,J:Je�?w�������wv����Z�/�`�̃O>�D���9����a'��y��������q�:Uǘ�k}�*؞�V�j��2��9l��]g	��j� ���6+諢��'q���`z ����n@��j��F���<��|������/��?�� ��~A`y�<�8���F)�U�p��~����_ ��掞�س�P�� R�o2ɣӇr0�Ҏj�Z��Ņ�z�B�g7����&ȵ�PתQd�>ș��KY,�z���Z� ���o%,��p�j�'��X��PJ�Q�J����R��.��/~E�J���
~���N�+?���󰭇���u����Dպ\�>/i�����k��hDEN�_S���*#n����h�p���k�t4f�@UX`=�Nؼ�sx��}Vm
���sM�$���-5`0�u1�l��҃#U������2�����;[�$3����6�7Wrr|*�G�~���l������c� kQ�Z���S?V?����yQ����~��s�_7����8r:�4�Ծġ�8�v�8&�oX;WK?>�\+��k���| ŕ�Q�5��������c�K���.d����������P��#l���l~�����͚d�����6W�ZѼ�2�k���LfN��>6Y ^��1�H��n�b��9C�R���E�| ח���ף�l���sk�w|z�0x�"@|F�@�mT���y�H*ڱ�Wjm�p��[� G~���8}��-��z��n�8��@@1����}�����~����$@��Ԃ�kP[���il�:����J� &��P�l�w15 �(�s�l4ԝ�+HwX��u�� �Kٗ ��$ QR�5 �3�KZ[�4+�3Ul�7 �E��������~�f�v�q��~��t#' �@�$���)�Z��k��~37"mk��C8����9f�?`��pB��:�$.O1���Z�z�+�`�O���ծOS�&Ղ��+���o���q����RⰪw�0X-��,�p��T�E+9������u}�{6W���%%1���r7��;_����_��%	ߢ#wj�py�*K�N0�2k@�`L�$C�n�p<�z�cBf�Aqޮ�oINN�������غ@śhVQ{׼���������fΩ=X A�X�V��0�����#�^�����h�ʅ721?z�6F,�!��#�-���Ѡ�;2����	����X�@�D;�om̉�J�`��������HbU�� )���[��ַ�}�ZO���o}�[߾�����|������$���&��������
���	�U`��� 4�b^��	����k�$=��$����@�>��V����*M[V��Ч&}k�Uk�s����a��*.ha� ����;(i��
RC�Yў��l���@H+@[�E��@n�v�)�P�Q0UX]μ�6X�6j�7�=�&Jw�B�r�Aڀ"�>�a.��B�C?H�fqo�Y�*B��c��ϊ�v)�@i�O���ʻA�YNla��Jf#L@� �����G<ToD֬�o�׿������c9>>�4=��'��Ϥ�nh��k�\�)0�Ff���k?�5�����;�Y���Դ%3#��䳏$$R��WruyE@������	!��M���V��}i5D���G�d������]���@W
�� w�}]+�5T .�Ճ$���|a� 0� n����� ��ٙ��]�Çj����ky��%�/�FR[*_�^`hl-�Y	�U�~9Qq߶Ś��r�����0Z��(,y0�:�x�>���|.g��^|�U^��X���	%L�0wR���ŋon�
J��Yʽ��1+Z�@	B2�i�v��j}u#WW�r~~&7����y��+�� 2=xh�Q1s|X9LK������)�SװFZ�\4D\����ٺd �?dr|�v}l��-�'T�@�
�H]i�8�|Sme�($��~�9�~��}	��_��W~����2�}99���0�-���f���~K�&�S�!�jigvqq!�_}#[��������/֘�[Υ�ε�6NJv�~,/�O>�8:??'q
BY+�77�Y�y�Ƞ�x�T1�e-kۥ?�BF���0!��(\SEG�X��4,��e`q+ۨ���F!���n~�ީz��E
�jx��WB�y�����3�a,�����f���l�ˁLxNy	�t>Ӟv]~�C����9���m� Z&i��NE˨4^-�x	�Sf��H�~B��#�0dvL��6�>
���9��6B��DX��@Ain�^+�Rm���l!77������BOv@`����e?�.���i�����7_}%`#���������לS�X�
�1*��
y�5�����,^��Z�5 � S�U��2�(R�&���2Қk�/*!Z{և�vLM��5(��;�����1����F����j�S�-�~ږ�$�6b�N%�OdcG_��=�X�D����(���v��C-��3B?"�
���U�/fM,Q�����ᠳ9K��b���Q[�v� ę�D5�=��QAT���3�N�����`�a�Q2H[݄��ʬ����.�xO�op�E�Mhh�?�{ �d%��^�������U��{ؘ9U�bߓX	�ȏI���uG�H�v����f/�9�(�>���y��Ǧ����;�2��������G\[`��c��q��z-术�;��k��}$j�ś4{���º�<�g�*�
_��X����s�W�e��5�����\Ŗ�O;�e?��q��η��F�	���!~����C��_9�U�*�Gk1�D��ǽ��Vk����o}�[߾��'@�ַ���oߙ�:��MԶŏ�����8nyҮG
� ���@�`�A�2'G'�pw/�����P���$ �F��ʐZ�ʰ�+xk�LOq�, ����I���4׌�H<Ċtj�������"Z	�0��|Ui�5lF"����$;oq�왋@ɆT�@�A���ӱeۆ�z�y�@ؠB4X@7���J%��k�f���݂ɝǹ)S .���z� F%�������d$���؆ߧ<H����hHlE��5�E�?���V~�Y�}2���}�*Zرdq*���o�C�\�jFU��Qo����?䯅���c�"�����Zf�{��T�?"O�<e�3,z���d1_�S��f�%ID8�iEeL�?!)R6�j_$t��Ҫ6R�
v#�a(�m�jrgʏ���sITEav<���p�ʏ����1�Hw)�F+#�5V�n����ȏ�{y����8���Ғ���r���U� q�����J���㠪`(� yv�F�� �a� <�$<�����7lNp.�=����usu����_|��$��˝c��ȵ�^���	ǠS�
ZY�T���	���h�X���Q٘o#?O	�:Ζ~[�"��_@� Ć����W$4�K�u�X�(������3 ������@�ͪ$��ǅ���z�
sx��D%�0�;��ĵ_C|��U����y;�������G�چ�H
|[T�'
����f�����T/Ϥ�}~u}'3��m��?�YLeS�^��[I6 �2��c T;_}���~�B���sY��.��d�k(���Q�v4�&�r/���1xw7�����~��С<~��k6��jY��j��V����Z ��.�e�3�� �4�^! =��A!G@�R��]�_�T^\����L����h ��P��V�,�:�c kr-�����@ǜX�]kP���Я�X��؂׻���j��F0�FV��������W�%F�[E8�l�4��^Ú���J\�X��EIG᳔�J��K�#�y}pJ�n������Ϗ��飭,�k?�W\'\[�f��$͡���Z�*�:��o_�z�u��P�!'U��W�Zk�a��ʿoE�	�P����uX[2��"q�C|[SI��?�?�@�.��,��j�G�SB��p�Y`X�
�I�K����� �����Ԫ�k+^�D%x����T��}���#��!�����@�؅�z�t�@ a���Pԥ��,��qm��0�x���V`:-j���Iܖ9-�q �Z\��կ��G|&�c�PH���kd �$���2I;�>�48Mh��S���*(��.��
���p���Z�i�ck���}T��
���{'lg��C(AV��4�r����6p��v�Xq���x�k0T�o��;�[�����T���	�xG~��u;(�Or�H���A�**���8�����o�/Ծ�gT���?�����g�k&|cBg���O���J#^����T0f��)�D�OWA�k�#)l�j#gUm�饎ef����ꎝq��p�SR�.^�݋%i�eID�;E��mK-���8�4�Zm��^�=t�3@�χ���6���o}�[߾߭'@�ַ���oߙ���a��_��B��ߦqޢ�]�� x��@�����[98>���#���@%������%�" 1�7�2�\&��H<�*H��u_�&6(:���H#: ���������Z��B�&-�G���
F�9����X��|�Z��%�Z�!TU=�a%B�՞%k�~ۨ�FaQ�u[�
T����JG~G$y A�1��-�/k�jo��� {J�EVӸ�(B�'���w�R]m�w <4w<&��Z��}Z�P��`�@�հAR@��Z@ �
�o^]�dx ϟ?�S=Ǔ�ߓ4ȗ_|E�*Na���&�%����qΪ�w�\[��3�����)����5A�G�3LU��
o���+�f��vیYA�1 ܟ�&&�	�>�r���	�\�f,��&�@��?<���	�]I���a��^�y�>�_�fa�aK�<X���9[����-e��|�_�=��ق�E�&����
����l�#�vW,���c�cJ��K��7�����h�o�,�x`97$�ߖ������_�R��?��L�%�A�����	�
`�����M��;�̑[?��O��^��v����;��/��kiS�w�ɿ��s���y> ��%AX�M�H>�q�x�=I��,($\�h�������!�����-�c�AWA��ğC�&@�l-MQ����T?���/t�V鏱�5���qư��}�s0�5���b��W��}?�e��2_�9���ne�)�ٳ����PNN34~������C�V�����o|��6���9<$1�s�}X���X�R�/�Y V��B�>��;?G�I��J�ѓ�d����|N���ܯ͓����g�.����[����G~۱f����l	\��,�z�Q5A2kAb�	�\cY���T�cߛ&!)el��VU��|+؁���]]����`*~��?n]�.n��^dC�zUY��C �~b������'�㘋�U�"T�`= IB�_�"���\�¾��l�H�S��q����N"�r�c��kБ?���d�c�H@.�__�}�d:�E?B	�u�PK)�]?ߡ�˳���p\�"Z_aMz��K���o���k���8��|8���ƨx����+��L�˹*@��.�xH��8M�9�t�A��c�O�#p W����~�4<]�������j ��ZG⺉~gд}!�R�t�ͪ��s4j�*SH
����+�+UK�2�����T�l"�(OHN���?�)/�u�E �O�fh��+��+�N`�Ҍ|��;��؟�F�:�`	WG~��u"�k�|��*z$l���%YGບsK��¡�>Gm�J�P��P��0Vp�@:dS� =l;���-/��#�V`"���T�P�bjl��5_fJZeJ��&�8�NIZ��Ü���R����Ѭ3�3�
j��TOd��T{��%��@�30=�0r�+��ه̆�� �&i��,-��Hw���-��z��!�C���?�ׅ`e)-�i0L����K����3 ��3Um����cf�`?y����l2[-���Z� ���T:�</�5��^%����U�P�r)X�� �Ͽ��9!ZLa�U\!��k���HA5�8�X�1��(qM�;т��T�^W[���+���V���ь$��8R6��9_�(��:#@�ud�)�H��~Ͷr��L-���C����ҷ���o}�~�� �[��ַ�}gڢ��E�'������{�!��$C�'=��C�>��K��O��&@��)Y�Ƒ���X]	�p<ӊł�i�Ӫ��ڪˤP �E;k-�o,�a64&�G�_��2R�FYw�#x,	Z;��|G�`�$| �-ps<�C`��v���,�l  �ʊ,����o�)�9�)+�V�eU��D�,
�~8���t�f{?�P}G����`1���
�c�Q$f�0��ʬ(����ZC��#ân���QF�lօP�R{	����f�Ѳr��O>��?�_}���wf$�Vr||@ e���Ś �5K�x@`�ys.q���@@
 �O?V��k� �X�]���D�v��Q�=�g����vc���Zu�Z���q��(�V}l*��O��T���.TQ$�0"4�ԑ���-cY̗K�b��?��$78�#�*�RG4D�@\*6[�lv���2!�SUf͂co�}s_Ԣm�?��&�W��+����U��c6�śQu���sK���'���
���D��p��P1��Q�"
�`�_]^�H�^+���p��(c�4+�q���� X���.*���i�6�z�� 䃔��; ����fq/��GC�c�@�~�H�����)	��S�1h�����F���I�n'��s~pp$�=�PFéVa��y�NM+*��>�|�}�]\�#��{�=c?`��E�fO�k	��o?KT�l9W��A�ʛ7���핌��w�����)�����)�i�_S�B ��u�ǨHn�մ(B�1�b��ak���F&/ �0f�_X�0���<v�U����_�鄄��ɱ�><��������� (Ǆ�h�V��{+�fրd�X�R����l��:� �L�z#G�Ǵ�i��B])��������X�+���I�*�V�f0_�pa7���Q�UP!���l�T�6���5��/�
c=��~�~�Ѣ�o/�?P]"k�����y���%	>o��c3k��pD��VinZ��'n�JJ\�K��JK�Yם%��;�V�Ӷ
�X}�����j�.�<X��t�E�6ZO&j�B�C~������0�ԉ����=h��։��Ɖ�,Ӊ�B��B�zk�ck����@x� �E�B�)ID��O6/�_������s�`�mY�r�p#�?"aYB��k�<6E�Z/��A  ��QI\S�h �2�j�
BVǪ]�86#��8&�j��¯%?�}Q�p�jXZ��31ǳ��*%�s?_����<i!��p�Gx��S��U��r�p���������,_[szQ��
(XU�*ƯA�����(e���:����ܬ�j��_#.�����|�?���5�ҏ%��y�;����Qe�
�
��V��RA�� �fd��<'AC�(qיEU$�Xl�2]I���-P�Ғ4MME�$m�,3�󰴱
��sm�/̔k����f��[����p|FT�!�,�guɅEK)�]˵,���1ɜ�1˺�Yk�?V�5r?04ވ�$3u�jv/���o�/��o���oI���Ɏ �[��ַ�}�[O���o}�[߾3m�ˏ��P�Pj�Bq�^���!�h��M��^R� ���2 �SY.���JY�p 65&զ�m���7+*>�w�A����ă:mM�υ(���h
Z<�ɔ�߰��2lb�'X�p;�S����$f�b�Ђ��`�`m��t���]�6�JV�īi��
�Ҫ�E��
��zQ�������_kw�v�*7j$��Ld��n��T���@;  ��*�s��Td�k`��p��9�D�j)/_���e��<xpJ%�t:���3�&z��f>��R���\obB�B���Z��w|��ݝ![N�=y"��Ǭ��
�w������v��
U��P�a&(x�'�X`��h�( ���v���l�o5(��d����>ԓ(�%	��w�;Ap�J+�F��z7@!h6���%��5��r]�[R�@8�b�טeP,�h��R�j����Z3��1I��g&KȺ ��`���fyS�e���C�X��+�5Ux�V�����3>8$��5�2��g�@� ����n����e��V'�90��1��\<	P�U�~^��l1{.��O9Fa��-6�x����S��mE5�S�5 J�y[����*�ք�瀪;���k�+R�/RҶF(m��5M��ő|��g���#y�����]˛7/5?"P���l�B�=<�ãC�� �m8��`��Y���n\K���g �0��������̗3�
)�W0�LU��y���oIdd3T�f�T6�iUd 4��.�A2V��u�j��V�s�fY��DY����y��9+@����gϟŜ?9y /ߜɽ? ��h�=[�ωC�Pl����m�S˭f|����̆0����. ��Z����f-�/�k�A�w�s^�n"��.��%J��P(���6��ʮm�%��f��iK``1�B�$0��jи�S������w��ᵧ5�c�q~0T?cM ����y�%B��aAW�lI��5��A~|+��>m��-�6/0g��X�_���v�NcPV��sl�ٔId`y�[Q�Gf�X�6��R��5�M}-�p�w�)��`�Y�V�n~ŽI��5�����8���P��Z�B�C�jvG�<�!j�|�R��# e�Fb��o���[f�)SX�Vt��T���
� ��1B�̲*���y�H��jL��"Jx�<�����$�>�]Gb��h�E��iXc��(D��J~������TF�H��&i��^E,D[�|�kW��Ɨ�:Xl9���3u��-d�m�=ˀ��ׯ���D>����ٓ)�@����H��j�ǉ<ؘ�����N�AqՄ,�Fs.���v�u�ǌ�]z��h�߫D|�yc�-�^��,��_"F����{Yw�h��˻{�{J����r��63T���n�f��{���=��R��]���U��V�"�k�_�|_BQ��պ��o�g��o�/~�����rv��s�dvGy��ַ�����z�o}�[����j��\�����Xݶ%���Ѓ�$j͒*��vI��V���D�p��ah$7�3V�&#��[�#Q�ϛ��P)HOlbs�j{�a��U��A��q��!$�Qٽ*�� ��Iۅ����F!����7���4d}��o�U�q�����GjVVٶ�6�*�F�%	�;��%�T�Br�5��>��j�R}���H�w����߳Ѭ�D�?�
"_���T��{�kfHi,�`�0q���+G��x��LGZu}xx$}��G#��7�a� ��jE���X�k_!H�)� ��g�B���7�`$�@ M�&=z�o�o�`k��t -lLF	��J���}��[ۥ	����+�	 ���`�Q ����\	�@jĦ�A5e�m㼪g��/H� ����WT���ʟL�<���q��PF�C9���fɸA��¨��$��D�@~.J�.�ʐ@ZK���R�D�\UF$*aM�oJ��xX�6�����\���Ҋ���P� �/+��V
��l��M*�YE��N}6>�Hk�J3r �b����n>�q+@�������l�?A���S��@���^�-�� ��������`���%+N�c�K��!�ӊQZ͋�@S �Ї:6*������;$4	F�`����'&��X�ө��7��_����V6~}T`���܇!���1�}����������P�xl�"9f�sB |�ٶ�-�V�~U�$nA��>Z���\�,�9�$ ];RĊ��di���P�!�@�0�l�F#?ΊV�늪8�%`��-Vَ�����ǋ��@�ҏ����ةI���J��,�b��:H{#�k�����L����O�� ��/�"
y�m�tk���Zy�'6%\Ԩ�@H6�����m��u~��b�Ɇj�I>��%�$J2V���,+(�N�m7m��,A�9X�q�I��m`lcA�}]e
Bc~֪~�5�X�Q����QBR��P��t�a�2��)K����uII�6�3vh�s��@ ��Rk���S����w�K|6�5�U�s�9���u�6���k��x�>�xn��vM	@���v�ޭ��s	��ڪ�1�^kqߢꙊc�S�=���}U�cJ޽��׻����.�'ҹc���C���Q�����A�Ɩ�`���#^�i��QP��R3��HY c���n�<)�_m��5�㓩qPż0U.F�Z$ETֆ�5(o�+N�7��~ �����$�z��٘B5�t�h�^K�I��mt�@���zd:.��T��D�SP��9�-e^�i�����<��9��֯G�$����e��$�PP�����i1��.uc1������h輒��P�#��X����zG&(�`�q�ʪ��,Q�s��C�<8<Ѐ��2�VK[�zT���#g��5,'���;���+:d�NI�����>Ȭ�ǭ�Z,Ǝ�&c��s�+y������N^�����<�i�&�ӿ��LR���ῑ���o}�����H��ַ���;��fănl��!&��x��Z
  g�~K��vD������s:�N|6j3���Qx�b�Xf�4bVWx�D�d�DFS��r�)iQ�	�^�U����foP�ʋ]�2����i?���C�0� �5+&���a�!��gT%*ء�R���J�@H�$U�i@kAk1Xj�0X ;A���J��zF#W!�����B�/݃8�������JN=��� X}hF�qYf�(YÎL��1[,�V��<N\��T�3�y�a��t2�>�^`1��E�,P��k<��E��{���=��xt O'�i�~@	����Ĺ����[5
h쏵r�ꂵ�X+D�\q|��\H�
��VE$(��ڈ$���̢D-NX�
p�2 4��:Ihg�0�2l��|-��^-�``+ȁƬ�8��.��8P�¢��Z�;Wc��������54f�j��z��� Yx-����+�+�	���/%���^K�*�����__�2� ����A��i��!ŏ'#�	�g��h��N�)�$�Fq�PwX�4F`�j�n&��J�s�����4�g�Ì`�H����;�^�~a4:>��X�q��ٚg�S���P�|�r[S�QS��g����g��?���v>��#y��߇�.W������n�
�؇�J�U�$pUnd��#(��R�T� ���m��~�dq�,wC!���jj��|#�%J� !�ӓʡ�tc���LK�"����H�#����`$2�%_�uX��� ���$M� P5�n��][J>HI��\��V�ے�Xn
k+APC��9;6��C�������r���q�+�櫽��z��?P<x��
�6THU����`�T )wVQt�)�l�'F$b��|� $����]�BİZ��>��ov���`�5FT�h�;
@Da~�l��C;����_�sI}ߎ�#�T��H�`��T)�;@�.��<��u�����6�Xכ��+���H�e �F�G�G���]���T��h�`�y�M�m����S��ဤ1�6]x��ɏ�.J�xg\���2�'�Ns�]Q���>8�A�����ֶ�gZ��u�:2(�: �uv[�?��] Q��``��Cqb]�0�?�Ȫ��R���t�/(�d	�����bL�v������Y_A&��UX�tT���Ի�*����&(�0�P��������vk��x_RRu�v_��~��)�w���
�}ҩD*��Gs/cU��Y&�w�L����P��zIV�U������ﱪ���T$faf��b}��,N��H����J�����Q�Q	��V�y�x�@Va	
s�`8��m��K�-��U(*�TN�����Qy	�4�����sF*����*G%�x�j��P2��-����b�(�;ɮȢ��
�>W��>�eT3&Z�Ü����T^_�< }�[��ַ�y�	����o}��w�!d�8�^^���P&�qZ�!��=L|�`���1+�SV��1�*o�v�/��cv"�.JJ����>��Qp!��8�VUU��fK@EĲQk� �Ң#?��*��:O���I_�V �����v����5����a���� �*_T\cPiG/�T�  Ȑ� ��VOĚ��� <9�#��u��6/��ΠDAFG���>�گ(�<.��J�E߬ߘ�CAO�od����}*��R���<��/�%�_J
����|�1��A�z���>$����ec}���̐��?����6p�Y3)�|�tr(_|�9�"����d���O�#�Y���{�1�`I�y���� :��+ڄ�EN!k� ��a����ی���y��F���FmLL�s���	�z`W˥*e Ҁ���U!���PJ���mk91s!r���Lv�� P�� #��s�D�?��&мR��M% ��yu�
>����G��r��sg��C87l�4�6�rSJ<�i�U�#U�ĩ�o�ٷ�{nU졲���Q�EPKPs�����ZI��+�B��<� �r���}?<8������{IM+�a�o�}���o��;J� �n�
j���u�f�#��i,�7P� �A� �1v�X=�p���hjVgcl5\�
��L� J` 谞�6����`�g?�sJZ��Y���@�`��?@	�Jj���BI3%N�x\�ՏH��)��j��@M�p���/`��D��o���Os�)���ֵ��HH6��[_v� _����x9'ȉRW���*s�� jF���-	�r���d4��@�ټ�uf�ٵ!�0-����·��]Zj�&�JHv�l��X�9��#Vă�!л.��=�����R
���k-�,���; !
vd�є�'I�XA�T�/�+U��s�ܬe6��}6��m�؋#��Af!9�	�F;�?4������땂�؎�!�
ۨ�j��]@��B#�}#�6�~@NO˱[���H���'QT�*��n������(�:
�W�T�qG�8Qu�ɟ�}?�Wg������SUGk�U,�@��U������*��G]Z�gi�W�eh����`O�$J��}��S� �{�7�Pȡ�vp\�*%�x�a�~�
$hk�rG�d��º��BEC%�ۘ�Fi�-Ta�{B�N�B�7�j�$�x���2���v_T��6*RKVXG.�K��Q�縃"b�$��k��Z*!���m�Rsa�ղQ ��ւ�U�a��?��Wsɨ�rF�՚��nW���i��/��1���_i�V�����EC�C�OlF/_����!�[-\p/��:,a�U�uX�T��|�H3X�q�TAm����u��F���
Qp?Ń�_��V��*t�`��[�̹�Au��1�	�٢f�[4_��ַ�����z�o}�[����jT?l���Z]럂������U2�/�:T�#$vx0H{��� [>�Em�X����"�Q��:�Zl*:�1�SM�]W�ۃ5����C�rj��Xv�>]��U��A@�2��l7� ���ȭ�]u/�&�y��{v���4� sg Ğ�y ��T-]���"��� ����hX���*O��m�Oh������C+�S<W�¬H�ld��>�¨ ��+�#``��kF�������r&'G',F�L��O>�?�̟x�o�ga��;����GX�7:�% �~ �߯�<���9��V ��p<���V��ZG�Wܦ��y��(בю0
����b#n�D!�1iv'���
x���	�5���A6P��7TX�Zb�$x� ��%�U��g��R�\�+?���6@泡XD����ځ�&�P�&�}B%���8%�rC�8��_Ʉ6V+�$��F�� 9�z4dG�ٍ�MIc��<F��B m��~P\[�4��ڴ$ �B���� ��4V�Y�;_b�WM�������2�1C%}�g�GV�D���j�`�4�<T�O����@�i�{�fg����w��-ɥ��\bң`: �c�믿���?�o���\>���������5����J�	�q�!P�XV��R-7\�R-�ʢ�<�D+�s�s��_X�c��ƱC��0���6�_s��(���S���@oq�@�@��s+�ۺ�H���gc�`�a���Su������

�0&��cV%��̬�j��0�R�PJ����"N�*ZA�x"��;w�jM��%mc0��1�i�V_"���^vH�8��Va��o�ޥSF��@TTa�>x ��Xno��V �H\e�=FJ7��i��oBr-X�����M�$�8�&Pj`�1h���r=�������p� �Y���Ֆ�*(@�����_�K<#r�qGl���س�b�M�&0br��_�u։q⺿3�#��"��"�X��K�CZ����.r{��qg�͸�K�'���
 ��@���V� ��Żc�1�����dh��ޯ�J-6�|���C�'.����-ѵ������ =�#M�Du��6���؍����ײ˧
]�Y���9�ѷ��
��m)��^���Ŝ����$͠l��C��0�P�4Q[��~��T}��Fx�4"B�ͤ��F&��@L�146��ǚ-��F7UK=fZ��$g�ץ\Cv�p�m���p?Z����b���7�i7�*S^�����"i� w��\["S�5�g!(��{'ܷV���6�in�Fd�͚p1-�Lꪲ��?�z?��y�W����[�6���9kv�ЃB�;���}��M�ڒ W(�xN��SYV���"�jA� �u\aCqd�������c9/��g���aܪ�(���\���Bi�ȐE-rvy�ƓI�_��QGm[��������?J��ַ�����z�o}�[����kAA�� ��lh���`d�q-���x(��Ǘ����xH�|4�nBPY���5�r�eƇ�g��`[�]��-�'���|��v���4`�`���GpU��Fs�P��W����|�Q*��˲ZS��!�f5���Em���X9*
�$#���@��~eBe!��Q}Ͱ%y�(Z��Qӄc�	 )Aゅ:�=�F3?�`
P���A�Ł�r�a�$�paje-%�� ���W����v.K�7��V7�����PU�����F�<~B��T���p��y��L��^ɺ�d�3�߷����-��a�N��e��w��(f�5@� �!( ��͍�/���=��.Vřu����(�O�=x�[�=�cׅ]�;� !y7TG�Z"�T�𥤭@�ܪ���?X�5���t�Qi��P!J�y��́��z�5������`M�
*,g^��}[о�/y>��(��9��d��4�B �GGK�\?��!����[E4Ȑ��:6�9߃�}'�z��~2������fȾ�['����d2��2���}��6�U���_O�6̓�Q��Bxm�jEk�*����ɡ�k7��[b$��2i�v6:����O��� k ��`c@0��
���%,1B��p��/*�o�?���`���ׯ�����	N)�>ө�"%z�P2���Œ��65P�e˵��"��������a*�Fr�>`>�k���� �[ΡJ�B��ˉ�)@���I� T�@薆Z$.`d9�oع]��\�� �:�#����͊s'v'�W paN��[��:A��ޖ$"	Lc�5[2� �ǦN�:�)=�Bm�jZ4���	$:w���4�|�Z�G�w: Ї~KM=���
���
!��G���^�ePD�b�߉?l�F�5h�T�|��+�$��YF��1"؋��r��2ȩ��5k<�n�r3��=Z���A��{�*P���Z�1#�F�m�ۅ!��+� �5�U��!0&P�4M��+�Ő����[�u�N+�S�����~�h��ߎ`p��!��:�f��\K @@���BC��z�vXs3�dw�*�����TF�+��k��0���	@}7֭`�s@��Pc��6;;�`��{�J�����T�kF�V����hW(Q����yf��`�q�{���Nũ���0�����a*7���z^��Ȧ-���V-�B񁒧Q7��T��BqK������U��6W۝��U �+��#7w��2�S��ˡ�W~~����4����_�ȶ�o@�Y:�`��vRH�g�Q�5�[���^
^�#g�6qIu,Bxa
��y%�*��_�!N�>�Ia��\µk���f�R����,��H�*�@p�@bp���VQ=�*����wJ��������u ��,�:)uRkM����
�J�$�?_]\����5db�#f����1T�+�[gnꯝ�!�G���>9:i�i��_�ٿ���)"�����ַ���o��� }�[��ַ�Lc5�5�&NF9�s����}� C�V37wA�� c��\ITe�Q��{�e���
 ��[.f2��H��[�V�!�b |�f�mx�]�vC�*%	}@�gtY�C~ H��V[�id�x$KY]m%�|gH��+�%�hC�����3y�V6�X :��P5�wj&_�c�6���� 	��6��(h���sO{��Ջ��~��K	l���5Kaa�PSl7
��9��Yh:���G��F���l��%	�VOL5��5B�+py%kZU�����/�kJ ���q��Lպ
�����@ߔ�%��.7�L�C T����1 浼x�Jf~<=z��a�Y�Rt9::�z"��b�b�N �0F*(����Iԇ�[�he5l����\i5��9ښ�y����c���*�K��󧰊�����hՂ91Y���'�{�ޓ��L�޼!`r}{)T��?������X�Jn�Ac"(ސq�*�ӓG�Oe�\���rv��%A � �ӡ|�����c�;��'_�ݛk�I^�B��0r|�D��@F��5���/̽R7�C���_�T%(>�*����>���)_�������`���α0���u�(��dS�i���"W�m��N%�'2�]�Ϗ��a+����������k��O~"[�~��u�$(� X�k�,����FA�
�������2�e&�N���������sߗ3����ԏUT�҂��"��m�Z��zx���~-�;6���}8���j����+��h���7��9��J>���*9:>��<���X�� )uqq�������/���*��)D?�\�ʣ�*�TBA�����$Xo땕û?�sb<������Y~��;����ϵ�&$r��m��߷�V���=�����ߗ�O��w��~�|��k�yb@�v�[�߯��L�v�5��J��ډ�ֽ4J���Ŋ�?�$\�A+Y{��/�#���ɘk_�h�9l�r�goV_-�ʘq=�������,�O�	3_�j+�_W�u�'��$��^:����+�5y�R��䬩�?y��ݔ��Ef���k�U{>-h����x�)��پ�L�1-����A�dTԤ�(f@%yl9�oh�]c`}�̀���	��,�C6�Y�8O������Tŉ����]wj��Fj��
`�~�FhJL8��񟍼�������ۘ��I��ڭ+Ĥ�q����0� ��,Ϡ�B{��o:R(X��z_#�H� ��F;
(X��Ht���|a~�F���Z(�X�N~������G_U��{��rO�v6�}�
)p�����"�8��n̐B�
	*,�5�)�����)���{ʜ �aǾM�S�/�)���#']1�{;�P1�z�C�ғ'O䣏>�2��h��v�9�����s�����] ��d�󙯇��K��P�M�j�5p��H(��cn����w��W���ƮE��{���5���c����v�(NI�z��̲��y�:�cЯSu����#�p���}�e"u�sN�3��I4�<7?o'���Bn3�JUϬ��2	��T��p6��z���uNO2�e�Z���7B�� j:��KY8u}��u��GGG�O�PV��?��+~��**�o}�[����n=ҷ���o}��4ó�����>�3UC���yz�_}&�ш�3A�Zݚd�ڱ|������x�������7G"��?�¾)���GB[
�� 0Vo�w�h��6@�XFȻ�TԈ�_�6IW���f˒dWv��1���9� ���Phk�=�I&��Af��#�#M��>���F��n���
�!�rΛ�Fܘ�G���>�?���p��q#<܏?�}��ֲ`\�[�d�p8RE�GhQ��m�P���Â| &P�	�� =B�P�?vY�=T�#��}y�?��`]���Z�I|}���Bd�Ù���w�U�qj�Y���nG'�/\�J.���4K���VwsI_tH��
�������㇬��ￖ��ny��(��,��0�_u��`���̗ (�@t�0�F�)	��.Ղ�"`!�!à!Gh����<��J����֍��b���q���s���Tj� �i4�w�aO�u{2�@��(>y"Ϟ>���P������n�UA��~����³\U>v-@���Jy=�rr2���K��z샹;6�#a�K��³����Ƀ���>)�U �G|��I���9�0��s�Z�K�VG 8���\�s�#�:��buG"�L?�2�e:�ʏ� ګW�|������$xz�!Ǡ+~�
f�O��e*��X�����w�%'��SH���w�xA0���훗���@�w� ����Z�AK� H�6hp: � ��h3Tiw����c�v�<������r�ࡼ|�B��������z��F��P��sT=��m�&=���B&�!i'$��y�
	��-�Jw��;n�Q�����$�`7u��R��)�'8�_��+^TVT�Dn��T\wɨ�95U/:_d�AD |fv�Xզ`�fD7ߏ�'���G�x��������s����?���Ν��l+α�����t�ݘ]M$��F��;P �݅���+Y�kT{hP4t��1����|T�źv�5�8j�L�h�W�kރM�V�&�'�����f�vfU����J�� �S���o�>����g4�G�؈��Ih���-�ڎ�;�'gn.�5��<7�N'#����qGNO�|{r����5�q�u�0��N����Z���@t��T-�̍�Q`TF���!�W�+���Q�,8̷�sP�
L��f�-U�����OJ�� O���őZD���P�Pm��V3�W0~�&�e�O}د?���׼Œz`����v�U��A�Au��Xy�"��	t߸�:���Qֈ߶�+7��2*LUq��ı"c	$�$lN�m���`}�*R���0��� ��M�2J���d�����u:,9FA/7[U�`� ���~�ko���_ўS3T�Z� ����؇���V�@+����ʪ!@���lϼ]��G}�w�88&�vu �p�_�_��Jg(�������x�%�l�6r��+dv�n�;P+'�B��nv+�պQE��q�}q��?�(������S���ǰ�Lܺ��mx}�â�_W��3��$q���,�5�6���q�Il�O���x�嚙!U�2P�2H~ Ks�Ҧ/K�w��p��S-ƨd��j����u�"��v6?��;9�p��s���T}�Mƣ������L���]�8��Ҷ���mm�A�� i[��ֶ�}���빜���xX\��2z�"�=�!� wwЗ�=���'���L���zɰM�g������C9@��d�/�BT�I �0�= ����s8��|<|����Юa��xT�:  �{D~�w�^U�DBezbvx0�+O}C�:�?O�/̒�z"($	P��e�e�8�q�~T%Gj��0k�(f��H�xH����"���-�VĊ�D�P�O��VYZY(<A�X�!$CČA��?�6�!�P��հZ&�唈'Tu��fr�Yʽ�s��NYA{qu)}����*�����vQ�ًc_�*ݽU�!%vc� (2�7�m�Q�4��#+Ecl�͡��+�U6U��t��HJ �F�$�m06Q�a�r ��ip�V^�(@$B�
!���@ߏ�IT� y��!���]C�	���D�DjP@t������ ��۟*�m\��;�H��^q���Cw��|��ɩL�#w�VTJ�GC��S�|@o�$,�l!p�1R���	->�����첵f��\ݍw�Q�M+�~�g(��H��>z��%+�C;% NC�lL�M�0�U/y���6��҅���ɝZ�N���~�./Y	<��e�YH�3@�;�{wlPb�uȜ��a,슽23��u�J�H������;dzqO�m.��˿����_���=�/�29�ˋ�O��K�x��F�M��ޭ8��n캋�����䓏����5�!�+ * p�u:;���)�Z"{#����>ɕ�t �gcR�/�8�Pe��g�˗��Q�x����D�\�����+�ẁZ�{�X�V�5�EKZ�j���սG��ß�?���A�$�������&��_s>��Ь����������B����-A��`��Z����r�2�"˙��H���Y:.Q-�����\n�Y���I���ή�*�ּ ͚�m-#	s��x_Q�R�ڦ�]� $� �;�f��P������%AEOިUOBbs��86�'c7_<���_=�V���V�q�N�؁����`,����I�ZQ�\�͎s�x:��ͣ��^��ZW�����S�Q���ǉ��rH%��ğ����Q���*>w��n!�r�8���5��C4��!������p]x�FyTɠ�_� %�W�s�33��֋�)~��,�P�Σ�\K'Sc��X��:&�*����`�d�ܖH��21Pe��f��駎�+���F�VoaI���)�g*��Q�SfM�<+�m�[���q�k"Ƶ�bA�o�4W��\�{�ҍ�_�ڻ�r­iת��;�~�v^�\�-��QZч�qRB'�~1�H�V�&*�R.��n>B�ͮ	/,?�-�/�Y~]�y?�~.�Qcav�����X��Eo���# #����;�u������ ^_,�cE(޿s�>o�]�r�������b~��>�L�}��;��G�E��;��PJ�yύ�¶9���ް{p��K?/A����.`nQ�ES�럕��b>��jCs��+�n�=��Rj���m*̺E< v�M������ed�﶑�����7(�(��X�=��twhYQD�w�"�'O������mmk���H��ֶ���{� ��Zg��MNW�8�
���
�@J[��>��aq��wkZ�t��6ڰ�A�u @���oT�y�ZE��˴'�Ւ@��`5���3,Y�H5C J���j��
�G���ʀ`�j�U�0] G�i��3q��C�=���� ��&���\��9!	��{���_�s�V� ��]V#�eS}K˔4�|� 4{-߄� 9�R�r�h�x����V�ܪ�4�z��&����3[�2�V-Y��c��@!X6��78�C4*������]K^沛�h���w�6��U@ =Dɝ�.2v۽,R�#����`}��0�/��*�c�Q�t8q\J\�]�]���[�>X�����B���%#W$�h�����w�A "�ٌ�Cn
���r'�͒`"$ �9�ǀ��	�Z�p&n ւ��r/���؃�
�J�`�HA� p�6qm�ܠ�����]#�,����#��ہ\�5P�*`��~��չ�B��_,�$� ���;1뎁
2(!*w��4��-�+�W�������������c�0j����3��B����fp�N�c�$���t2���Umm4T���y��t�C׿Pk��kDK�!ͨ�Gh+�5[خ�9#�h�u�����������9;?��������y�v�y ��.״�H��s���D?�/g�SwVr3{�͞xx?�$L��ςcCƋ���~��� G`c��;��7��-�q@ɷۭHt�N����y]�S������y�q��D�(Ah2��=�Շ1�򣴫}�T��f�ϻ��H>���J��R�޾%i
%��9���d����v�~0��l��9W�>�9杴I��Ӽ;�����K��G5<T1 G���l��B����3;�1����ʁ�r�h�T��}遟��I���?�)(�p~;�V��R��w���l*ݗG�? �N�5z_UP��'�������S���w�O�X�^����ݾvV�c�_a��!�P���&���<Je%TkU"�J��a�Ѿ)�-�fr�Q����ц)ӌ�(Ψv�5ب�Ce�����@\���}�q�;�M�C� ������CR�h29X�P��u����bT�&��EeC�T�2�kE	~m�.�6效Q�˷��.��&�y/�|F��7�u3��.�A��s���>Q��{�Dx.VF���WT�ƶf)�H�a�ྛ�d�$]����+-��jXyc�߬v�w����vN+��U��*���\�*�Y�����H,�[Yo%c8*��RR����T7�kǛКI��@�Ryi��F��p�kggn�=������!�ǔ}�l���G�}����}�7���5E�O ����} �%���4��N�wa��F*�C)�[o8fFC-��{����B��PJ�W���E�l>��EHn{ۍ���1����{PA��Cߋ���^�A�E�[Oƴ��c�'������w��L�k�I:9��H��Ȭ���	��+�Ϋe4��$���tW��ad��
�Աmmk[����n-Ҷ���mm�޵��E�1��K'�è��k�><��І�5  �v�Rr<�x`^�b v)$�_u�����tSF�
8����5Lݶ{T[��zC�"��{��%��x��`����U枼�`wES�k%A�|���#;�(��V�,%?�3�����aǴ��k�m�����X�ɰ�|����ű�@�� �pu��
�#�K�B�A�R/s<$k_�D��MK�XY��J~�]X��D0�<��Bb&�U�P~ �3#p�l�p���������ljy.!{?y����KY�ֲ�f�Q<��!aLr�6`���XQ�t#�߱�`�UC��P��{x�Z�s�Z�ς�P�� �oJ�$)6��咹e�����
I� PD2DA��Jgų�AvF0�p����z!��� �N��/~A������o~�;%�t�%���� B�V���A� {�����]k3��@.��5P�z��z�l��\_�e��/�)m>���k�~w붗(�A`N���o�Z�eML;��!�gS��ի׬6�cX�j̇l<��k�Q����G�
�z��$踉�\" �ʇ:�T���9�1Q����},����2[�����r�� ��e=T�V3 ���k$�|��bW���7��d�AU�� Q��_ ^�:Zܭd���؝/6������cwa�nM�N�JD����|2��"���lO@�?�R) �n1��Z, ��Qq��%6�%@*�u�q����Q�*��\_V���^6�0�8/��@)��t�8�A��ܘC�5��T]�ۑ�׻'; X{]7���"�_��z'��D��)�l�z�Ee����H�+T~��qP)��W����} zo��OHj��#+V��I��n�K�\[�^'�6_'�(k�#֘�ԇ9�r�i�v��]g�� �֪�Æ�@%~��@��+��}��w���u�?5�2]#�{e��-�R�+So�T ������\.�u���K�@%���t9&p�.ܜTG)�i8G $q����xJ%��ǵ*"�ȡ��^��e���^c)�-{��&,� wY7U�~=S5�2��y��a���Pk�B�p~�؀]Uf"�
D�#��8�< �_I������>S�F����$"+C�ִ��I��+"�P `�H�>��g���[�+��$�F�^E��������<׵]�Z\P���=^ۏU ^4~'��І���ד4n�UQ�}���"�,J��Rۭ���Re}�&ù@q��cQBY#�o��­��D�M��\BU*U!F������J�8,L�
�p,�5�|y�U�����$@���sݰ�a���{s�W�=�'77rM<^�@�[��:Ͻ6p�`?�"�D��D��x��2��$�u�v��0�kf�#���װ{o�ͥ��:F���[��dͽ��P�b��*� B�Aը�*��.�_Ҁ�1%�0g����MIB͸�L�6��s���\S��=R�c�s]�����Y�:��mIk��ђ�=2���i�"�,7QL@��ؽL�u��t!6Wݤ��mmk[�~��%@�ֶ���m߻�DV��e#gWP#�C�XM�l�}��2<�,+�KP����B6����|ƅȮ��X�Ux��}'����nʇx/�G�D�i�|������3`��>�͎LYP��"�Cz $T�E�5ۅ�`+�? ��w�V�^m�2�' =|��0� K�yeu؏�j�~���ɼ�}�m��R��:�xx��jū>@�<ѡ���Qu�-
�)a䭰��E��΀���9��.���@�����@_,��!i��>����L�&��G=9;;�����9�h �_~�� )�@jk�:�[��
��<���@� �s_�Gy�Y����<� ��*_�o���~�%f����i��U��X��� ���*>����Oڬ@z� eb�l߄�R��~�RV�	�'O��_����~mW{��_�]67k���s��W' a d�6O�?|��ѯ��J�_��-F:�!�K1� :�t���o��˄���Ӊ���*�����V��$/}��n��`r���jWh�TVk�퉜]��d|BO�/����7+���2F0�x����� d(�ÇW���-ݜQ2�',�Ȋh�E3�	k������˯��W�٭�vy#�߭xĝD����)jUR�29 ��<x�X&�Wry�1�&�с��F��� <�W�����Qw)���ț�9ɿ���n���* +w���w�����'оPaSS��K��a.��� �W˵dݒ*�no,�qG&�Ý����l�j��Hl��B3A`;�>ں~�i3s\���T��{��{��-���]ñt�S�ݱ�r��D��P��cXs�xD�3���2��ƍ������-�e7o`\m@��
d�/1�(�����rZ
I��;�������f�}�Y }d*I�$�F1��Z�E�+�sn$ $_�*0�@��|��@Z1�eA��� �п����2�5+��_%���?@bR=��Nh�;m�TI�p~\�_Z�<+��{#\u�Q����[,	N�8a?_��6�~�z�B�OO����\m|@>�Ћ��p��R,����Ȟ���ܬwt���I ��%�t]"��\���d9��t�eSѾ�=��E ���>-|0.v�̈OͪJ���U�\���\đ��,h��ʟ�W�~5��(��<���?�~��X�;��om�n���}��R�WIz ABo��s��Z�N�OӑԼ�gC�p��P�b��f����ڍ��1��6s>�DR�B�,�|dI�R�4V�N�,���IC�S�d��e<oX�HE[���B����/�&$�(�Cf���[ZE�Sմ�ǂ9�,c��J�n�ǫ
���[��UC(���r6[��HF	_mLjJ�$��Zf�}�8"U���^1�d��<gy��j��?Tɑڴ�^?z�E������
.�6�{]�\���Sn��J:EW\��s��j ���՚j��������v��I�(:t����쾿����|���F�60М5|^���s�Zv)��ym��]��A�������mk[��ֶdk	����mmk��������Q��Ռ*�N�}�R+K�BРE<$j�D��VK�$�#�����f�QK�9���JY�V��5���>��-�������(��w�6� �j
�@+S�7W
�V�'��E��A[Q�cչ�Y' <�jG�Uo�|�! c6���� ���
Y5�\�@������� T
	�Y��@|~�8�b�R�v�8�w:����=+��	%
3�ڔ��� U����D�?��T�.���JJ���A�D�TB�>E5�� �����F~����<` *2	����9��o�})��L��-�ۇ��6]�Z���+`�f��b�i� �ҵ�s(+N j�Wj�Iß �&��m�񚇑Z�F�뻯����1~�������TWxK��|.ܱ_�]���s!n�����Y݄A��.le
VO
J�jS��?���߿/��D��N������Ky���
��fżd�`�~���w���d"�~�s��2����"�h�&á���=%6b*&�|���򭌑;q
�'�X�����ӑ;wn�.�4H��r!�͒
�Q�/?��g$����+�~w8�0H�zc��-l�j^쵎G�~�Q�㮯�áFݦ�`E�*%V�s��
6�& R��6���Sw.��sZ�U�U�3���5�.5	��]�Q�']ج�=w��2�LY<�[��f&I?�뛷���O1��O~�S�8�^[������n n�8��a8�0��y���\^ܓ?`n*z��M �6`U���ϝ��k�Wȍ���MSx\��܍Y��3��jx�h��}��t���>�$L�'�����܏X�!��;nN)ۜi$r;[���|K�跟}���,�=�B����r��*�bZau�L!�I_�.�H%�JJ	Z%,{�<�6�y%�N�m��a��;�P�����vYaP4��b1^T�H{G#$X�R�n����%�������)��z��(,X��BQE
:�
�h,��Z�N��ݛn�O���3�+(�*�:�kAM����{���U2U�kFs?��>Ř��2�PB!͊Њ	�в�*�~�=�*� f�e$��j��9�zɱ����XK׿;���;�$�V��v9At(`�6~�J��oT�1�U�r�ѡU�{bcUdQ5D��$��Tr�eSD�1�q�G�S}ﱓXe�N%M��U���� ��Ȏѷ�BL�Q��S��@���3*��g�(	D�ʑʔ|��<�E��ψ#�l��J�v�ES�T9 EHb��
}��]C�+">7Q�U��=���"�ù�����F4��yL�Hhw��O���L����d��J8�뵭��Ke1	��QA`g ̱v��fM" �
͘�8��uSJ�`�XGGRf�_U����)T�)�C�:�`����S�jK,���1�r)Y�P�zM��r���vZ���{(���*M�=��Q���
�9w��Z�2�'�F�oj-Pm�9.8�G�fT2�v�/u��T��d�]m[��ֶ��7����mmk[����i��ڬִ�Һ��T	<�d�F2����T~ ��$]A�@�y���z�g���(���]��6<(숒!���RE��X�E�kﲕ{ԇ4� @�G�D+�Qq��(jl��c�������$��)!උ
�A_A�=���Jx�JL��RZy #��L�`u(4��y*a�*~�䃐 �B`���V�z�l*I���+�-T,�EB��+<T��Ͻ/�8P�_�O�JTm��pV�J���|���?�5�$�p�J`iy�f>  ��-Sr���O [Kyw=c;@\x�ê�����V�2�<�*��DIO��� �ǹ�C��Cc�r\i\p�VX����>�Q���PB,�*�֛�[]+'n\�j<s���M!B��Z^���4x4J4ς��n�9��ײ����́�-����W$A �L�'T�|��GJZ����6=���^����ɘ����=$���g�ɿ���N����N��������"�e���; 	��~w('��N���c���/�P�k T "�x�L&'�rz~)��|���G���K���/��V[V�g���� ��DA���ř�7b ��b��xr*���yo��#k�][���� �ST�'�7
4�VPP���Ux�d��WP��W쳀�T`9 �"���B-R �(��>c#V���9t}�?T��z�U�ӳ��|�L^>{��p_���G��|(�}���,�G�B�y]F<��L��]���Kfi�_^�M� ��6�ws�W/���+�z��B�<�M��&�� L+�w�#���V$������ّ �3��W$l� ��!�7���׌VH(o˫Wo����׼���g��n9C��wk��[-�2�i��w�Ŏ;��&<�&v�1���@|n�� 駼�u��6���w�����̜CZ�P)Sj�{�,�5�:���2@O�S��Q 8+5g&��<��9u�64��+��}�9	�on��?QK��[Sa}�s	�`���O�� b�i� ��xB����R~{��V�q��2n8��X�\� fX�qF��!���kT?P�0K�1j�;���R�Z}�L��	�����s�*�BЉ$�r��`��b�Y��Gw>���1�=�@��.���7oA��ۈY�NP���>��@�~U���*������Gj��֮k0��.��m��u��|���uqA�ݝ�V��B�(�]�0Y��%�d+��SҐ��`�UE�4�o+����*��!:���մrDބ�U��	<6�"D�=��sUMP�`���
�H�'��$�;�-�0]��h�r�3(fy�����Np�@-�$T%i}��B�]�M�ۅ��:��N��9�,k;v�(�o*�c�WV�SkVo�k����?_�k�r�zM`.�j1�M^�$�'���轭'U<�JU(��*N�E���Z$`�:C�V�C�J	(K,*�%�W-J��#vstdY( ��F�Ү30�,�������`^YAUu�Z��IH")2,�P�>�}(	���6t�j��q��v;�%Ѭ\Q�!��"���h1����mm�o���}��ֶ���{Ւn(�.&H�p��x-����*�Q�=M����j:rs=��f+���n��V<��[V�]V��� ��6��Q�������mh��Vi�˙��؉�F�0���~��ش�(�jX�&���z݀fQl�t~�~��I|*��bC|����R�X�lT�����JV�@�	 W_͉J?�;1��u?Q��A�i���h�}A -Dr�6��I�����D&�@��T�}��ƪ^���{������J�Kd�ەYv��,�b������J�L'c���zU����4�ځ]FI �ų״�@�G���IXXG��� 0���l�!���Rf9t�3Y�7��"`A޽�G�� �Jd��B���G@/���-1���ކ���#Tjzq�R��6�MD�L��[ �ɽ�	$(��Υ׍e0�bu���T5<�k&x�@��s�^�����!����ݽ�:*���L�<~Lk�J��9U��% T���I�v��w��~���cח��T<zH�������Y�?�������;�Q�#��Y��rs���eɇ}"?���d궁Pn�JQ���2@y�������<��������\��lzJ���c��Q��5�!ܧ����u2���k���g�K�����'|�wo�����`�v��7���̽�rcn�����p*>�+5�Ԝ�
R��7r��k���́_ i�����ݭ#������@�SliA�p����p8p�>�����w�w}y���X�ג���cy��Sٮ�2�e<��d2!��j#%e�@i�D�ق}:�3�ʹ�CP��|$ӓs7�P���j��s	,�:)��\Fb�^�L�?��Gn}����ۇ<s�",��������M殱D
7UQ�k��ͭ���|�'	�׼��K8�Cф���P-�Џ�<�GT���d�O���N����f�!�Iܓ������T���z���y�g=�������g��P� ݜ����������圛�R��6B�O7v{n�n>�|)��@�S:�@�5c �S{w-��������$@������9�������4�ɢl���N��M���,�� �~�= @��.�dzM�

� e{�%����ר��3�8='���7�r���㏸���07���"O'CIݟ����#���J����X�P9Hۣ���xE�����y-
��W��^�513º��Vx,^ �l�MJF�S��y�؃ٕU�+��w�3����Ps����1�+XF҆��Y����# qc��^%�9��%8�(�(�v���WdVi��7~c���;�J*� l
5��[��u6���7�*?M�����Od��Z~	-���i��q�P��@s܏����1 *�n���a��
K�o��ZIU!Hc=oB��_M���d���FY	�H�,n]	�.�'��B�*@��f����my���C�[�?c����8,�X�Pe��@R(p�����+7Vn�wh]0��?(� �5�S�b�
c�À�� ���]� �Ca�N,�O�&�)�u���� �����M&�@�rɼ}b���kh'!�\�Z������N�Y��YY��5�q.�W�0#��Kj٠�����Kb�[���l���
EJ��A�� ��� �W;�qG�H	Ĕ��V|�x�cU"n6
OUhQ��}\���Xܑvc����R�p��z�QD��ܡ��7J�m�}��Ͽ������o��i[��ֶ��`[K���mmk[۾W�iݴ�5�TO��V���Ǩ�E�UW޻���F�I!��Fv��_{T5��<�K{�`�ƪ�$����s�	��X(���|�WOTC�YqZ*�Z�#���Y͊m'�0�јo`A�>���`p�/����E�F�բ�yk��l���I�yXDpW�����������[M±Ox�DT,�_<���7�X�m�	�)����?[9�V�f�\� M�vST�t����3 :��`;E��=d���J��y s��_JP29*��v a���v6˥l�+� w:�.�H3KDK��@���>
� ��5�$~�m�b jTEFꃎ�~�_�V��A��A�lB��ڀU�Vu�b"���:R�T�C�������
r�-s[ { ���B%Ic99��z$�x:"�����sVP�@"�*DQ��w����h9�d��t,���d4����3� in���`@�,+��w/�ݻ[wN.��~*����`�����l6+��n��7���ky�������ե����}3~��'O$p���_*�Pr�
����D��/e<>q�9c��O~���X��/~%W��d<��~'o�������"w�֋�/�ۧO����2���<�����9@X�w[[m�+�*Xsb�H�1"4��I����j!C�ˑ�Z'�p���N��9�כ�;�@ ���Kw8��h@O��Z�]%sׯO�~�~s-/^��q��i;���d���۷��vT��_�/.]<r�x��U�A�d{SbŬf�8�<���9V߽S�q49q����=��E�`���+q?]I�������]7��3�[ �-N臞e30P���j���_?�V��\\ޓ�I���ʧ}�#��q�e:>���)��s|�pHԆ����璊2:�3�T��U�q�^� ��/��/cVB3��ҹ+�sOBjK��0���٪��� �v�M+�Ќ�Z-hB�U��
�2��b�6@&WT�E�o����IX �׍x�t{#��Z��J���*�/��>���pD�d4�k�>__����Sy��![P^ ��<4������n�����R���P�K]'�g��@T�혽�(bAQj}�X/��JѯP*����F�H%T�'��_�VVp��32��A?D�eT�f( ���Ƈ5����f�� ��E2���r�|Q@�}��8r�ܛ2��HfX�9�\�:|��;���wEy���W�����{'^����8&%b0��K�����!���;�D56��k1�Kb�Pm+��,"a��*Tr�](��R%~o��Yl�6Vi�$�k0��Ҭ�xÏo��1�����[�#�.�[��U4��k7��n���U/�j�UZ����5�K{��@��X,o-���	�Z%y�>�J��ᵆ�)�~K�2�*AM̓��s H�nfTq�A�-��d5%�cܺ�KK*LPԃטL��A4�9
�����������q���{����wwTQ3?���6�s�Ü�y���\�N�9_߹5�n9�2��tB2ۼs��<���Ћ��}kwlw@��Η���b��f���&�ܚ������gA3�*�����t�T>qÕ�������_��������%mk[��ֶdk	����mmk����͗�q��pTٜ�O�Hhu�2*2ܳ�z�a��/�w��i�/n�=�u�,��5�ioR�:V���x@/*�[�%�*V�y ��O�V�}DEu��
GD#S�h�`�������^�h�f��'܀G4�'T�!�r���� �&�
�8`����(-h�7U��b�x ���xwd) �h�{P�l�;��}����}o�ʫ����4�G�
@ B��ռʑз���o��뤍}E�0���.���wVN����~2��|�n��J�D�Qu^i�C�Ѭ  � 4������\�'y��{��v��"\��� #GѨ˸�4D=��fEYZȽ�r���]v��40_�@��}�q�FyK�&=�ҡ2Y7����@�C��w�@��1��BF-(�y	U9;���ړ�S@%g�+f6�IGgwzjc�q� *�A��� @��z HWWWr~~N�����JCUx�AϬ���p�3c��@�
��w�[y{{#I�\#q��<�Qmq~z�~��k*+~�W?����O��'�[<�=�c������ �NϯH|���k485$����6�s j�s�w�k�C$� �����|A۝�bt�2�5G�1�� 9�q-�mB�q~y�dT6�>w��*��k7�������alRI�%!����5���w/e:���!u�������ǲܬ��u��c�7$�	���0� ~-��e��%K�Į4(٘;��$G:��A�`���oH�@9�W1���$�Dr����իk���?�X�A���J������Sf|(����I-dTi��֗���VbQ�҄c���S��᫥1G�:���nx�[x�߮�K	{��6 ;�׶n,x�p�J���"�h���`8�I�5\�7a>f�G�Y ��6a�697�������;����D�U�Z���P��l���~¿1����/�a����SAqvz.�|򉜟��� �p3�Ś
���]sn΅�a0�q�x%�&�z�s�.�n��`iv��6�@~��B�ɫ%�Un���DH�֪0
�܏��V��u�%��.�����X��~��a�Bo��,\�)1.�ȺQ�u�еqǌ���rO ��[!�~�;%�	]O���>�{
7@}�bU�h.�Sd6ee��wHeb�[W%@����c��}o�_(�ƪeH)��O�?���b��j���O^�:��#}��8���I��f�C�S#��$�&�~�U�^�@�ڙz}s�x�o��Z��{@e$��8U"���B޼}�J�7oݿ�r29ef���b�֩w$2u]�:E�%?7r��z�����,�zn	b%K�P�B}Ƶ���=!U��;�6��$�W�L\U��L{<.(ݶP�B�����q]�;��]�����o����t����퍼}w-������2�L�,^8=����;��̭�s���Ne �c�Œ�b4D�Õۏ����z�y}�s�"(~0_�������'֓��-�k��'���qX7�/�?t3�&�����?���,�7��o_J��ֶ����Z�mmk[����jx(���K4<��K��}я�-���Ї��~EՈ��]�}���^���lk�}D�Y`CD;+�AƟ]�^Z:
[��	��U�/��&����
���,��P�C=�+�?�j�%jsUXif�3.� �HA�* t����V�O Vxp̎��_�D-�:�zw�7�7�yj@�朆��M|�dh�桩c`o@<6,5���X�)�j_�j���VS�dP� G�{��AD��FI.I�R&�C>�?�R޼~'��������� x��|��%�3ˍ��Q��+��(T�!jt�d�M�n d3���A���ϑA�9�Nv�Vş74�.�U�J�<��#88�k�����`�'@��@p5���`U�f���S��uZ����?�>���ڨ�GB��$ļ�$HXiށŗ�j�V��Y�����7�LO	� Y0�u����
�����2^�o�;H��z���}d��/�� y�d�X2�!�#d��{2_.�ͫWb��[j�A�	��oa-յp�R~���O�쿓���">&��f������i�R쏩Ҹz����/?�;�=�/o�\sl�`��^�3� ܡ"A�7��CU��c��^��r�d���/�}��M��dB��t*����gCE �xM��?==�����n-�;�,b ��:F�D��ryu�����︝ӓs�w�y`7�%��r����nlaέ4_��2�Z	�6���1�]� ���n��ε;�"usB�����h���۷o�B�۽`<��޻�ޅ�_�*�����F�\	����+���8n���8�\��-E�K�>E-�`�ӣZ 0��ڔ]ܖe6�
�'�V�:ן�ȥ�	�S1'��,(����0����c%�*Fr`�B@��x��S��W��L���ޕ䛵�,������Ѡ/���rqy&K�&�u�۳g[V��G�QT�������0�}�$���� $��T���@�GCy��*˘e��z��k�wxr삔L⹄3�+E̱�k4"�./-��*?<ea$Mm�Bh��)��ē��\0�}v��9ʸj��․�g�(��@� �"�h����a��=I6�%��.�V���ā�B�F$m��~��=\���j��`�8�ﹶ�}�����bo�sBB���K��&)����'1jƂ�Q��2VHh֘eg�-C�`B+����!�<	҄�Gz���D|��NE��j'��Z�#0�{����(�v�,۪2K����p_g/��\?y��)t	�����߉��q��o�g�B��ĵ���_�.^��r��=fJA�p�浼~�Z�{�-ׇ7��:����dz���b� )�pM�B����X"�
����|��EZ�R���r��AO�Ͳ4�^��a`�[O@Hb2#'��'s�(|��$���X �K*�U����9�E�ݚ����n�n��c��nݙ-�r"��7�B#�1:$#:�m����}K�	� #4E3�c��#�uc���7�
�R �S�b�}�ϸ�@��Lb!���^�(*U�ǔ��{&��t/ȓ��d�0 �� mk[���l-Ҷ���mm�޴|����[$6�C� ���cڛ����X]����G������}@֐^�;���>x&#�S�;�]&Q�p`���v����iN���b��_�Cy�T%��8H�`�N�R��Y�]����lH�u�j����@d+�AV�xY�E�mIx#T����A�*W%K��WlV
`��F�H1�C���zG�e�YtT@#U���_%-!���AP��=�[s���\��v^��S�5����a$=���F2 ��u;�G-���Q��̼���ݖ��{�W{ =���-���5���W�y���3@5e��
R"���}�`b�;
<��Ȋ���xʇp�s�/�
 O/�Շ�#��i��-;*�*����c(F�,2?�Y���Hz �XnO�-�>ެ����Y=Pd�\�f�����9 J@~��O�&�������8g�4yw, ~`�\Erw7#0�|��} �0 b�*��}�|wH��gP���w���#��4"��IdqnЖ�ިh����/����+,�ְ�Z�e��+�`W��;��)"�a�X�|����wr{3�a&��[��<��{�'�Ϩf��Q^����[��>���-HY Ț�7���)��bCM{����L�ps{ |F�'� �#!�E�����g�n߆��Y k �K�T2v߭9*g��?����|��׿��f-u`ߝ����Kf��X,�`=����\��ҍ���v�8�n�`�6��b����;V��<�Z�%̋o�2�����>�q��l�\m�J�a��@�p��f6 >X<ἄI�*k�*�٫���A��N:�o>�/�s��;˚��6l��e�2�C�!�y}����{����n�2u�Fv`�ŚZ�E�7~d�5�B �q�
 �V;7�S xK��}	Em� �A���Ǣ�v)_��.6ă���^vc�E�2�,8/"�A��L��r��9ݟ��9bA�P}�yd0�I@`L��5?��uB���7r�l���s�'(@La<��<L�Q'B�tc��椱;7 �� ��1lݵ\�̱�{�1����.3�R��Po���W������J~ �Qh��4j<IGoo>�����^��=ص�G�C�'���"S�(I^)�����$g���Q��n�㱁��w�h��r¸5�A�k�c��G�A��Y�i���0\y��B��H%� ��F�;��ar�����F�0$�|B�6�qPP��98n+���Z���� �fO�{ l<��i�}Nn�^��Z���`��efI��C���tZfY�5X�m Vg���ȸ�
ta��6��"���7߸��s��*�X������&mOq�@�G�Vp���g�f�V�:6�iL�d1�yl�|���`>;��,�&@��W	Uw�A��k�9
�A��q�A@�������)���J\(�J��!V�X˳-�3a���b�!�5���Ν_�a3D$8�f#�*�:�,�M��u ��Ϥ�M2��f/o�kf���E�*a̟z���8�8Ң�:�8�������}Z��%��:
~�$z��P�q�����~��������mmk[�~P�%@�ֶ���m߫V�&!�C*	�N��? L ìDO4Q+.SV��k��/�O�SY�v�&��{x����e�\����WS&,+����C����*Q}ȹZUT��WӚ�G�ժǲ	!o<��g7ņJ  �>��9� .;Pfj� ����j�>���mPj�hɌ���9�͠?��'~oQ$�,����x��ٯI̾�����:n >�:#&���fum.��V�)�������4�Ԫ7q��<�n���a�])��W۲��*c�q�*h�u��w�~ ���7�$$.�^����~��z��{��pc�����ޠ#�~����^L�멶��Cb��~����o	�UH�ʕ@� �@���s.W�N��+� fԡ�$@7з��U�|	������y����=����Y1�5�K0�����E�}wZ�P� `Z��-k�C����e����E�z9c�?�sT��!+_�z
*x�W-q0$�=� �N�����(���������m���Dm, ��ң�y�3x�/V$\��'`�:p)�.��$9�)��ܹcQ�ӗ�J�����2� �3���hz��T�@�T( �r#�Vw���l��gϞs�_^]2`]��3V̒$��矪�P������e���>t���V��G$UL;�?�㱤��k�~����}�
r ���)-����_�O�3���������g�n��� �pl��U3�@����g�drr�c>ٝ��<��`�5k.�p��<w��C�k�� 77o���6zا��w22���V�'$ �?xVg��P˓���i�� ]���`H��c>Rз�6�<��4�>�q��|��w��2V��z�`�6�8N(�֫��`�VVAE�OPͅ�m���ku�'���C�^�^��w���yt�L�_X� w��>�J�8R���;���jmVw�~LC=��?�X!M�W<g�9�o:9����_ ;0�!�j���?�d�B��>�6kX�t:��@z�= �t.�can��v;�.��w}p���9�ʭ��Fv��3����9aDڇ�����ߎ���I�&��
��p�,�)à�^O��|�&��u)����\Q�g��{�PL5����l��Y���'��͔(���9�$n�`r��PHUl�Ƣ��{U���J�;\�T&�~������x-�s\鱄fߨ��0�Cc=0'�s���'Y�/���F�Gh������Jh�6�UA<�����j�������#�f���P�`ۄ�!�+�BS��x%_�}.fY*��R5-����o�믿�l:\�U.9�q�q_�LU<X�P���U%*kdh�~����A�W�>�������y�Ω�Onv e����-����9���xo�M���|CN`ˆ���2�4w$��=v�Y��ʌ$�n�k����"#��m�s��kKm��y�u�=�]��P~IA�q���T�\[����@Ta�)�g��djJb
�NE�m  ��IDATMe���V����.&n�����U%���_��`��KG�ֶ���m?�� mk[��ֶ�Ms�R���VB �K�U��� ��h�S��g�#��A%�X]WE��`���0<�`��*�n�X"�J�C/�6u߼��*"�la�~0�=��a���Uh�Ǌ�V�v�T��,NI��z�Ŕ^q�ݣ���<����v�m��Ъ#KQb%��YL�*<����� 
��R<0���zL~���<��j�>9<l����W\z�	}�u{Ȕ�D��P�74�$����uBHN-iDH,Di��oI;!T���!��f����듥첊�4�;��6C#�s��,�+Z+�</}%jm�X������k�ƞ��;�Ԫ	E���
��A���Q[�Q��V( ��LbAY��DB �ES�`� �@*�Ng��a���-϶����z4���R��|&���w���c�N��4l��w����{/��7�X«|MB���o���w��ީ�E�Co���U�v�X�i_��*��޼a��.J%>��>o*"�������t:�ư?�y�v�LF� G�����Uδ�@�kWA��j�����	�t������~Cp���є�C��҉�r��Ŏ�JVf��s�w3�! ]�/pd	2T�T���vRIO�.~Գ}0�K��� V#}Z;�x��q����B�.��n�g�6殎���ь�?;� �q~y%��[滀,�Ր{N�޼&�����{TR���e��Q�C;4�Y1�n��8䜙t9�kw�@���8"����GK�4�U*���
�=?rzJU�h0d8:�>y���	�Ix�*w9������k(`pB y��y�Ҍ(X�p.�\���d�ܸ��Z�y(UE٨|b��h�M`���f�Q��l���Cњ�+	��S���$>4;���{	MY�� �e��	u�	B��!Ƚف� .�Gګu�8_��2v� tE��ʍ��;�X;T �hPj\]�w��5��#7�����vN��w�w�@>G)�f(@b��\'���1��,ܺ�����Y4PY	碀sC�A*18^m�J�˨J�1�<��绣,����朑H�_P1Qej?h*�ױ*H|aE̜.�i��,%+1z��c5�V����Nh�f\��H�ǆ�R��sb&�{�CU�qvLi�2uT�6�B�6"#:�Ցuӷz}����M�9T���u?#�Vb�kS�*��V�V92B)���X����gA]�P�=+5��v��)�cFx��2-�P�_o#�}�<"{�!T<'x�3˒�Ɠ�y��v}`6`��7я ;-��A�PU�e���=Pö����h��X���џ@+0+�	5X�1�ˈ	(�`Zfɚ�X��'m[+��C�z!�Z$���?�
j�+����8��
.x�s��k�ZՒ�-Ω�|Py\i`=�CœVj�����а�ľGINU}���x�W�:,Թ�z���+�H�p:�I�E��`l���4�]���Jz����N�VznN�����Һ/����mm[��ֶ��`ZK���mmk[۾w��|�a��.��r� �Q��M�������t��!�n��CF!����3q'"�v�ب�D�?<��󺱛B%�/��xa��w��C��>4�܇� |��n���(*�ū;�&� ��@�{K-O4�<��nJ��Q���<rE�L-�`-�+�[��0R�|��"�-�4p;��}�U0��R��XiX�7�*dt�%���+
��<
,h��>�4:"� ��ʝlwC �:��l����Q�
�Z�m���`wKe�X4�JV͎V�c��c�׊��䄤�p�ݶK��ljugd���)�,��s􍷅�����fM�u��1tL��c�a�ъj��|�HA�P+�9>c �?��t���6A���D< =&p��- | �w�&)��d_Vru/'�<�����N6��9Ï�f3�!$���~WHz�%���	P�@�������y���M�kH�0K��( �z�0<�K�;�%5 ������{@���-�C���M�I����Qh}Ҁ�ՖE �<��s��o�LO�$?�{lv]
J�*y� � H���lx����Zo��ed�>�������9=;�����\�&p�?�aoh ��K@��n ��'�I?��y�07�ʍO�`ECK�"g1 ������п ۭ=���/����&�)ؿ$�9�P��oh����s&v�(W��S��OO���N%��oXi!Ǳ+(?VU��{c<�K0��0���ׅ��;�5i�m�q�[Ƈ��QP�������N`�9��(>���-k%5~2]��f.�Dy�h���"h�L$S�0���՜?{��Q����J{^��-=��FY�
�|��č}7IJ��H��=7�'${f�L 7��2����o�4�Z���Z���	{f x62P��լ�Q�Η�%�\�y#�}��P�������'�_Xl��nGU��=�ډVU ��4�Ą�)���D�����i�3'�G\�|X�p ��4��b_5�Br����y��S�s/����
�B�^AA���Q��_"���x���%9�(��L�\	��=Fa�{m�vXM��4����s6�<F\o�����+r@��7O|P���U���� -Bڽ��{pϑ��7먒��[Y����A��p(j�l����>
�Ae3lG�Ȑ#LKT_K#1��E_Lr����Ȕ(�s�����*�1�x��h }��f8m���l���w;aw_���xϷ�}Ք�#��SEkQx�M��Seh6Vɂ���N����*�*�$N-�踹5����A�~�-jc?ʢ�3���ybm
Ht�Q�\m��ć�G���,��EK�D	k�O�uߓ<R����3��B���Tu�mD��"�C�,R
��A��>��"ׁ�3����c��9$�D8z�w��5ݲ��>��mk[��ֶPk	����mmk�����a�x��Q��'P�~�A��!����a���J�o���Q���26�/ܿQ��l�ݎ�R͏��I�htl;%?��K�nr�j��}�1(v��L������H�
V��/��.'h����?�Ձ@�v;��>�������𠉆c��Lu$>KD+)C��J����f/ ��pv p"[ �l�7��{U�:M�_V���ܦ��{��O��{¥*�<��McU�г�㎷���ޕ@Y��x~���CP`�0��\�(5�V�@�j���[Z�Q�oʚa��a�~���.o*�a�����aCf���Cj� �X�Ջ�9������`_h�0�}n`�9	����� �N�S�>1u�~J�@1�l �����?�/7@G��˻9�~7U�7.�F���ȫ�od�k���> �{;��j���媱�����x(yV�����1��j����aWt����U����U����Q���@f��W`����t:��|�~�e��
"�A~ຆE*�K�j<u���%3G^��8��Ҫ
�?��i���D	�cU��#��@�0��� ��[�V�9�.	���� ����}��W��*X��Z���=9���dJ�j�!�����B��:�Q!��w��qsmҕP�|��>���o�e6~޽{'/_�vc�њc/���צg����Qr��;��Ϛ�z(`�|�2�38P���',�ȫ�=��mQ5��
�������<2q�۽�W���C��~ߗ�z� �`2��r��ty^jVP����ȍ�n�y*���5�?��,�,�4Ue2M�.�!2#x7��������b�Sx�ZAAT�'��O�o��U���%#^B���q ���uav���`iغ���8߂�s�!� �2wc�G���f�F97h땺��IǈL�|�	���T`aƓ�	��q�bI��s��5i-}w�%,B������ͅ�~��U����뼺Q:)!�� (����ʽߝ�(p�2]"^�������lW斡�� 20�b=��Q)�ہ�����P�:�����\��Z�H�R�F^��DE#_u(IK9��>�;�kP4l���<�fM��3>�}=�4�ʬ�&��q]G�{iC]�� ���9iqB��ȣ��}��Uaj@]�|ȅ��X\��/aط�2���Q��ZJ]c�@
��F��5�(do�W�:	ǆ��P�����|Tr(%à��;xO^eV�5��E��4�l�zev�&��>B]��i����ޓ�� �"�5Ԍ�\�^-�񳚽�
3����X^��-����Sd����ZO(ƒ���Q���\�P�q�^k1��@y�Z-CnJ�j���������Z��y�qL�MF�<�R+>Jُ�?�z�]��
S�@��&)�SR9�M��u�X�Z��,���J�c�ON�D��'\p����G�-;7/`�I�b�����2�gSQy��B�.��f"��m�ͿQpȧ˔t��u����
j����э�Z�͌��j�mmk[���Cj-Ҷ���mm�޴���{��cV]zl4��V���{�Ym������ c�H	,���gU<�+;�`Q�V�C�pՖA���Y^�� h"'���+=<@��ac%�3:"�����!��AG�0�}T��z\�FEF`���>�j��m�%f[U�Wɇ'Vl�� > �!� HU6vOI��|�pJ}��>������sKjʹ+y��VD�[	����E�$���,�r�.V�����<ԧFnŴ�ll)	`�l~+��"77}��fA�z}��*2����BQ���9�	D���b` d3%�<�8��J�G�6�1� +�cx�#���� @�a��UB%6*�Z�w��S��"J�R����X$��	@���$��b��/���v��p_V�E�3i:����7�丒�nl�g����4 ��p8�đ���hIO�y�h��I�4z�^j_r�Unv�Gf5���88�8����̈�p��0�f֗��󅜻��
��uw< "�쿥5�j�F1���� R$�х��l3{��	2$�q�{��i�{Y�����k�6ȕ�������ꄣ�C9<<���x�
l�*��fJP�pq.S�V�<�m�}��t6��ݎܹ�u}8Xߐ!��{���P4��I:��g�'�M��Fw�S*��+�"[���\�w��!~D�'�O�TI�p�"�2둡H3�J���] a�*RU���W��+Q�P8>=���#9:9f`y�� ^����������Qe��Vm���(!�Ԣ�!+��q���f�[쁠]��w��w_�B�0���e�r]p��8����]�u�r9YJmH;2(����1�ǾV5L���o�'�o���Uu��aᲘ,�ޠ��UA�c�/� b�C����hQW��
@�LWk���_ZH�*{0�5?�㎥�c��kەȲ{~��7 b@�h4���eH5��A���ª�����P��9�z��~��S ��ܕ������P٣dd�c�� �7 �[�U�s6�����c�n�s0_pa1�scd+�X�'��-g�,qN��������
�l7��F��5����C��1���z���-���]o�P���PE`�H~�)b��.�R�jy���,� � 1�[_���ʲ��\�����%���>T5��
;�u�E���$� 66�Zy��΋��O�����/T�G�3lQ���"W��\�qo���Zf�YY��� oy�^���Y8�2�v��𧜡۫v��{Ol�y��
�{+,�tZ�Y �/B�W,HAP�81���W�O�US�V�*��RF�(�QUG��X���&�-X/�zlA�N A� u�eޛ��7��[�ZriH|J�$�z�G;�1�d�֩.�/1�%�<
]i���f��ם{pC�fDB�/���ڊ��42u1�X�Y��EWɡ�_����9e���	s�R�)����|�P�-�r�����s��Ox��:�h����sޓ�8qّ�e��ғ�"���E��%f5�̷��S�?kNY��Ҵ�5�iM���� iZӚִ�}� 6�^��lZ6,H�\}���
��Q�͇W . ������4J���He��d>��z�"ؿ$? x+�Ue�VRf;Ԣ�ۇ�=x!#!\�ǫB��/��gx��Ĭ��@n#k�H��\��R ����F�[|x�kH����������ޗ\+�x��}�a���择����ZM�{��'���+�qk/�R,;ei%�!\�F��⺯j�v ��O�C{����^؆݆�F��/%)T�Ҏ���ׅ���i�-�g�2��i���pX(ml]�d$�0`7�A��y~����4��{Cp��c��Z4å"� 0���Î�u��xS� (�6�7X���0��:~����2�^�' >�Y_ۖ��3=w�$��X�ݱu�-��b�eT��g�\��U�V
�2c����;�K�o�/^ɛ���\��h.o�����}��$�B�� JΤW�5âU0�j�ͭ���V��T�7*�����M��Tɋg/�@h��[y���
D�bN�7+��� |;�n�S�Xg�{2���^樌'h��x�w(R�'�B�K�+���-��tQ��1�ǃ��UTg��
��������x@< D��a���k �bj��>p[����2����SuGY�K'�^�,f�a�Dm��ܖ��o��p���Ƕ��i�5��U���m��S�$�B�ѱ�>7���c_ �'��� �(��lh��j�3��c^���|��a�����u������eD�i��"X�]�i���U�E�Ji��kI�������	������4��&��C��p_�g%ϣf����9=7V@��s��^%�kye�gE���Z	�+� �3�m�]�\��w�z[,d��*I�.[d�X�l��qR�Wr��zPf��L�+b�9���9��8"��J5͇�k�C��Q���*Fk�+�+��\����� i�y$s��aa��I{�~�2�gk���̯��<����5�[�f���ؔ�?]��V�V��� Tѹ�|�-��T3)Z����fi�,ҙ\iŕoJp�ju)+�f�mcVP��u�F��!�.2�FV�c	���2�b���۵ j�_~�W#F���"��3`A�?�51��%A3Wr�*����:1���.���Y���V��չe�H+7-r(�זL�6�UI��Vm�$�B)�!���m6y/�r��1^)�4��}��en	�0�P����Wj�
`�zLbި���l��y�|)
O��1h�/��`�����Y�n�t(ܼ�����'�mmrn6o��A�P����G���K�JU+8V�;�z���u�}%CV�g�}it\=�񆖽�+���3�
� ��y[�}H������?�����or��ݺ�	j�7o���ٹ���d �h�k~n���ZL�΂�b;��Z��}	p����9.	�9�z��΃6����ִ�5�iߟ� MkZӚִ�l�(�ae:��`X1�=�.]
�����L���T�U
�*J�F-:�b�1��� �Sj�'3�['�5р*YV����T!+�c������G�J˲��C_=m��ՋI������!� n���C�9a�!1�a�}�}��i�Id���ew(�}��"������^E���	������T+�HF��/�@���5��tx�qB;��x�cV]�=n��J�����VOj�lI��'�lO�=l�v\zr_���X��*3��;�@���R)������eX%�$�硪2�[w?O�U�X���S�q���6Dq\�,a4Ε;p΍\Q[�(��P1��sfӑ͑-ڲ0�u�#Z�E-*z���U���oY���m�"~�JV�`A	���Wrz|�9����N/�2Od�����;�f"X�Ǎ�� ���vfn�<D�V!�~�
xN�8Vd��P9<<����2�z�c�����Ⱥ��[��g<� ���	̕��bu�����T+� {Z�N��SҎdc}K������l^������Ʀ$݈l�		$W�ޥ�d>�wT�W��EvM�G���m�D�x����YH��9Um e���tM[�Y�u	����[�;RF����<��K�����j�5TĂl �P 7�'T�@�d�$<٣���z���{ֹc�#�����F�ۖ�X�A�u��TǫZ��� a��<-�8�r'%y�3�AC�s��~�z�`���7��B�uwww�d���͛7y��q���I���m%�|.G�����s\�����:�X군0�D���,`�c���9����܉�����N�����x�U�K�"��@l���)����+�5�����HNOOy<[n<BS���I��Vh>��t�jr%�Y�N[�ȲRB�9�q�J+��ZF�u�m�k sd�s�'�:�L�\���������	c���5p�P��_�h�TF��v��*H���Z�ZHū�? ��J��Y6�����eK�h^��g�J6��p4����6��P��T������t��UM�� TH��μޚb����B���z�W
���������@�.�����Jt�K�$T�+)k�,��ᨏO%WU�uG��U��L�$���h�R8�㋩L�j�jI�����{� j�D������Ds|Z47e�JPd�i��~�
7��T������q�iw'����׮�
	!��S]�C+��Vm>I��"��K���A?o:����16E�K�XQz���Y��>��Zه�����B�6��P��j�I#�Z��<��
���."�:����
���f+�p��yϹ��.w�ݓ{���֖Lf�z��ݸ�����1�­�ݞ�O�t8�AK�A�ٶ�t��`��^��V���T�[HU}ޚִ�5�i��� MkZӚִ�dC�1B���*g|P�
�� DT�<����&�w�h� <��bQ�
<�g
�s�~��WV���# �� �-<������=֪1��תS�<���X�(�1R%OZL`*��h���eR畇~T�F��U��J5��b�$1���=AXcx(����*+�_���.Y�_1� @hU.�`Yej���h�5P
��[*Q�1�k�&�<8fkE��N&A���(�����j�P���Zti�:�W~(��b�w�%��`tx��$՜����A*���C�;j@D�a;5䞌fj�D��*%r��@d�[���?3Su[����$%UP�<��I��������B�9���k������T
$V%�p��Pk��
� #�6�Ҋ�e<���F����� �Ξ� �h��R�8�j��@�R�`�t��}�� ?޽y#�% �4S�����Mw��>]�~�@���Z"�����<��P�~�3(���!�( b;-�ڸ%-��[������k��̠@��;��������`|�uO�_ە�A_�ߕ� ��������k���<�E��*I}�u@�:f�?	K7^�6�����i�� `��g�����O��@1�'%�b� jZ��>�L���\��rvz$�YF�cVNPi�W ��X�	�.��3��n߾-��<q�2�!�J9;;�ӣc��w�y ��m��b�Y�����wQ�P� ����
t��u�����������(�r痎uȳ�t��}�/
Vo�P" 0w�G��1NSi���n��uB�BV�W�K7�q�Tɸ1�w�<��!ǫ�ю���@�-�X:q��%	�En�D��=��H��8,�J�U��?-f$�V��` శÛ}5^Q�qµ��T��\8�,��b�~�u뎜�zb�u��E�������e�����DI�DI7�A^�@�LC�<�֮�I��	%~���=�On��*Q|֔'m��da��H��x�
dt[-˺�:�{21���T"^s��Z9fZ;�
�K��+��צ5o�6�������-ժ.�,�0Z�mU�Zh�$z��E��	h��XJN��}��8��:��nG�N�� _�J	W�;��X�j����V-ɵ�>���스���x�JR�I\��2�ʦ��f��m)U�?���D��B	��1K)�w,���T���ē�$��8�(���q��@��d }�k:-��
���ad��\��r�����M�\ܹ���w^	��U���m�셪	�D��i�dF[L��x,�ﴻ�wj�Z�jD�RV�{�B�8�ca,��+:"�/I�vp����>HǶ*t�L�p$���"�Tم���pQ�D�J~�Re�b���	;�>�$��đ�gF��]slU�މ�r�J��<�������ڵ�����,A�ko1����\���s����E:���&��sX�����L���cs/�*UQ�$כִ�5�i��� MkZӚִ�L�_���?���`�FF� �V�W�HA���n4K%�d<Y�~X�3{x
Y)m���P2�e��������.��VZ(��C��C� �H�ï�e)��<G�]Sy"fk��D}�gҲ
� �fk�Z�Y��Vy�mQdiœ�XQ^ￔ�
Vc�������7�p�Kd�J����A��W��Av��-�U͢���숕��㴸	rY�T�krU͢Č���l; �#�2��uP����]�;V�{��{XFN�?���J�OH
�[�/j�R�~����R-D.���M�t��z����6!y����!�4��Ee������L���l��D>�Q"���{��j5�R���=b��,
��A�Ro� �����4�������6A�(��߾q������׏e���aGF�K9:>�b��!������{�P�c�%��KO���765H9����{���yZ�3 �Ǔ�m�Hl��黱�J�1��
U2E���v�%NJ���z��oܽv�J��!�5�q`L��@�u:��A�8Ȁ�����&�ф�ֵ��]?"A��0����YQET�����I�@���B����/��o����}�.��<��R�,�� 9P8(y�0Gcck�y'�������1�阫����뙂��OffL&���N��p,���9Ƽ���� �t���&�u��`n��HW"�{�ۻ�:A�|�]I��ƀ����0ǅ�]=Q 8%����_�l����*%�1v6�7���$c,��JL�e%P��}[T)G*�AZhU��D�:)^��_R�Jthx6�
���D�����H.JOF�h�EYL��F29&$k"�Z~����ѡ�z��]/�6��
������q�UmU�s7�l3�͹[��Fƣ�eU$�J���
�+]��bK�-�h7���ɂ�nF��|a��e���$I�ju\���5���C5�P���\����۱+�Z�[^��	�%�Y+x��-gXY�.��_��fE:�T(�C�d�����k��ʶD��0�A7�U�'5�}I�X�:|}IQ1�/U������[a��I�Fd��T%z��>�zm�j�-<���+V�˪�#�SB% �}�~vn�KU��;:�H"�n�����7�D�� ��6	W
N�����5�G��@d�����3�Rj.�x��g��>4���FX�1�+*�4Z~��-��'!���J(ɘ�Ң� H�V+pנ��5�؃�����h��9[P�a�A}:O�5������ʪ۪sij��j [���A�՛�P�&u�)ET],6��z-E>��P���#�a�j��ZறCU�eIp�)�����>\�0A~�����ԻLe Ú���`���tח(	�9MkZӚִ�]k��5�iMk�w���.�0���=�-,P�?P�j���J����:��Sa�:t �xO��l���OhU`༙{3+#	��T�c�� ��sB��*SSmT굼�
�##�� ��>(�U&��D�ګ�J��(K��J< $bn�[ӫ��o>��[� SB�e�e�lb��	%�qV
jT;��|A�N�jR�VC����d:�MNm}����fDf��=�k0~�UQ���'����0	�F���
�^���P��K�5n[�V��dXt����\����� `T(>��n 3��di�z>�B����:�������Z
]
��q5�$xH�! USҹRS��pl���2T/�@e9�(�J�ňLi�:Vj����39;>���M�'�$�%;����D��o AP��,Z�Vi�#�?��cHu��H~q��$pڑ$��vQtM�9��� ��߿'����E��� �OΎi1�79T
�J�XX�ۡU��&��r���9�G'2wǎZv�{�Lf�Zg�h�Qi�G����.k=�yk���̍չ[c����-�vG擱,��/J8��:�ר!�i\�s���}i']9?~/o߾���n�QP� �C�s������f�Jƾ�۪�
0)�B�NO囯��?������7��w�����?�'�>S���d�}���ٹ��.9wq���ȍkS6�01�p~N]���i�y��,X��>���'���s�HTq\�f��v�qOC�+��X��A����\*P��`cU��� ��������@�����_��R��ş���P��?y��J@d:�����9�3iP��U�-l�޽õ��#�=�M�?�b�ь�������sȋ�,�riwB楄�U�����-�� ��P`pr�͝��W
ƫr*��ހ�w܊i�W�z-�DY�����^⊖��@����֖��'?���/���}�����V�yM!������B�pJk6.�P	����Ol�ma�L"wޡ������`��Y1;��8���Mkw��µ����*���F��h��q�:7���-��bi��]�E>Kˀu_@�s)��?�B�3��H��O��Tz��˕�� c}�ȇ���y���9z�ӿ�;�-�yb
-��5��MqiVt��إf��_�L�MyQ[e�mj&��6��?��+�����y*u>Ida�uk�%(<�� �\�V�����2�ߋe>��cO��_���4[����2����*-�g����m�Js�*޷��Zn��S�b����
C%�Ř!�jN�#H�T/��7��4fELI+=O��sWN�(-|ƌ�'�Ŕ/D��b9�}^{�!EO���5w�ۢ��3^Gw6wi�W�>�B�gX���B-�y���� �O����grx���|�1��Y����͕%n���C���nKɡ<�U$���ﶻ�L�/�v��Ν�T�17�ժ� ����y��6��Աf��98:;sǾ�yO�Z4���*��j�'.�Ul� �ZRR�Ui�� ��x��7
n�ִ�5�iߟ� MkZӚִ�LCPq'�HԱ�Z�`s9ӯ`	 9X� �`<��CU[�^.'S��Z��{1�7p��L�^�%pP��ªj�8,5��>�H \a�T�a�F~L�Z?� r��R9��[�0VV H6�_1�n��Z���g�{@F쎡�v�+I�0�����+�W�܃�8˺
�����,���Ň�2q����Z	��%ǣX�:Xw��Y�ya�K��%�`�������%	��ӊQ�Y2IQ�R���ՠא��ڸ���4k ")R��Aj�<@+���gu7"�(Q��ٱd�ܬ���֥���-n�3)�y�����ϼ�:�+�Yň*� W���;����-�l��.����#�� 1�Jw ���BV�p}�ͧ�\\����
�� n�mUr~y!��Gf?���sǅ@�n�}*5.Fg�ܼ}��9�g=}��$B�Jq��Z�ܔ*��J&�)���o��|�  ukc(��T�>}J���DA�
�s�����{M�!�Y[�{�;�}���wr~1b�:AD��m�9-�������BF�rvr*�m�q�\\�ɥ��t:e�y�c������{�k���Mǐ"&ry:���-����3���|2��L=�G�	��67;�Uo���>O�kC7���y[ЮD�>d� ���R~���ȿ��WTD`~?�\��}�P����)wD�����)���l�q1wc�)D��#���P�1���o�~#Sw����Ky������>��4������Tt����M���4B���V��p����;���;��ǲ�r/��"Q���d<�Z��ȍ�o�~"��<y�D^�~��Ñܾ}K�]�����u�,���L���y ���pc,��d>�ŋg��?�ٍ�Н�r�}a��Do'j���t6�~���Ĺu4ss	�e��)Z�������y%��*t���1P��v�8 ��Ү(P�K2��-�<��~����/���0�q�i��V����۷妛����`�%(��'rv|&�3lnqA]��EqNВ63,h3��; Ū�CJ��/����>�c�
���T���?�s|$�{ Y� ���$K��eSs'�����1x���;3�0�aj����Tw�Z1��.kE|[�8�e�$;X��.�z�=��$Ѻ8���F�* �b��,�Dr�a���+6?E��1�۱V���%�]�����Zs�*�J*	��ŭAT).������7k�W�+|H���Ѳ�?Dv��/ig�mD�#�tX�Ơ`~��+��ZNK4=7�n�ʆ�����|�eh��
�Bj+(Zs�~��VKF�c�@j��/�a���Y ��l��)��w}�B�j'���Nz�q��u/��Aڱ)NB�ʖ�AnJQ1��PIa�V�Q��x��G*_|XK�Tɀԛ�s�R���ڻ9��~�_��?�/$�aa8���2(fk��c}mC���s��#������{������V>��s��S^��8���=�
ē�?v�q�gve��L�ǂ�a���	�Mp8w���V��`g{�ו�u��H����A�*2����z����?�T���������שnWU@>��p���R}cj��p�k,��������µ��jZӚִ�wk��5�iMk�w���f0t��\�=`���P��v����C]�����{`���=9����������%G^ r%R���	��^&7�(< 1�1jK��#P�u p ����ߧ��Vq����C�$�(��I�e ���(�������j%$�6�UxxN�`9˙e��Q��`A�@V�,�i�y-⟟��\),1���!����W}w��>`��*UT�H�N��d������u���H����VaΊ=�j�zH��v'��<�+l\PM�>g�+���d�6��|���X�p��^�+�  Dzu����\�L��c�?'mV1�D�W�0�V
�퐫X5w; ��
՗9��CE�W�+�L� aS�E�����<�l�v�;���:����
�"�%<7���</����N��=ܭ�w��g?���s�=�ywȹ���-��Ab ���#M���V&KV"g���h	d�P[���_�s̋���k+�˥�]��A������\f ����ѡ<{����A�����Lt;&���\�4l���| �����Y+(
�O��T:��VT��X#I���B�����Ƨ 	6�������2Cت;�6���C��w}
��{�%����Lf#�g�>�����@��@!2}J��3��ȡa�\���@�g���z����_����7�q?�����\8;<��/]�����o궽���\\�H
�}Ϟ?'@��7&���w�F�ݗ�[O�1eU��p��/�̍�k�;$ϐ����Sy��lm��ݻw�E�9����?�{wo��%_~�LGSٽ~]nߺ�q�5r��������_ݸ�dv��
@h�!���s���+7nܔ���K�?���.O�}Jn�*��?�'�w��~�#��n�������ܿ�NH��2l����I���[o[r��=f�����>g��h>�s��J��8>�ŵܘ��3��W�F�-��)�_�< �5�s~B���$(����,E���8���eX����v���L^�z	d+I��Ʉ
��t,�p]B7���6�ѣȿo���y�2%A����?��Ė'1��~oMÐ��󾢂%��͢ q��� �TXぬ|��W���Dvo����.	U��]w�F�y�v�m�DC�SU�`.��ֆ=� zf�+��퐠$@���`�փ)��E]�W~D.�;��[�@Ҡ�`1��E�9�u�~23\}%��@�6�-+DH9Npw��G>����.j�dA�J({Hd���K"��R5�������ü����W��t�����%�痒Öhy��ɆV�U�EZ�1j]V�F���V��ad������+�!Z �r׫�d���'��/Y�OVP2��#��T���qKK��
W¹WO,�����BK8-�`F��'�70��:�~����n��23�JUh����q*U%���켔��˽mh	"3�q�,H��(L0U������^���qwl��������9F��ۚ�u+�4�;��l��I
�w����������}�[�_��Xwql���0Ϡ���mTTJ�n_ەG?x$�;[��x�j߭�)�z�̴����'�Қtt�ѭ3q��{i�)q�
��{9�iI�b`�޵=�q�{�;w��g�}V[.���f�	���]@!㮥?�����G���w�>�� O�>�ӓSy�~BjǙ�I�,7�tH���U���\���j��ґ�§��r��5�iMk���5HӚִ�5�;�� �0��5d��l�� h ����A=Q5	��� p`Y��Ks`1���R-��Bɏ4-�����ļ���Uu�Zn���r�B+��0p�Q���5ϣb~H�� 6�U�,5(>����_�r�U��������2VB���k�m�;��RA����������
�x�u�f@
�"0[,˶P;���ȕcY�I��Ci��j�����a	
`�N��T�`�b�Ň]��U׹�C
1k�*�P̒� *��}��T�т�+�*ǱguȺڜ( ���juSք�o�[@%���XB�1��0�l+o١�q�/�VO��jB�^u;��P筻��F:�������;����//�=�C ��2K�4��9��J�;DUV���];N���	��2���� p����,�*�ן|���O�|/_=�w 1.�X�=O��rİ[��A��cڃm��Ko8t�fH ��ߥVQc�Ȱ !1�NI>���v���"#`��K���G�8>>���|,wn��*d,X=����BƮO�*ps9��G��lF���eJ��ڰB��%2�+Ӵ���1��V�な���vc����֓ȍ��7�y�`W�� �_���$��I�'����h,��$@ ���K��?����C��m�v}���NZ�i����=y��|���<U���i���i.'�����O	2�P)}����N�Z���_H�~�+9w߻�!�0���ߋɥZ��XBX���b� 0�(l)����ݘxE"�ݻy�~ƶ��yG1<����˫��叿���q�<��`~`󹂥�;_P��ܹ��|4��|�Ώ��/S7G.���H~��y��7\81^:�᷏u���Q1�ZH�.h�kJ�uh<���R�բ���e��;�yU�)�z��_�s,	�D�;U-s���֒��C*�0�A,x�L�����^��)2�$"a�?~�;y���Sj��,^�HL)�a���\�r�\�0�g��ߙ�E`��-��ݗ�p�J�Kx���n|N"m�y���)`["YT��ATښ�,s��������W�)4��yᎁ��O(&𺮝G��2� �b�����bJ�:\u�����I|&u������#�eU�\sQyN�|��3P�ۚ�@>(�ܹD>�>�ksG�nL�o
7�ٌ��1���'�_	͊���*O�k��*	����L�Q�*9]�N�V��t�ܸD�T�,�1rE�rU���AW�|�ϊ�(ȇЭ�<F_H��l���k�(�j�IK9�8�(j_���:��2��ᔥ��&�ܠ2�MgTp�F ;�q`!�)��4oN�S�m� �U+~�G����3T0�A������P�ݽk���D�p-w�u�R�nxx� X��)��~�������C�s��f��t2��xOK�Oj����=I,-,*L�"��ԹZ�F�.����8�{ݗ��?��۷dǭUׯ��I�I�B��!�=������lo�4!
U��^�=�Y_�7����D
7ǰ֣?p�x�b1�X�f�ǻ>	zRJN㾳[�\׃(���@�ִ�5�{��iMkZӚ��i�TD`�1U����Rw4T����o��@�x0���� *�T�\#eT�������>��]Z��, V܃ᄕ��t%d3R�ZeQ��dQ���jxB��\m�����2sE�C�6W��u�2u�=� ��p�E�x�sU���n��;�[��<��g�w��Q)5�j���T� �,cVSG�������U�b����y��@^ܯ$��kV����$��~P�Q?�U��sP��FaE�{P[��jhȯe�!|X�!42H_���C�����<��_����d%�|�f��*M� f͜		&�f�f
XU����o9�c���$ܾ�{҂}IH@U���OeogW^�J^�|�
z�{�8L���\�Y�	p�C:_��w>��l1'к��&�- p<v��y8�k��p�Ϳ-�u���.��e �}zzL����9>�\<�ؑŁ��u_�[�dE�0�ma�'�3s_
}��
�x��=I��E{#�zl����ũ�fSV�B�%m9��
e�P��4��uXͩ����X�(��I[�`���1�/z<oۮ��k�rmo��`rYE2�ؑ��XON�_~�K��'�Wؔ�Frp�gI˶TN�i9�>\#����.&���;�󟿐�o���/���W2vk�,�8�������-���@ܹsG~�_�\�h@�c�����X� V����;� �s�:F�	_�-������o���b��m�#�pF>�G�h|!��g������1�sy6O������oIpc��[=��nlv��^��5V'_��;o�$Ґ�r�ι�
腜P�-H8�7�ƭ;�ɧ? q�$0,��~���������Y�9��U��CU7d�^��-Z�����L�_�D�:[�05Iw����7 1#H}88	����8y��[ۙ��`Mq����[y��
���>����<���?�	�����G������D���I��J�C�@�b�0�v�6Aм��$��ہ1��ݻ�d��-Ys������]cy������F~���<�c�-D��a��dp%�~O��S	u�Ď��,TM�"XK3s
��*�p�!�)��E���\s�
U�$��B�`6Dz�f�6�����0�}.�?�nk�Oa���'���C�k�P8��j��9.��{|�7��������;��Aq���h AZ�����F���C�[
Z��Y%A�ȉ+����,b��(�j�'_�6(��-�ڪ����'?���j 5IǕl �ٜǼ��u*�k�!W�%Jf��!�� =GA�ٜ��hc%�7��$���J?�%���,| 	��*���J��l�B�bn�Œ��l�y��j)�d�[+h�ǆ�,�	�Nq��z��w�޲�í��Z��ޯ�x��-��Ӽ� 	j��?���FM'ӕ�[*��a��	MsU�!�+0�CY���+�)"�� m�ӟʽ�y}H�~��� 8y��9�*|}�3��Z�����-�oސ��<��
 �-����Q��=��Ѫ�ɩ��l&s��b����.
w�F��Դ�5�iM�~�� iZӚִ�}gZ��
-b5$+�E������ XՒ��6>�U� �!���Y���d:��P& <i5ѭ�W�z������!8�=���Q>G m�*����Ls4�/��\	^����YjwuE�!+��ڞ���H��65p[��3��-��K�`����$i�2�}����C}�]j�cfV���"|��S�e>��u+D���*D2�$�����/s@����WM,>�B�Cr�`E��,�px< K���V� 3?��`52l`�{�`��	 ��9L����(�~VSah11)�o�G�����c�U��H�bP`Ы:�m"���� �\֤	S�()L: ^P��m��P�yq�q쯭��s��k���w�ߓх��BB�ٜD�XX��� }��$)4[�����M"4#S���{ݶ�= zA���]2xYm�0�W~�sF�1��W XJ7�X�����p���DU&l�〜�r����#*A�3��%8V�?ݺ}GƓ�[G�ֿ)�y�}�\N���||,q�'����@�lnKV�2t�";��m�5Hv����a�w�y]3B r���s���%�;�2p�H��;�R��5y����}w,[�w?�O	$��w3���dl�擩��IA�g�/̝��k�'G�f��ܑ��k���+?�я�ѧ�������~����<G�>H#آ!�a:�ur�>�~�\N���_Y�ɬ*)�t/_����S�~���������5~.�L4�2��&	�
೓sy���wt�흻�y�Rf'n��T��sww�s���*�N�yv�=w�})���c7nf/X�`�ιFA�6\G���ܻ�@�߾+}&[ۻJX�;�����6[�љ$њZS�5	v���8 ��ͥ���ԇ:g�sN[��^��Fb�n��+�m=�ގښad���\�@�P�wޟ�x.{_~I�����}��Lr���[�w�k�����L&�\���)�L�-�ƣI}��)e�{wl�Ì�v��oݾ)����(?������=�k	�9���ʭϞ=�/�������m�^�}A��X�9?Uҍ�u)��B��/��X�+S���0�|�VD�2�:�q�o�����o��P��K �ܑ���Ԡf��Ɲ�y���^�L��:Ƌ:|�ҋ�\K��6_h���P�1�9i�ܵw;�8��,
�. W�-��z\��R�4�+�E.�,�4�C��ֵH#Z��_��H�ug���͓�ׂkcl�2yiDH�����cQ�k�����]U�p3�Q/�*3&	/�J�$P�[g9p�I�z��(�z�q�pO�\g��{���bYd��N���i���^�CT��+b�9.�	~ͻ)���5�I����L٫
�d�2�jIx��e]� sI�V�{\+�o`����3\A�`'�$�q� ;��G��,��������R~`E�����<0w�5qss]��R%�����ӏ�⹫hgXa�W�Fa����ju}c]666H|��F;D�����~������I��_\�0�@��9U�^ԐMkZӚ��mҴ�5�iM�N���%�_�F�u�#���A��yfvcxPY	�VJ�@ޔ�x�^ܢ$���]Q9@��L+�=�VB��6�`�x{�p	���	\�P��	��b�A�D^J]=�K�L`��[��@Q�%�������4	�t�uCa�I��{���ן*��p��=�Z�.S}K*a�!�*�4�}����]K�g/�:�!��]������8n3���vH<Ó4z�
P�&�~/��\ڂEU��WXDXqY)�BK�"W�+�xGSm+k��ո���@�!��G8wA�R��$9�4���5x��!�@���� �Du�F0�R����Pmz%��lGRP}-�ٍ���A>�Gmx�=�C����;2� 9�O�ϰR�~B�<�3�nܒ��-�� 'X	�:hX(@���@VDf�
����; N@<������t�l�e��<-ԫ�R0X�+Ð�:!����@�XX9*��nN�`�W{��5��!�iu%�癿>:���hx@��,� n��4p���W��rf�ܹs_�n�89xC" 
�mol��ε�p�	N�v�Cz{,�PЈ̃�l��(J���k�Hs}�hmsGnܼ+���>�9n}B8��ryqI5�-��8���K9;;W{�4#�srz"Qǭ����\��>��}���[��H���@�9�����ɤ��9N`AB�����
Z�U���|��W$���J�<�eX�u�C�}�����?��-ؔ��_����s��AJ��wn?��~��s�Oy�����|��K��1�%���|�_GG$��ތ.'<fӤ�a=Si.T�j�.h{sSܿ/�~�Cy��ZBay[�ؤ���7�_ʟ��R���+0+=Uj�=o�o���F?�d�w����)Q��~T��H��MU��,�Q[�ehyU����*��|nP)�g�n�|�k!p�7n����Ǵ=�=<�Ar}�ŗ���s9>:T{�W �]�^�����H JY�L��ts-u�;��ݐ����~�y��C7�:n���vL����k�k0�AY0�#4�>v�/1��Ӻn���X�v>j��,50�E٭+�I`#�˭ ����TX�5ס���6A Um�Ut�ڭ���1��5Utj��@�������W�3�n���%J�V�+�	�;V2MĲ�
�A��:r��:�\���k��Bǭ��괻nݸ���k��-�w�>U� t�U�c�˸6�݂�)%����aM�����\yŇ�I�;��Z���Ռ���R]��!^�ado?j�F���g��s�[5d>�>.C�c�˾)rS��F�,��Q�X<��MA[�ފ2�06@|c@�C�i�ׅ(�[�P���� �%r�*�ZT�F�
�c$.$5)uӯe�)��	���闣s�N���b�[V��C�
#��7�$!g+������EF�2<r�?� ya*�@��2�{[;�)��x�x���9<_��Um�௭���{�6�o��r6�����)5��T|�-o�J�T�����|FR�0��@La�)�:��t�h$R�,�Xhҝ+fnӒy�=�)��Ѵ�5�i��� MkZӚִ�dK�3����4 !�ł���V�%�%�6�#��v�����{���b4�<(5���Y�**%�� �0{���� p�I��hO��mBK�V�Uެ��Zi�� ���}fz�s8�?��-�G�� �T9�g�� �8ҿŦ8H�>���c���v 4J���W��]^�p�=B�<`���{�0���,T�¢)�_r#��\��jǐ�JQ�Z�0��έᇜ���JV�B��=
�r�և�@*�w�3�/�W�>X�����[Q�T��s��EYW%��N0��ցz�W9)vV���M�2��8���,y^���yȣ��\� �O������]%�jr��� %d�P�6?_�&U��������0�	���l��KX��f�T�����}�q�~�\c�=8��EOv�m�'����ߦ��m��!}�=����A��j7� 8��;9N���s2Q��%�@�)�<���=x@?5 Oʌ��ط9n{�<��8��Ȼ7����['H@;B�����i�U�ҎUq&���Z8������������������S�r��]nl�r�������k�K�I����>=�w�yA�@!�]R��t��GX�����ݑͭ�?d�[䫎�Z'%Y
�܏��lA�T�E�<������_~�̉��s����7e���>����jS�s[�P��"���a�8���u��X�`k������:�����$���/t�}���u�;E���d !�@�no ]����أR��͛r��=�w�up�_j�=��N��������ג�!�.��t��r~"̜�!�U��sO�&P1�\�[�d�a��R��Y��	c��X�hͺIjˤ��κjꚢ�j����" �^���'X�A-�,Ãܻ~Sn���~�<�T^<{N����2�̸~3�k���k�2*�B�ȿ��ƶ�=��s���'��O���;�o�� X�' Q&n�<y�D���K9t��2��Pf��r+B��!4K#5G�3�èLIh�F�$���P���&2���j�9D��\������j�\���őYz�*\��h!#+�k�MPp������� X^���Q���H�+��$�(�maw�!OA�m�����1�Z�F��ݼFp�YW���f�ԖV^��Z�Pџ4�op����n��eg%j㤊�Ю�W@3�y ��^m#��%%S�M�*?Af]+�+׸������"�氷���c��Hm����re��g�Z<r�
T=���d�O������R��Yi�Ha(�8��H�Zb}Z���2�Px�.�{��ͯ/X�y�mPI���5Xù�W�嚭����{��Ś����/嫯����#�t�թU�!����CQD����l͕K���b%��
*̈́�	�/�~D;x�ֵ���F�;PK�^�0��XEA��nIKNd"������[�3�k�wnq]��")
�!�zN;���!a*Yi��U��e�-MkZӚִ�Ek��5�iMk�w������߅�V����|*��}�ֶ'!+�3�  @?�P���`�����Q��1� �"x8Mi���vN �PF����	����; H �E[&�ɒ$����i����ros���A5�&ׇ�$@��N�m�ڝ@�'&D�xƇtm)TQ����Hh�DAU����I e�ڠ�Qѝy�@�9U<��tb���F�jN�2]�re� h<8���62F�">�4�q��H�8h>|� �$�vVV�,FL��uF�sa 9����?o ( h��X̖L��Zu �ƣ}nVWP�t���H��X|���`�rQ\Q@���/�6W��l�̞�l���a\*aR�-
�⤫�!��Ls�-z:�뗯Ԓig���(�b����G z���!�6Nn��s}��K��4+f����W{0��gf��	>��p�0��
s���@�f��'#U��Ah���xT����	p�XV�B)b}J���D��JH�,����d��]�׭�<��@���#	������W�UT��	�J1�Z�h$+T�@���v�"(��#oFx8	/^���͟l>�e�H�L��xɱ�M�7��퐸j�y�궩����~Fo���-��,n%�}fG�_0k��kݐ[B�Օ�چY�d$��w�������sV	c]ػvK<�X67vd�>pǕpȆ��`
�Ia�3h�<�:����*���]����v_��ꉼ~���\�:�HD��������������{pWvn�ʭ;�Iz\��UTG�Đ���Ie��o�ȟ?��|�?�1�;�6��G��,�f��4�g��F%6BʑI��Z�mQm��9o���G�L0XS���n#���>V�
D��
I(�=�G��%_�L�b����7oߐp���
�6q��Ļ=�vݍ��C���*z�w�紲�Zs���;��ǻ1�Z�p��);�}����_[���k�{�Ab������J��n_�����o~#o���l:g���ݼ(�ŵHI�cgn�R�@�R�>����u�����{�<4ā�$����׮N�9�EO�B����.��T\3I��
�C������*�#Q����_]���xkJ�s� �?��y�'Ǵ6�6{��$,aI�QEMDT
*y�p����V��7�Ϝ�Xc���1=E���+d�X��������GFGD���ʹ�YFR�j�:��J�m��]y�I�WHlӳ�eX�ǢR�2�|N��*�՞Vq�Jq�<�WT�^����+��rI�| �q�[#2Uo��@��x��%4�HT�����sL���Z���q�AVM���'jO�=⻷��7��y��=U�m�ֹs��k��D��&!��:�E|2%,�쵛��n���P��c�}��}��=�jx�����z܃�u����t�/�n���ۺ8�t�"��˿|�j���G"�Oa�5�P��g�̊>�ʔ-z�@�DDm]������{y��>A�9$(��=��|\c}�j1��oМ3zO�>1��5�iMk���5HӚִ�5�;�2�t���m�z���e!��ʷӳS>`���� pQeJ4%(I��pE�V-���������|QҪ�vV�8%v�)�j�(@�vG�4@�-�DK��j���)k%���r�V��q�uhh��Xz�ke1�B�,�����`�� !p��  �@h����	`kN3�ya7$�A��*��@�L��������2�P�
�v��Ӭ�#���L�Po�T�Xj��<34���+��R[3{�Vh���;(�`a�L�d������kH.��=@�������fՀm� �}��t��A�Ɖ��$I��B3@p\ Ba7�  OI����泩�9��em 1�����\gx90��T�{8VX��`eh��C��4H��L��)K��2}�q%js�J��`7+���-
�D��dx��� �pL3w.0V��X�u6�Ӡ�(s��P2C�죥���LпM�� ��2b#�ud�>.�.��v���Զr�w��a��n�y%��ků?�-UVg�DI(��Ľ��}ë0ΰ��B�u�.A�7o�˗��������~rr�ֲSX;P��w��ܺq[vv�d���>�v�ܺsSm�H��U	��g K���[�J��u^�,]����z�C@Vf���[w�]7���e{o�}�ܑA��I��I�sTc��=�k�Gds0HM1x� 82Azn��.�Y��u�~�;�y�j��M�yۻ׸�k�*P�L�7�/���>��S��~ත�,�U��I�t�1A����o����o��������\�7vd1������#7>Oݱ(Q�e�Z�P�����:�C�& C�%F��5&�N�b�*%Z���
�c��i��O�;�u�S��=���T=F2���M��
k1T07]?D����ڍ���/w����wܺ��~���;>9��C�B���:��#\��Oe}s�*�	8T�Sw.w=�L�܏���'�>q�m�`),��m�C�:�������l#��X�Ś� 
�Te�S^�GKG7~ �����X����i#t����Q����Y�-��X^��`���/�WT���$�Kd����O�ׯ�Su��������N�md��y�r��T�N�y}��HצԭWJT���zE��ef��Ӣ�R��D��6j��j�(���e��W�z`Y�W�m(}N��;�PV�A�Z\�/��W��X*B�������aIzE���E���W���`BB�O��oIM��ﻠVAnh��F�*M�ͷ��~�=Z�J@�A1b���Ŵ�R)�?T��Qȑ�#k	}IP��QGY��Ԉ�(Z��������S99:Ѭ�|��Ҷ[�7���l���~��Z����	�Zf��Y:�|���b�\$�_�!�bvx���1�r�-���{�K:�ђ
E:�gg���e��#�:�`5�wMzkCw_җk��I��7�L�5k>����Sy����.F����[�9=����v�d��,W�Ͱ��Vnki~e�T̏R�X��5*P�z��k�+��ִ�5�i߷� MkZӚִ�lYI� *�hR�K�2�X��=h.�� �����Fu�*���/�� �$M���HX�����B-�B�㚀X�;	a��e�}�!�%s�B���� �2pn·�9��@ᑦ
���s ET����=�Ā�؀�J螂�(�}�S �"���m��#�O}�]�QY�JI�������a�Vo#�˜��8Foͥ�����>�#�
�H��v����f� �QrJU2��3��̫JU.d9�? j�f�	�Q�>��;�A���R�WX�fb �|u����{k*YJ|Vy�$��}��$�ǅ�,���#������ "Y�A��P�kE�۾�a X�p!g@�4[v:������)�
!Г��ܿo޸!7�=ZD �D`����B�(����̓��k)���}co��5@g9��[��B*@�@]���g P<؈mԪ�V���FZ��
 j|x|ld�7�Im�dL�a�-$���*����M���q��/q��q�*OT�K�j��M�6��ӽہ�FE`;� kS8Q!��X"S�(��ӺfA���~���8x]���'��@���Xf�[�F���y�N}���[ ��ܔ;7�<�u��g��z�I%"�n GfϠ7�9������Y)��X�+�b��/ +U��m\���Ms��@y���7�s2Z�"���rK��۷�����V�M�% 퍭�
��7n��O����@Uj��I@��bkc[6�7ꧦ"�ڂ��qk�B^?.O��Z>��免Q�K��9\��\�2�ҝ�x����VV�
}���$O�BRPq�uk&tP���q>[pQ�R&i+�6r��,�;���0G@l�n�:��T��{�V̧�1�J��B�� ���_��<}�B��'?�I���=�/C�P������r��M����hUe�;g��g�*���\�Md��X�#3l0?�
f<g�~��1�������ǿʟ��'��/q�_�z}Y0s� �e���}�eT�^�0��n��(�����\�2E=���uU:�K�J��A�r����oN;�P��H)�R1Rrd�����Q=N���µ�NJ�`8�Ȥ���0\�hSY��^�5�׃Rm7K�FJ�_^���E�[�_x�L���(fv
N!��EJ�@����F[2Xz�w��ކ2���Bcl.�3UǸ�]���|r�\s|��	� ?�����r�jL1�-\o�Ԭ#�Nч���.\��7`�T<��]��X�����Fj�WˬE���'�K��5�ψJ�r%�g5�G?7�l�Mj�Vf�Ofq\�~`��`+J�اY�ڵ��Ƌ��Z,��)�8L����P�X(����9@�f��?�n|��~ >�X���*k�I ���L�5)����L2X|��I""�V*���JSָ}�=
σ�X�"��B��%A�;����v�
Sw��ҹ���9=9%��vk>�? �qz�����?˝�]�;�0.�:��M��o��_���rp�N.ݚwq~��w!�)��}��ٜw�o�}��]+����RO)m�L�J���;MkZӚִ�gk��5�iMk�w�����H��B`�{ ��C�cx���N�m�b�L!؊_(c ��7pXDT<�Rݡ��m� ��!��B�I��!N
��a�Y���$�]J�`K��˭��Ղ����Z}����Ҩ,���A��d��T���h�������dȅPi�ڈCYVA��~�/4xݲ3|���Z����aW�j�P	!�k�
�j	g���'���"��x
|({^�$^��MLm�RiX;���@x�!�8oUfʌ�0�B�jX���Q
�
��AQ�5��J1?�J	�ȫa���_1��CB'!��O|%g�� ���ϗ^��dQ�f`�P����V�yJ jV������3z�s;n��y}���q�柴U�$���z���c� K!�9�u@n�|2�|�
��$��tƐk((�g�*C�L ��ְ�Un|+Q��aa��2,��X��ݠ]Y�*z�/�b�n;3P�?5�U�^Ɂg�x��š��"Șk��
�A���aH܉�"��o�|�L#��f�㶅���ٗ����aQ���7��:�.�پ~M|2a?�~���2d�����������Of3�j ��@�=�>� [ v$�\"�#0�ɟ\-Ђ���]�N�S�+��k� �>�#���|6��R����,��Y+a��*�a����E�	��i����9�:�[<���, �ПX�a����S��w���~�;f���<��X�n�M9<>&���ZPR������&P�i�>��c����Ę��� S������,�G�}�����O@������J�ֶJUU��(T7~�g��g�"�)��r4�OOO�ѣG$<��J�����'Ȕ���T�n�ػy��*�+ �õy�\����h[���Ir~r������׿��%�>}�,�d�@����p> �dG��=���S���2cii�s� y�~�2%.��Cz޳�7���g5�^笂�*�<��kB�s=��+Ub$��h^�zS�W^	@絍y`a}m���^1U�9�¹�c���_����
�"�灠ӂ��� � .s Z�
�ե�  �p^���T�� ���k���+2����0��2�+��a��[�.��)�ڔ�������Ԉ�%b,�\�	M}� ������XC��+�.��^�1$�j{0����#ԟ����粸B�nx�c��"*<�\2-�hܮk�*�"s�"]�[��c�����^k�]�4��\� �,��en��!�g:���ߩ'>Vȁ"]�d�{䇒�lZ�{�] ��A�
�t��Um�h�vxrĿ������ۼo��Z������ݻ��}�۷�Z��̽P6�׹ ���/{o�,9r&�@.g���H�qh�4Z��M2�����Lcv�Ff3�{Msg�d���Vwm��%�p�� �{F�}��b�ɓ���s�I�AP���R�����o��b�m�l���ֶ����g�Vdmk[�����i�Іj��J'e=��� +��>?��&S��+��A���m8������ �4��;�Q��FVu�͑U|�`B_�^�� ��QՃ��K���$Sd�0�>u�,Ǉ�/��R�ح,�z�P��̏a*�겅����X����4����ANw"��E�й 6��|�i��ú� P"?�d� 3�<�RQ����4�������-h2�t0
p{��4a�vݔ'Ij���>���&(G���l��*�����Q��S%��6"FR��@6HVu'2R�^�o��;)���ű����k�|$�K��j�]Q'�Xy���H�9�ܷ-\U�cL�J��������}��~ɐj����ͯIR`�����믾1�7XN�x��� ��X����C���Հ�U�I�}^~�=���wT�����k � ���޽��c� ��~s����)qZW�����i��օ ٙ6L��A�hw����{eĉA�s��V$�T�B�$�R]N� X,�ة� �WAj�^�`3r��D.���U��B��[�Đ��o�?�ro�d��X�h%E�al]�,'�_&� <�����?�1��o�3���_�\G#w|�mn��f`��מ��J<W�M�w��C  �����ZX�t�߰�����~v'٫`ۭi��xk�ݳ<�no��T���
���;��8ϡ|���7�;�k��;J����J?x���������������=����~��7T@<����(����C�Ab���VcM��䎩�I��$[�ɖ�D��&+��8�����F��*��י|M�j�-3���y�5; ��t�$��
�T���H�߽{˿��	���o��>ǜ�<�E�-��tV��$��vu����O�n�������}x��5�ا�C�����/����s���� �IW�V�3��T"4��Z��DH;9AH={�z������X�
$��+E���Z�+a-Г�Ő��g2�6Ub�u��H�X �T�������*]��~�I}�����g��֋f�xs�#�F�_�+��Fiͱ�� �=�l��4�[�t@�R'�O(�蚖���ڠ%q�@��]T?�j�`��62끇���GHf/-W!�5 n�i] 2=�g�F�g�,�E���Yc����w[��U����$�hU�fw*+���s�%s�����M7�N��_�h@$sg���r��G�Ԛ�sU���x��
2����;�SJfI����Mq�,+_m��vZ�.c��s�״E�̲�uݽ�yf�f��ndHz2�8�}'F�,�"���@�@E���w�|��{��(8�{�*ρ����TO�s�2�Z#%Q�EFm��0u��t�����P���Ԯ�6aM�}}U��umk[�����l+����mmk�I6Tk��~������uآ"�J�exs? c�F~/XA�\�C>���tf�;�Y��ܨJC4�4p>���+������E���5>x�$Q�w%��}�	Z6 ك��(i�xf�3�yM��i�ZV^�J����hJ��Aݲ1zUǎv���f[�s����j�h�Uh�w���L�=�^:�\�]��T~�L�P�%'>�R�Y�,BKU����,%q(��J���3��� �N.K���#�G �*e�K-�-�Y���:df8���JWMe'���$2�?H�����d�"���Qi\Uٸ`�T
Ce��(p;V��v����+���r�2_��������|>����W_}�����7m��/EP|��6:��n�)������;�P�܄��{|o�>dE����՚�u�����}�vGP9�c|�ͷ� H>t�=@`LA��޼{�[����M�‖GgY
����*~ ��y�`����1 }��ႪR�(V yd�?�����q[ g<gU��'�Ҝ����6���sv?�}��LE�D�S8.d� �����aow�k�`WU��� ����9m�>��n7��'��N
BƱ�&��#l|&��ؽ0K�
6F�������������˗��o~������g�I��� ٘�N��	+�o�%H���v�����}�Ͽ~�6O�R�7ʽ���\�����-�r&N����pL7�m��C?���������7�[�d��:��H��m��Z1E5�[�y��g�����u�|��>����)��O p�Y�������W��#��W��|�-ה�w�h_Ek&�)�r2�ݘ=��m T>�T��
B � ��Я@���Δ
�=�kX�3C06h�ǹ,�U���A�B1������d�+\˾��e����7_������oï���7�7�W��C�k�_"h��Ӡ�`Z�A�RI�R$�_~I;�W߽��>��o��q-������c���R�B��P"<�kʟ�Fc���3Ǽ�In�>�4l[멾�<�-!!�=���_�py���Z
{7�I|�Bs*�:I�NjX<&��r�fEd2J4��X;�9R�I)H*�:M[�U쵯F�7�1[+fush����c�l7�d{E�I�]7�@r2�YX6N3iΧ}�ZA��T����|���3��j) �8�Q$Q����B���z����(���T5������^����������F����d�ı�Rp,�e�����k�5�%�IHL���N���b>�y}ߐ���U;���e��o'?~��t�FA$+2A�I�4Y��R�b�`�����P3�}>�:��J#[4'̖J�ٲ��(��ujl]F�2�sI�.�K����㮸d�H���>k+�C�v�p��"s�y�ۙ̚R�Y!X�Ii����S]���3Ҳ�DH+.���Տ۵�mmk[��m%@ֶ���mm?�f�	�=�z���r �Fvu�̈�U�,��u��[{��0�1�V�_) �J����X,�X�j
�jT zM�-ث4������Q��?����  �Uq�U��Uzfsb�����طi���r�i��Ce�Ĉ>L��خ�N��A$X	$YP���CU4F�|Ά���~�|U�I�0��.�N��R�ܑR�j�a�D5��x�S)R�&KY��cQ��ÿȤ��L��AB�\���Ԫ�É��� %Wcxȵ@Jo��Ǉ�:���3��i���堽[P�2�����Y-�#��M�� C�����jz�hƹT5tE�������!�?��d�T 0�!|��g��/>�1 �]�ƛ���D��#����@Z�b��,�`A���Y&��&�"��w����L5$Ǆph�Rc��UN��ho�G}�4M���!x����!D��z�#t�x�z�� 9��>&#�
�n�n̎Kj�	,e �~��9�+���,��9�9Ŋ�ǧS>gSޟmx���0hWK˫�<"�Z��¾Ny ��ѳ���7ۛ����o~�[��>|��O~��~�q�P�`�1�SQ���	a^_�����_�?�s�՗�H�ss>��Oỗߨ����J?r�0� s��7��yۚs�Ju us{O«��bk �6������@M��ʬ i������Ndr�v���~��|��>b��Y���y��c;n7D�̩@��������߆7y;Pa�~�*|��w�1�%��o�9ú
��d)���J���_�O>��D��Wo8���xǚx�����[����H=�r{w^~�R�T\'*)T��j
^H�o4�+��[Cq- �U	��`��3>Ut��%ia�-ɘ�J���>@f�9���>�Kd}�����5�����O���U:�65c���+��-ֳ<�ޝE����������3Æ�|�*<��Z�9ǰi�
�6��"����^� e5��p�)���T�!#�VN���^�MVXPY�FU���z�2B
�e��N�EM�
?��w�ߪ�7���?0�=k�ifFؚ1s�r�</��FՖ`n^���:���sV���QD	VC*Ԋ�*d%Z�!��N��Qc>�~E!���֋�Ya�f��5ϯgTD�N߹�<ܾ�y��J�"�1בwABa�gX� �(���Q�YM]U��尶�~������M��@�]&]\�o�kN�
��P��<�~�MI*a� �b��[��k�F�c�b�5���a����֧�4����M�K~km���{-�ٔ��R�'~/*�W�]���M�&m൵�R-�W�O/�RQfPu��G"K�z��O���L̠�d�Mm=L%�Ec�[�"�2���/��`����/����++A1r��m����,ۍݠ
�ˁ.ŵ�v�Pn��[�p�u`2B���^��7L�z��emk[�����h+����mmk��5T�M#�B�M�j����Ѳ*��T(�EO!.�ҟ���, �� �@�H��D$L�퀲$*B�3 һ�;~��w����vKh���YY��`�f�_kv���D� �H�M��thp�m���r#���G�g��28���i$�B�l�Gz�ϛ%��ӫ�;ܾ�Y�-�ۛf�,#2����E�����-��q��E�L��$EXY[��#0U��ŴJ����~S_�D
*�+����L�F)_���,u; ��س1ɒ)[�6�^�����Z��>���+x�����-�a�]Llb���~c��fG���!�惾��fOvX��`�JH��Vn����Y��c���AS�q��hT<�JJ�kU�RCE��t��<�> 3�}#�J�([�����"l�&" �< �V��ڄ8aܞ�v�9���۟���J�q#h+$U�$��`X0�Ƣ*=��J������������?�0��y	���]��ϟ�/���� K|pSm`���!�Med���L�	��3��Բp���/�2���������܇����?�؁b��˗����<_���8_|�%A�7��R���pk@g��S�5\םl�	 j�Y�$Y� �y�;�f��`6do�B�p�Q�@�]Ky�.���ddG��e'6C�c�!�	�V����9�`=�͗��NJ�g�C�� �~��%��ܟ?�4���9���1|�՗�իW,��
��uw�#�5��vn�cT��P�}����S7�Á��@�6�<�s s�sNj�g9�`[��{��V��C_�=�Z Y1��`�DT�� ����)��S:@p�����H��Z'�(�?�(P�`��>������	�w�1�y�}�����x���/�|@�aLّ��p{��������o�������?���px|C�1�;��P�Y.����2p$������薇�Z�M��ʯEZJ��܏��{ʇe=����<@�D{-Y�==��� ��5*���(k�R�JS��k<A6����5�h�87����jS/(���)$���!����ө�:o �e��6��/�ca�@��
6HI�Ԣ���@�[*,'�cQ� X� �!��2�X'��r��%cg��.�W�e�j�SC�`6S�{"�moV^4V�`��kR�KՇ�����-�
������CQ���r"�����J���hʇ`�Wn?5�+w�J%�˿��)��Օ���ǎq&8��]\�G���&R���Θ�$��ו��PO�o?�Ȉ�'Zg��h�ܢ��jX����������"˿�?gJ�7������j���e�R݉�*
��0ß���}�k�����a^�A�]��y* �z�v�A߁�N��m�5�qC�/-US���,�FC�9Yq��������������k[��ֶ��W[	���mmk[�O��.�@`T&����q����j֪n�m�/�t������ �ӹ�2
lzhY�Ȧ�y|b\T�%=H�/����0�_�j�I,�w ���1�5p����߇�� Yb�Le�u�ݞ�U}��� �ra�>��vY�Y�I��+�uw���Q�`��ئZD'��!bh~P����lHD?N}K�nq�0�(>aq&v��*;�Iq�[��]�[��e��F �錼�>�{�x��~��,�C�G0~)@͓�ɬR8@w4���H-��my%Ѷ儆��o�|�倌��hD���f{�ir��1?�o�?r�l.�6л��q��u~�oA�Y���[����	�N�h��B�;��z� :�3ڪq����2�� �$K�TC�t�>	rn'�8N|96# ��u�� +T��ߏ�!���S#?�)oB��n���D>Z�o>��!��:��d��k��
����A�~�}�,�}�蓏�e�HP��c
��&�3��]Na|�9�i�2�$�0���JR� @�:��)�z�.���؃�џ��/>�|� ���oh%�YU�^�t>P�Dp��b?7��_������d�ט���&�mNM�(�}��P�d�E*��$��nt4Tt}�>"W�*F���m�Ӣ����`��=������7����O\ǟ={�?<�5�N�?7�����<v&���3z��*�B�p�(p9&�ԟ"32@΁�~x���y����w�`���/S-���5BAڳ���?X�1/��s�u�fP������O���-�b��D[tՈ؆ȩ��&�=�}ΑjN���#\e��ߝ��8���5)irx|G������>����СT�������7P�<X���/������庴��������X�.oH�i�A���f2aSn�kR�0��
s��d%��' 2�^$�@�S��hvP�U��w��[0�9�T /&��R��JW��3 QC`�}m�
v�
�AK�|�~�Щ��fc�`��1��Īӡ����1�j�}�۸�
Fw%#˳���0W�fK;XQ�����H�3IN�N���"S�z��m����J R"l0kW��>��sȹ�=�mg&i�2tc3�}|�� ���3�~��PMb����>���Vi>5.��Y�!�7�Ϊ�\�ξB�n�U���2ď�ږj4[�ENF�B���}5�.E[��4.�9�dd������k����~�?G�8��X*?k�ɭ��L�ؕL�������-�Y9�Wt�
E��#�ogJݼL��{:ç�~������
���kÿ��?���?����˯i�����w@�����#��"�ٖ��QXk=#/5��S�I�ocb��+<����mm?׶��k[��ֶ��l;�C�G��	��L��o�\����x��s��뗬hf�2�	,��J���u�X�s�4	V�)��ʨR��	f�䟙5��f� k���� n��o*Uι�@$@�zG��޾��T�Z�R�8�T�!�/*�K5cX�ki���ip B�[�G55���A�~�RR(����P���$Pԉ"��{�c�wi�6q��#��{����Y�U�	p�/P�xշ��Wf_�I���nDɛZ�I�J^X]�mC�@So��UT�+���x�U�"?h�c��.��k��j��� U�Ѳ"m�"����q��dXK`@���AF��~�;�����Ju$B�b���dAцգ )�$������Fx5U$y������Dr��D��< �!�.X��y^NCg�!Ϥ��ю�E^���cZfÊ��@!T��˻f����� ����g R$"�1t��ܦ��|�0 ��P3�49���hRx��Y���~>��c�K��7\X���[�FV���ľ"d'�@�D�H(@9 �	(䍼}z޾���|�^����_���������W��7E�әaMS�b��V���	c_�;��g�s����)���1�ĉ��k�,��x�������a{�p��e�r�*�χ��H�� |���5�^~<�����}�]>_��T��8�\߶�)3@4�RJ0�{83������g���3�
��\���
��P&���ͻ�,��+�a���$̉}>O��A�P�?��, �T�}��kc�9��&��5?�z���r�JRX��[ ���� �f�yJC�^J�y���,!�G��j��3� ��m�#YI�֥�}���|�0�޼~��%��H2�#�ʼ����y�H,V���YP��B&�n^?�ea�b_ΝUh'Zq5ۖk��5�)
�F���ʴb�[��p��`7r} ����8���!,LH
Qw��m-���8+h~��r�@z��R�����T�')t�K&�>W����8[Ty��$��,_�d�HXcl� ��eE���`�z�g}^��3�U�FS)���6k���I�w����L1�?y�ܻ���_� A��rAҽD����|�X[.����\)aA@s���?���m,�z��������ӆE^�����n�Z��_��dOZ�@��� �è�8YAˮ�!��.�n�l{�ܔAAԸ��Gݧ��v�D�x~��˾u��$��uF�,�YM��ּ�=�gDQH�q�\�������.1Kqʬ�1b��xc@9B��˳7��o��^������߆o^~Me�_��JH����t䱌�v܇b�?�ވ�彐]�$���,���<Ͳ0`5��\%Q���Қ�۵�?���e��^��ֶ�����J��mmk[��~����1<ᣏz��2,��0��?WX+ �{XV�G�~<�ޑ����3�n��p�����h�E@  ����]�Ɯp[��`�s�U	�)��e.E(��<���g	T�@[-<��Z�3:h!���| P~ p,O���nX@q>X/~�j�����$��h<l�Y8&���ݪr��H�LܷzS�0�A�v��'�<!�T���źx���|'�32_AJ��Tz���Ԗ�]���z���ٔLW����*"�}��o�!`G[��J^ eȕ���'��{���Cv��ΊU��؍��i��  �X��>L��Iâ�x(�ܯ��1&P}-��@�G$�`�+��������n�J�;�?! �0����Q
ȑ~<���vA`��@p)����+���B������7y�oo8H��_�<^/�p��[�Z�� zC���<7 ,�vv�{���0��E����R�q��ʤ'�I��`	�&4��`6�N�1:]��\h���˟űSm������9t�3Ua�֊��W�> �sM����>������o��?}�y8�o��ڴS'P�܆Wq`�G=6��ϖS�B��:O}x��ǀs�.o����sd���:����	)Z��7px�,�7\Fl���{pr��>j�&n&�H�/��@�d��)�$U�(?��.uS%��n2�H 1��? q���X@��|�Վ*wf_0��H�Ѻ�9���(_N��aHx��2�m��h=��&��6Rʨ$ Q
������Ǖ��#J����@y���
����D���-�$~ gA8�t	/�{C��>����믿	�|�}x:ilam)2+��SN֧�~�k׫&�j`T�u���ʲ)��r���a9�tV�:�p�MõjH�O�Z�ek�r�<PI��h�ZaM������<�MRm�۪D�N�*,Sg�������ޏ;*Y���u�u��)�D�)#�<��
�9��,�du9�9h�.6S��떪�Y���-|�.�Po����� ��s�6e��~�5��x�m\	`����8�g����9��h
�`�Q�8��S���,��(ֽ�֟
~� x�/��_K"��QE���J6VŷT�$�[f�T����QcY>)��t�Prʒ����?#�wo�e��z��H%��c���FͶ���<i��C�1Ҕ�2|?����^a�li)2�|8Q��u�®�6����ߍ�*���՝�`9�a����a�gb�I�e�ԳB�DI��a��i��i��/2 ��0N��-�K
�q��^`�����Ij���̂,zl��'R�s>�(����	@+�V�"�O�O�O|�;���ρE�[����fF7I��>;���ݓ����?�ӿ���uD;����S8Φ������l(�1��a�VY��V���/�2��Q�v�u&)�Hj�|�{�ɝ�)��-���~۬�k[����3o+����mmk�I�3��� � ��`����!�( �Q��<\C�RK艉����Ve��eDlU�ʊK�i&X[n3�y��4�:��P��@��Ǚ�UES�2,���F�1Xe�f`�?;�ګ�o@t��*qE�0�� Q 0	`?�z���y�������)V ؆BMk>8;���c<�nH�8uɏĹ?��n�n7���ޜI�#H������{(�]���[ly-����	4��Jܨ��U+D�i3Hd���ի�VR��ja.S�sU)ٚCQ�����X;�'W�� �b�媑T�S1�x~�|��_?��Fe����������R� 4��׌���}  ���Ⱦ��.��I�5U�,���8����5O��)c� ��AY`� @�*�ۘ�LeĒ� ���� ��k #�UNJ��Q/��,�DI9�W^��C�m�`SoH*�� BZm�	z�8cb��*�ZCq��|�:t����c��/��������>��UW_�5-��6#A�ȵad<����6MɈ���'dM���rO��]�yD��"��Q�̩���B'�ٙd�Dۭ~"h<�^�������J~�)��Zzή���y,L����o��Y�[��$E� ��䎓�R�Jw����<�Ε�)\�^�}�����,�7�[w%�'HB��77�� ��{�k@�Y��`YV���엶���X�q쯏��7����V��C�:�H�ڸ�����5`j�ڲ`s���$;�e#���%@[yW�c��d��&�B���bI��I?<��[Fр�=i	Fv��m����$����E�A�9���}u�h��sm|�bP�*�>΅�ϻ+�P��V�"{E�4�=��q\KQ�=�U��'9�L0��1��M�W�|],< 7b儛��I��p�d�%�?�i+g�W�0�c�b��n9�nUiVm�m�3�H�`]lu��1�O��U@�Fc�A��s�l�`�o�[��H�7M�쟕��QfR��D���^����P�(~� ��*Ѯ�~_�k�u��"�d,����r��M��v�>�<r��T��W�(㭩�ŵ7ٸs%�|�1�	�x'Bj�}W�߳|r�����֡��Rm��i?��[c����6m
O�[�{�:���6�dwH��Ff�۔���Ǜ��eF�{���n+;:(ں|���:x��]Yp3c�<�/_MEB%�v�;�o�v��NʺɎ��l��#I�s��ƀ�>o"�(��w8��H�I; ����T�%��o�^��b���ݯ���RJޕY��ֶ��m[	���mmk[�O�!|�@��}�W�!� 2����>�r�����ë��J�*��ɬ�@nL��oa'$��BT>>�~��T�`ܖ�+��9D=x{��`�����q����C�����
U{0&��D���J������#	�cm���|�%؀*�`��x��5�x�sߧk�*oR�DJ�@�٤����/^؋Gt'= nxp'���ٖd��L^T�h�ÍU
8��e 9@刓UFT`+���^��M��+O��y����9x,,W�>����Q��b��-�V�ץ�y�j��}7f�f���W6���/6dp��Qe�h؞��go
����J�a(6]���
Q(2��L��<�����lB�%�EZ�1̽����>s�����,0�]%��VeW���.��E���ڪ�V��@\ f��]���g�!*��	�(����s
���T0<�<|���fw6y�}��g��!���{ �@%T] !A:BU�n��6<=�x<���~���	8�f�̞���ɔ,�y��r�f#Xzm���������Aw�[6l�����ʂ��=؇4���c4���W}_*u=ӂg�>W�mPe����)�l	���� �yQ�� �����N�ʛ�]N������B����Ӊ 3cp��l��A�S喂)�?��\�	�'H�������� y��5��H�*��_M��W�Jp�&��s���]����+?c�H2g#���Y��m-���=�c��' �7s�6�3wb�ڌRT��@ޡ� p¢��F��@U�T*��C+���P�$#�bQ�a� N�qbKQ����zz�V�P���b�!k8/^(N���۴�o�>�����T�ٴ�
N�@���_�="?�p���ƮF�W��O���q�y5;6$׺�6���� #'�v�s6��~b��@K�:�Te�q��G6R`��\���Va�V ��wQ9T�B����ŧB���qo��5K��>�Kc1�'����@�BQ�sy�H-V5T�E��V*��ԺQ`7�|�{��A���դ��?&�)�H�Ⱊs.�IJ�M�t/�G���k���yJf����}��3��<o�>�L-�`����1+����T#�ξoA�,�9ܪ��%&��!����.�7�
�)�r����n��A�,�N�6e��$1���c�=�l)�X�ι�6��j���$?��ȹ��ݰO��tyM;ȷ9���4� ��1�FQ��[Y�I�%*s����o���Ň��cؙrdmk[�����k+����mmk�I�g�?�C�V ,��xvw��ޅ��;V8���7O��p��K��?���<�Wp��M�*)o����z%(�۔��)��-�óg��}8��1���R�-G����W�s���nP8��M���bQ�U�8���N��8x�.*��~C�����(�X�t8��(;��`x,r?F����� ��ܜ����Y%t�d�o,V�u�1.����,��Y*����(h�P*�A���.�ҫQ��9��m	�u���$@(��#o-��Aư�b���ô !�`hy%�k�Ϩ��)��U/I�e�?��9)�͈�<)WT-*Y�ǵ#��o߂qq\�����M���1�[@p��ǲ&\'��@q i>��q�0}�xJ(�U+�B� 1NV%�U�� /�g��q�������+���U�R(�!��}U��mKۺp�} xf6Dw�c�Q6�	VE���l/��^��\�p�o��O>��,��������m�?<�s���c�}ۦ��������9_T}�k�Nx�}FE��r�i�	p��C|M��i����4����A��T�UZQ��C�xN�<߼�#H��yA ��*S���N���!�R�`�V�_a��*����߫䞴&Z5=0�n���`�\eFp> �`����"�g�1�)@b������u�����~��y����5�DR�R΋���3sT�C��q Eח��g���N8W��U�pk�a?LR8��+�C���R!�D�G;N�H&�^~�|a֊��'��:�`�0M3�\o�&���g ����~O$<guP\�77wF�ua7f�&+6�%�?��襤�(�2���
�KU�T3��nC5��~K��G"&�r�y���@iY4"Ծjdq�h+8k6Ze�`6Uv?A���֥z���XExթ����l�@��:=�o��@A4�rYG(��c�6�y�����k�������8gh�q���8��Ś	�n�H�T�q�((m�v�xe����i+��mx?��C&��eui�"[�8���ԩ�T���1��1��aL�bF�jsv��q1Ms���=]n�JV�Z8Y�Ǉ1�,�0{�ҭ������WU!e�ä��K�B^�k'<6u�~������p�^��2DD\�d���N������pl2[),l�f�+SuSu�+Rd�P	ĉ�)���=�B�'��o�<����ikH0�k#H�-%	ݨ�OR}�	,=R:��?�ǻ�6|��C)� �N���x]��ֶ���<�J��mmk[��~R-��d���An�����t����Z���H �e8m���i�.��!�l��i	�@$m��S>k�R�,#l�����|��� ���h�SO���09�!<�=�d;U�^�A�h�*n��M��JLK6->Ld ?{T�R�N�o!��İ\�"��T�x憁7+��b���p�	"Fb!E�����Wc����T�k(����vK���"��5� H�/	&�����lʺ�s6��%��Yk$SU�+���M��� ��%�BH����z*������	�� 9�+ ��m�K+-��?�d xc�e��C!�U�	j�^�Rs��b00��G�6 �0c�i���{1�p�.&�a�O6;5�!4ϮQ�={=l�8t�D��}Cr��"�*�,Ϧh� l�T�|/�r'xdoT � z�TM���Uy }�> �Ң,�<���K�����q8�9����"���������N�´�<�ޅ��}�����ߟ�����w߆z�xn�[��axΰ�j�x�n�A�TO�T��N����,C���,�PaP��}���
�y�*�n�޾�*ލ�S���/kԩzK^՟l\��ͪ�I(�����f�� G�m�4�Z����l��1(H��8��QX�YOUa���A6'�Y��/\DDب�2E%�����{n�|�p�8h;���X�̋<���77<&d�`�c��Z�r���ǧp��x�� ݁`8�B�>�6��N�Si"B�=k�0_���a��s�J]���H���օK��da��'6TX���nG��I�;�y^+3X �>�rd0���~�l�����t]c�l=�Do
y�5�p���l�nnn�o��'K���릐_�>s����R�)��P�*c� D�ˡ�ρ?uQ����C��e_��T^,��^��^5�T��"}�R���1�o�#ɧh�V�����a�5+�q/C5H�R+eL~?�@`�pn��s��<օ6���o��7�+>��S!FS�В��k=�iey!5�%\[V���''~��*��y��[���*/�1}MAVT}}Q�x�����k�J�s7,�~tVƬ�杙�7��n�qj�����"�:������7E�"ޟ�qQ��(r	u�cWT�:���^x��`�V������|�+��]4��C{�6]�g�\+{��M����5�-��<�3��Ny�V�\p?��U{4�{e/�*��lE�Ľ���7$ ��c��99�A�*h�J�2���
o���>�NǾz���7%y4�ۛ��⃏�^ܓ`ܭmmk[��~�m]�׶���mm?�VW�|X�n
���n{�8x��iT�����}�#0���������B��m��&�*��;���gD�]if{V��S# U��O� ���3|S��&�� ���`����v5�[ �`%�8Z���+��n-��@�Y?UV%�m&@�3*g��
>�:LT�8��(7O��� ��jv�BDF�m!I�a3�����nq����ev��SM@dRd�r
}�C}�u��.'��Zh�ٿݱTut���B������e �yŏ�S��1f����P,j8�@@l���$`�'�w"��3����~HUԮ�H6^��N�� E�'cK��y8��+�9�f�'85N��W�����C�fo���vA�� ��r
�k�݊H2`��~Y��_�� ��c@]� ��Ȯ	�܏�fH�'�PdѲ-�fe�`sT���1Ga�J�@J�U�xSޙ+`v� O���e߾���7!����� �_�կ��p�� �҇f��j��o� i_��u��ߴF�XG5��e���'Uc�B�5��#ρ� &#��b���Z�+���ϊ���X�9�)"<�9r�.́��׿�d�/��z��Fҍ�H]'y'����D\f�O5g-0����p������&���ZI�:�b5�����SO�&�w6�jS���D�c~o*���#ע��������}����߄�w�\�i)W�bs�6p�s���NqPS76�]�R od��KQ6��D4i�`���kZ2�2��F$��V-C#�fsH���u�C���є����PuΧAa�ۭ�Y�ndEߝ�=�}g�4���������\j�O @\A�6�uN�f* 2�2�k�zS�q�&��XBNscZdD������A\�,1I���LJ�d[,�;�����g�*	a4�ۯǘ�nO������ք�q"��ˏ���y�uؼ>PY�� ʃ��U������w��r�і�A4�hx��ݼ_P0�N��������n�i�=����O�e�>S�f}��l�����f�ǌ}�b�[���JSRH�廗gɯ/��a�W5U�/ۄ-��xqC;)-R���W�l���D�
�j;�c���q����
;I���Ɔdlm6���2�R�����}�Dz���E+6Yf��v]��E�bH�f�*۹��	Q`��{	�Z��z��r����Kf����`]`�y�����S	�p{w���^�����P�a}����
v�I�M����\ u��1�g��h�U������ֶ������Vdmk[�����i�;fs���*tT��:q������M=�q�uۖD����?�(���U�7|Hz{xk���Y<I!�<������M��f%V�g��h;�6��vr����g�@&=t��pp|7#*X%l.�*M{R�:a�����Qz@H����i�a��� f���*�da�!�~�&�~��� S�y��'T?�@a��������4q<��]�;Il-C>� �^Ѱ�/2�S�j曭J��٨п�2�������������<%�O#Z��%�
��B�v��a���[��`��8�����1Oz�*(s�K1�}2$�.E'A��e���J~Q1�j,Q0�2j]�0��;�p�=�����p+|�r��1�T��f�1Ж��EZ`>&S�(g#���2*Ux�I9 �{�s@*���|PGOt�K����Wɑ(6Pʯ�����*��������� �|Z�v�Bf�0k��ܩ������V�+� @C������|���nw�_|�<^_�~�{�*���w����ʳ<^��6�-F��=���F"j&;��(y���=t�b��#�i����@�iE��¡d RU� �k��8z�J]�	�5{B����ˮ(P�,*"@���R,�BW/T�=���@O~�aY��MITE1 :�ZH0�hP17����齕��jxW|Ly�c�c�
�cc=�՛7��o���C�{�5�U�� ��f4��$u�2���͜!�� �m���$�`����}���3���6o�Fp/µ�8q1�
)0�j���0�~L���Wܦl�x�8��i��Y"�,�F~����d��X�xP��<���)�
BkG+G˜"���f���R�2c��.��B$��i�nY�����"��h3y�(wd0[/ íg�PJdO��'T�Ʋ��R�=1�������+E""�l����tL�
���!�5�>�"�s����G�8-�D�U�Y���^�\���.q˥���T#B\sZ�-�B��̨PP���mR������d�����+y���n���]�&u�`IAP{�t72��uOH�-Veg��AлY�y?�xk[�����V�0v����ϲ�xM��
Xv�S��R]B� �&�R�$���`F+F�1.�)���'��h�{�ݙd!(q[.�7Z�ug��6ד��È����B�R�`j
䒌�Mf���@�z���߼'zC�����/�7�)�˖��6����!^�!��dA����N�K�㦱g��<\��|]W�5a����mmk���� Y��ֶ�����&ކ!�	Mu+�F7�M`�����Ƿ""N�ۻ����×_~E����0���}~@:wۅ7��qj@dE�<O���aw9�v��4TLR�t�*��>j	�ң{ZXHl�.�:�V���,�C�pzaU�n��,�&Y�-�X`R�^�İDxx���m�w �����09(�>u���:�}c5(���E	�Z������ϟ��U3ƶlW�j���!�,���T~U��Hz�"��VR�$Vf��$��,"		쿎�����+xs�����(^{�a0 hϞ=0�����ʬT�^ZPM��D�c,�"�q� kZyp��j����Z�w���4t?���컯��EE-�����
}4D�YZ1�+�9�/*��h�6�-`�$���TU�J����XM9P��Zu/�����Jyٳ����u��蟦Ao��:�-Af����	�P����t�^��ꢂ<o���6��˭�dI6p>�&�zscMx|:te-��Aa�<N_,�P�8|���/�*��߅��gy�~C��Wo_��T)7�����g�����f;!ز�I��=h�pQ����+���=8g�Áۻ���9x�T�K}�I3�3�^��N��
�y�RU���s�XUl��{�_a�2����o2%��u���Cq\�a�1�1�+�<j4��5��9��5�7�'NRzH;�ak)�X��%���HqoR��.l������pw{�k��w�����A�N%h�V�!�$�O�*T%d�L�b$y�N2�*`�B�+��+`W�6aW��	ߊ$������B�x�N��1͹�gZ,�ev��n=�u6���ӈ�q [���*���W�Ɔgw��a5��]������̊��o1���>?.��V���칖M�U:�����@6ٳ#H�7s�S�����`��VѢQ!崟�~	�l'����>�D\��*��T�n�R�XIQ���GD�>�#P��8c�{�3j4����'4���Ywl�c�#W��P��el��m@���n�YGS8��n+6���~��*�'�8H��ŕ������k5��F�G.�M��R�ڮ̟1X6D��T<&n�l阉aE���D�3����P~7��ps��ސ�&E�Y[�΅杩M��{%�N�]����*�Me�;+�|�h��o�b��|gп�5Sv�ZN�9/��
lp���|��-o����=KŇ��>�~���vZH��~�j�ó��_��{*�V�B�ӸPx�s�?�>1��n���@�16wx�Ѕ��B��9_�o?�k[��ֶ��_[	���mmk[�O��T�m�+U~ }��9�@�����v8\�J�!0��w��R�r˘�Vx`�L�~�z������Ǥ
�qh$�[�`����a��h��C8�O����a�*XA7X�d�,�@`���4�}��	�������aqt<�Ꙗ/77�a��К��t>转`��jNXl�3j槠�uC0�)��+�m�·�X��x�zZm�
�2@� I���@"����@	�.��@Nye?<�^	��nv�;��S����O�7;�}v�xBXqG���& i���7V���`�[G�D��� �퍥j�P@J��Oq��nQB;�i��z������' k��$�Eu�����G��#V�����a�s l�;i8� ����Z� ��IH��[63[��/�����U9 Al�h) R9 v�Jƾ��'�����O � S�1�ſ�X�	�[���}�>O�P,�b�0�<v& ny�
���%��3�d���@(�I�<g���������P�������혷u���tB��}���R��@���fG�ɳ�,�p�N]���F`��@c�X%�'t'�������-I�?"$���Þ��j� �+�$�z�we;L�,�4&�1PHi(�F���[�:����QY��$A����^ ]1o�4r���>j����a�3�ğ*��T�O�fv{dh�j]!�=�+H�����sߓ0&��z+�w�����Ň/�9~F˕�|��;�w�j~���\%R�6b��k��)�8&��Z��Z�Wȋh�R�Lf1�n�����D:v��Ҝ�'��:����#�e�?~H�������;@��z�5��czImJ�b�Ԅb�Ck�i	nV\�)1Q��:2*Fq��������/e���6M�՗-R��� oL`~d_�T��Ÿ��������x=�|�E�-����,4h�q˥�';��l�q�F\+Xd�C[�dև�����Q*:��{؊��0��
fU�U�O\�Z��4�N�"A�p��
/H�TT��$�c �z*�:^���.嘂�jeֵ���P�E�s���}��R6WT�8ᰰF�9`��Ac��-l��ڈ+˔|��$��}m�h�$�"j�3��*��N�.���#ڹ��U&�C؋����jWrY\�2[�I�CR��U�~�8�,��ƶ�L�80_
��@6%�{0���)�xX�T����a�����Fy^�����֖�]�A:�\A{X:ԅk"syVw\���׶� ��%S>�Z��"]�{�qE�Võ/�C��[)Ǫ;�^ �����~��&_,��8ί?�&��ۢ@�}X��ֶ�����J��mmk[��~2�c�o^%X�S�������={FO��{E�b�u�>���� ��v"�|�+UE�t�9  �by��S�x�,{���/z�/�wb��[N�Ê?y�� t2/ꁕ`������¥�۝� <�oE�k|0�[f0�x��V�����%��U� `��6h�ej��,9�J��z*TjS��a���6�}ۈ�@�������H��՜<^l�}ˣ�1 �l�9s�"v3�U��� ��nqv�V�{������!X@��([\�!P���و�2�N��sTѾȁx?� Bԅ{�f�
s��<~U��AǱ�d�3�Uʞ���=��(�_���r���*TY����,:1�F�������-3^�[{���|; ���_��W#��ɪ�ݮ�K�n�s*�t�
�U�|[�j�������x�9�j�ɳ+柝��^�T�`�j�UhSI��xʨA��Su�昿��+���O~��}��K*Ӑ�m���|u����<H>
4t2����f�4"�m��,�U�fSqs�sU�p����$T �P�!�e�*����1e�9jJ,|�`䁇�o��>l
q��W���:���k��3)��Up�M�R�Ӑ�U��H!�s!�f`�v~���k���h��<�0���-�[h� ����|�A����������,�O��@2�P�Ԙ߮8оX���%y�SE��2�}�ġ��������m_��}��;\�s�k�)c2����e�r��F�9U��$������H<[c���Y9��]X�Զ��ذ�Uf����k)�������^p���u�+�F^WPW�B�Q�B��^�Cr���^�W�?��r�-ǐ�<�B�su��RX�) �`��/�FI�8�b�!�7�� ��8׼�=���3���^����yO E��A_��/yӧtF��XȊ�ŝ
�@����yI��	���!-,BӲk00qa�4y]��b���d������UmbTO�Z }L� X���H�p� &b��kQ��0纈��9B��MAj�'��}�{�i��I�,�ٌ�R\��B�eM:,d���d������ͽ�6�����k��PP̱����n\~Mr�{m�M7[di�}M�I����RE>��5|�r��>�Uv#�:f��|^G�m[2g�f��y-9��5��nֶ���mm?�� k[��ֶ��\i��'"�	_MΪZN�ǉ>�P� �x��� �d�p"���y۴��<�i��_�C&@���T�\���>�U�-��C~�-QY� <{��kQUq�
uV����=����*�4c	��ɼ�U�����#�ujD� ��5M
�@� ��VT�</$E�V>��"�{T�ߢa�Qyː�+~� �XY���J��p.vmUL�V��DI�PU������'V���Dm~�9��S@H AS�#�f�x����HCA��
zl'!��1p��Q �T՝����M�A�}��e��[�Z�?��d
�h;��B������XO���17����83ŉ��}�:A���S�U�7e[��9]Wj_�����a��M��&ۘɀ͉��6�5���1�����?^dG��z35���GU�$�@xT�®}�i�����R�v"�:ھ�x�q�����'����{#��'�G��[Ta�����Z���:�gZ��7�c�2�MZ�E� �S�H�
��)W�T��R�OQ�8x��f���� P����+غ���B��	P�l����٘�9ڶ�}ے�m�^�E�)� Z&�	&'��� j�U��WM*��jb����
�`�5��؟y̰Q�P���3��@��
� �h����ga۫�?�O���-��@�b��L���6������j2�~���k9��;R�`R_M".��΄f��Sہ�Hʐ:,�#e��r�����1�������Q�b#K���VH�Rc��n�dD��p�I*��f�h��1��c�Jf��:Z�;\��$Hݖ�װI	~Am��n�1�8w�P̬	�$�<;G����7���P�.癝A�����������޿�P�h��SV���Xl��I�ܲp2KOܩb���R����|��:���Z>��B����#N#��͸�TU�J��K ��e�\Xb�d�ؽQ��2-��T	�h���|A��2�����)��J4�L�i� փ��v~]"1t��@A�:��,��߹8��jSm�P
yA�P���d�p,5ʁ���rX�;&^��fk���A5z��{k�IT݄�Nk��I>�����)uj[�]}ļ-�_2b���<��3E���5�P�����W�X�l5��MFf�ufD��*W����w����k�|��۪�s;\�Pnt��h�de��B[��N����k��n�7Z��}��ׯ��ֶ������Vdmk[�����i��;l�+�����S��#�t"�A�遶$_�5��_<'�I�8�$C����~���m���i�7�d�Č�� n�2m�"�B�ח�"k�(+T\o7Rt�J��Q��T #���|`�Ѭ��V|�0�[pXA8餐QTN!�e  �J ȉ*Zd�~t�k�h>�"%PA���P	f!`���6��0W�y~�.��� iA@�B4	:�� � ?��T����l�ǔ&{ �	��=�ě�z MÂd��	�l���m*�@�<����_�b]*T�x�r<N�-�y��$K��<��H�B �쁼���RaXu��S�,+���������2fT����1:Mz���f췇#{H�����Y�x ����#���Q�X"l����㮘��DL(�XY���,߆�_��I�	�$p*Z΃e�~�@W��j-�_a���CO�ߴ�k
h)�]��$`�2��?ȄoĞv(����'8fd�m� A����qE������m؀��T�>�g��<"���U0+�a�l�0C�U��A�6-l} <�P�6��ws�/��@m��+�5>D�(;�*�	�Y�Em�I��V^̚�bk��:�Ti~���B]��T���>Z�}!��N��W�4����km�ߑ�w$uCo���@���T��N�W �P`�������t������v���C8�x�<��w<.Z�4M�"� �i`�`P�u�!lȾv�����f��L��ٙ������(@>�H*�ײ�y���[e�s�x�j��"�=�Բ0�Z�ڀli��ץ��}߲i����m�ݫL��ۣN�nZ;�Tv�@b}�[�g�q&���O ��rSU��[��=��:�?�^%�1Np�\�}�QE�o�GȏJ�����I��t�%���'IPLQ�`u ���tev� �@&��Ch���Aa�>��������2jdՕ������=5�m�� `��K�w�K�� n�UԤ<�xu�4-�����.B,��
)���KT��lZ`��I�~���g�ܭ�{�g?͊����dT����k���r 6����������4�P
b�Q���
R���%̈��(�j*K3����ꏠsC��(�F!'��a���9�to��e�����:���y?��m1�GVY6��`k�2��^.�`6j��f	w�&�ヨK�lq�Rc��Ҧ-,�#_�-�'���?��4�+*@�!>׶���mm�� Y��ֶ���d��X���H`�������W/_��ǧ� S)8?����0�Ã*�jY�~����50[�����;�B��iC_eJ򭂌���|�M�*�h��/�������$R�<Wb{t1� ���;i�����g<ŝ��!Ѫ� T�ȅ�ӔP��U
��/��3x\�G ^� ��`9�������vR�fL ��u�Vğ�$
��U��U�;���Pۥ��4��� �����R��H�T�Uy�JZ�D�y�y_*`|��z�}�*~f���x
q���*�d�� �E�<��(�����$	��3�e,�b�69�r=|m�I���C����L^�w��aP��!�s ��Gg �'���X] �"DD�Ay���9�j�B������Tn�w�������N�GfnH�@�W�c�;���I7J� �7�hX����@u�T.R�l��{�EF�g���fc����9�9�1�l�<&�Ƿ�a���ŉY<+�$#޼{��8��Z���QMp���h�6`����J�+e��6)4x�D�%YG���@2�d
�<l<WO9��s����� �v:���X�E���a�5��T�+8f��ͧ��$gN��l� �2O7�e^&��"�v�"�D��=;�ch��DS���e��
T��)��D�(d=�C�$��y���݆�ݞ�����p<I��lA�]�=�+|�VX1�Cl�N׵�N�H�6}��\��W�3 ���{i�7��	*�������Ʋ�:��ϣ/t�8�����-��M����u���ܝ˺�k6,�h�e�k$���f�Ĭ�b= ��@�1�2N (C�=�RF����j�3��3� v�:�m +� an?���w	�����������-�����Ѳyk�=$WAT��<C�>�YN,�4��GJmw�����Q�;-3��&'�*�c`�-�,�	럈
m�k��y6�q�	��Hi���t�5he�o�y�,�b��Ep�+?�afA�m*X�F�$��`��t�V�1K�<�ک\#J^ȕ��5yU-F��Tv�-ļ/�bWd�I����@VIAcJ�~b��l�}d����H�a��y)�6������V�b4�ʈ�����,R�gڕ��h�*��
�z��F��n�lM*B}�2.,�m�X�����;��߸5��������䃧��Z�`UL���4�C�'��hi�£���zҵ!�hI9d�'EV��ֶ������Vdmk[�����j]:0�psۆ�t��[�'P�oc61 ���<���� h-@�A��~y*��ʫ�'>|�c.�<���rp��Aœ���jX�6����� �{���:���o�?�~��9�!�wb�U����$�b
3,��8�� ��Q�\ �;-�s8���jJ��,���
a�d�Nm��|��W�GVC��)xl6[ٸ��6-��`TJ� a�s�]�cV�����������#x�؛��� �mls �L�c������H�뜏TCL���l��f�*n�r�}��0���K���g���=K$.�i�I�賍}^vi�;H�����Tt0��,Ú&zU��K}��9���'�cT�o= ������ � J��U�f�`�Q*��H��?s�o�ޅ�D�"R\�w�Xk����&�#��\&Ɏ�AU#���ْ��+���i��ص�q��cTMK Ġ�K�.O'��x��i�<<4?ܟ�۷o��o�=�0�v�E��jx��D�@J�u�<�b4�E�4�)�(�CYfi�*�BF@&c�B:��r9s��<��oV��U�g'��@�L���� ���D�k��/�BՆ��|m��/��V�p��1:Yh~�M�ʣ��6lڍ�'&a�Y"�|�x��[#8�7-�r7���? �1�v�]����� �`��L�q�ס�ܢoG^���T�^	����U}	 �W�R��l� �ym�m���.v.\��\Yj��NxJIc�h�f<� 9"��3����{�C�͕#ii�l��;��z�A���Ȋ�U�OE�&��P����r�|��R!�\��y1�9H%p�q���2�-���+��b�)T|�Z#�{_3�o<�)�+3���o�T�~Uq�.->X��%_$���,�J��|�u�e#�}S!$�9)f�{�XB,��<7���z0�L�-�h�{Q�U֋��&�o�����>b�6�3&f[8��)J�F��֔ʽU���}�<�܎6�%�kQ��b�
�|��SA�J��*�d�"H}oZi&%=��m�|Alr�6�B��F��RDb }M�,�?w/�	�^�_q�\V�\�k�߄H�ldC���������}�e���u_�y�kB*���}>�R*,�{��=�숩5��(p;L���ѽ���=� ��xo�{d)��s��p���͇��x^kikF����*�^���q�D�˸Y��ֶ�����J��mmk[��~2��c � @M��pssǪy����p8������!�x��Kbp�&x�������8 
��*�6I�Z������@{k�@Q̍�a�Eo�������Qi�]՘�&�MD\V��|�m��G=��{��Y�6���=�"��e��~ƃw�����-�=���U
p����Y�"��H�͏�E��nYD��}�y(��b�a�[��<NonoHb�B(�����<���z��7�����"��<bT��C����o���
|���*A�g�^�M�4�������<~X�m�"D�5�f,E)�N"���]�XV�JgCI��U��p�"�^�7���8�R�>�N-�^������T"���\��^'�,���?�N�C�y�b�����X�3�t��*ͪ������x`�/m����.��D�z k:;�̥�C9 �wy�ip0��y�R!>ߜOasx�-C���vgdHNG�)�����Nա�.2L�9�d�����������8�Q��GuYo��ԙ�G2~4��±�T��Y0n�$�t�M����{�&�q�X�xd�f�W��k{��/��{���|E�x��� �����[��h��ʌ	 �~��T:8[�Vk�>��|�+)�H�K��<#���	�E�ZI�����[t�TjT�Ì󨦐�7���!)_����m�&���O`��j�%P�A�;�B�Rkۗ$�ݲ�9�ɫ���c

#�������|�Z`�T޿�Ƥr�z�6��v��AR��ξL$%�Ɂ�NN�i�AB]c��i�D���"��i�\���ϱ� $(m�3�s�. ��)a��dk�9n=������\D�5�������

���~�'M2��ш��-����+���R}�����z��|h��{$���I�Y5;,�@�lC-po�g㸪��r�u��}p=g(y1�)Rkʷ,�>X���}M��Χ�r�L�I�,�[���ӕ��&�k��_[}���bmV1�|B��[3)y�_?f���0�Fd����!O�}��r&�-��[��uI�'��mL�Xm���5�	���R��Ws���ھ�A�B�R�Š޷t��n�uu�q2#˾Z�O��-v�נ|]3ߤ������z�/~T��H����e��h+��?�I��{ ����*	��G����dHhy�ַ+��ݗ�y?���И�z�����IEG���'�C������׬��bI���R��M"�GΧ�qN�L��yv8M�ubG;�юv��n� @�v���h?M�_�p�$�e~��B;����%T�o��8[���Og>p����<_������F�:�V)=/�����$`�AɃ�M���iʌ1���9�as@{&�0���\gYK���!���F�%P���u�ʾ�!�?CY1^�
S���Qp�_���_�}� �D<�Iϖ�p����?LS�d;��ǵ|��Ƞ�lU�<�����ҡX�D�0a��|_L���V�k/VY�8�2�Jl���K1{C5�IRh���]����������)����Ka桒 �2�"W�I"p�] lK,�Œm��s�̙��<c���C�����J6��fV� ��mգ?�G�� �gr��K�~'M�+5���/��#+b^U��mZ�%��:[+�5l۳���ԬYy���M�,k�L�������s<�`�cZU�܁u�S#�̋�ۋ��%�ɪ�M~�}����@>n��_������R_h3���}_'�At�:q���J����8�˦(�����=���~_�F����rgX��)�}}�>��~���g�@} R�βy�/���=O�~�����,���l��0�G-h�L,�<k��MYe�g��NV2�{���z=�V���J�R��3y&�愃e��{6��?��Y�K�³#�,�,ق�+�<�V
FꉔD�}�_,��q�s���+�z�y�yn��ú@��1��Ym/����,�|�@�d��܅����e��Bl0r^VXP�Q�g �4G�Kd*�Ԉq�����*�]铍�w�I#�Ev2�ۋ���MF����>��~�����"{�P�^Ui46 d������o�ȵZ����}<_���ÚU�}�m�|�F�Ys�?��[����8c�R��z}u��?����l����B�^���î@!����\yJ�;a,{Fo�\��ftD�f��I�����[�Q�:S�	����T3=8f�P�|��}�)Ë�zW�a�m��P�Zg�d�{ŻQ�r=�~����=��sp]�|�z���Ֆ���
]W���/�e\\�j�<��S��b$��i
��![�b��\E���֎Ƞj�O�]	^ kHxS��nE5�z�t�ʕa��K��P�P�k�T�U:�(^C��6�ᣴ9�":˫��IR�H	�I{py����a�H��PI���-���n���ɾg����ׯ|`��=�n$�t<��H�r%�Y�g�_�"<T;�;���q�p�Y�E%�	۹�]�9v����H�x�6�a�%��UAG;�юv�?G;���hG;�O�n����/��//����'�x�z���?��?�I�����À��;,Z>�`�C��m�{��-�F����]>�,3b��?H���lV��o*�;Eyk�֐��i�os�=��p��8Z(��2?�^/S\Y�6�����ɀ�7�o�� �iXȘ��I��<>�e��_���������H�����������JA�=��@����Um`P����xV������l�bۋhZn��=x@)-Ē���@�������۷����q H��n��� �`���/�p�>���a'�g�S��{�q��c��"k'�R��æ P��S@P=�����w�$B_�,p�URl Г��l��ZM���tp��=Y��ZN*pt����!l�/ɐ!�*i�����դhɔ5�M)D��e���
̉�M�А�G �Vt� �eiU�-{�1�oK^#��sN�T����m�e��U@첉��[K�โ��5H�� ��}a�v�lS�l"�@�px�;���"o[�}�)���X� �0	<	7�y�O��6�h��s�g��;W���9�p"�����;�ʼa<�ۿ�V�B����6.��/@ЗU��2�bU���������.���$]�e��C���}3Ӟi���$���F�Q@�2Wt�; �i_??}��urFx8�4�6>�p��������j&�s:%*������a�O.�0P�dA41kA���e[G������ ����� �}~�D�}�z��c�����s�~����>N_ߘ�R
ꭂh��TK P�5�+K&Q@{F���;א	ʃt�~��w�����.cE
3	�O���	�,�~���D0?�|$i����ir���S��κ�k��kG�W)�do�X��H,#�`���j�������r:�e�fM�nq�kB�s�٨ĺ����@e�ړ-���A*��8W�m����\g̏E�(�g��[�c��W��>�Z�g#D����� �J�>���D�M�U�@e���7ƼT�f3�.�A�'�DE�	�,oTn�i��A�Z�6Cp��*6O�?�b���Z�t�iX�C�-V�"�Xc���;��)M�_�*��A��\�bRH�e�\�'];��(fs�Y!�RԊ���Ԭ���%��/0��d�"Uy��z*��L��q�v��Ë���ۉ�Æ��������ysXo�5.X�F��d$�nT�d��4��%�oH������HXc��e_����j�u��儏Y���/
�=o�C/�pW��-�D3�o;Jǽ���>H�#;X��1+�U����F������� �����x��u�9\�����`=�:���j����oK����|y��;�uߴ_�3�m��gS�⚁>�
�o���U�7,`�<(�0��M�G;�юv�?i;���hG;�OՖ�K��>}z���Q9z����,��Q�|����ӝ����`��@�aY�U�J!0ҎD�|�A�]��	��U�: A�c >�i6��@�쑶�$��4+�g�� K�� ���JՈ,����@��.wSH"b	���"��7��I�#%��G����~�}�=Խ�!��#��\T՝��B�jkc_VH��0��;H(W�Ld����Z��}��1+�B��[ ,π�Y�yp���i~�RA��n3����j��Ui�
�fa1��Y�������
��q2�P�����_���u�u�A���W�3��VO�le�����=<>�:����{H��*[�N��8��L;�5�9��	�k<� i-B��� ��s�"����fM��m�U�z��������-�e
�B�iC�	��AC�u&�~pۣ��+�V� H��&Є� �lV)r x ���e!𛧅`��c �Y*sj�A�� ���>$6P
��h�B1�U�OE �;c�Έ���vh2%ן����;6�
���.�·Y��U� ����bs�~��������?��mul��@b��^ˌ'�,��ۣ��.�ǃUL�4H�nN4��/T��י��'�;�����^��4�-c*�R�E�:b�1i`���c`�������sH��:`��Ϯ5˼l�����ޑ+�y�յ�m˨�>w���T<����-�р���P�w��g�vhFt08�R�^�`ln���3�f��1�ȺIVO#U�-j؇�� R�󜄁��R��. 3Y���M�e{��m-Q�S�.r��P@Dڌ�U3X(�e�#j�4�/��ӯ���wq>|��Xd�4�O}���zєm�}�K�4�Wa
�����qޯ��ό�!��cERBt*�U�h��o
f�E뿒+����:�L�
�$e��":Au�����#��3���S��So��C�����$��H����.H���S��j�fyZ�Z[��U����7F����*�=|h�m3Y�"��x&��J�N���J\O������ǖNm��L�Yf����qb�W��gW|�Kѭ`�1��^Iv�^��F�C*E�>���I���U%�#)�`����쟤��d�a���3A�"����3�J�v���h�v G;�юv���}��^���������z<�u!0	X�B%����_h%���kx}�K1��OTUg�g��#�+_�'p"|$@N���E	�*��Cd�\h%�� �O*�H!��e/�������W�&��������oQ�_N�����z���ܴ����*�a��h�1�,���4O$ h�Rd�f7hv�F�+�ȴ�rV�8� ���R���Q��$A*�mx+����@�h
 5ߟ_+��	w+E�_3;VFF)Y�S�����:�׽���b������F\�,�Q�w2���+��@��~�Dv��}��������ag,��˾��� d���Iq��dF��\�}{}�x8�B��1���}6���c���;n����<X�����lZ"=� �X�n�S?n�U�[�x����G�~�c�H�x0�W�*��{�m�Z���	 L�j'1�\�8��ϲ�zp�@N���.�k�� ����� �`/����H ����I�m4�G�,k����Ĥ�´a�%�ο�;Z�؇œ�#�O$軙��{�FS*��2	�����(��׷�~�3�c��#�
'8**���M@�݁�ܔMNtyöj�Mj����b�Q���B�A�"k����F��p����>����gSNm�eI�����m�d�ꩌX���5"��N��o�X%Qej��9W�r��z0z���X��GL !
�D�jjG�޹M����gLT�Gs�	�~޻�+q-��g�G���ܮ�ף��uA�F%|V�=�%�1��$U�����>��,�pܩ�,
P��;�Tި�"���x�@�j�GFP�'�3��@W���X'�N���=��,�24��fVO��ݖE����!��`�cjHq��R��h�Fm��b'��>��Q��휸&�MeĨ�d��K�u������}�g�0x)�}
�d����:����n�X���P���_�sQD(��-w�����H*�b����ۭTU)8��*E�
������}�;��j����n�hC�O�r�������v�S�u)E1����p]��)n{e���[���Y�\R?���zPz�?�wwG�}��d�TX�<s�,�_�ؗ�g�:�Q��-u�.�ߐ*u�E+3����d�V�ǺB	\�x�MѲm�p��!scV#r�]�v���h�v G;�юv����Nx��ԟ�|�TN�i�{\�I�jt ����z~�����|oo/��~�~�#m��U�3� !��+���"*�����i �ۮP���L�d�����%�;:��[��F�c����n@I�]ML+��eu�=�4�Lg�z5y�W�Vy>X��H�Y�X�h_C���@uyF� q?r����e�=�=�50A��6���!�%�xlb�����S���9X�w��H��F���H5B@��G#����BGվ�8��}�c=r0WԀ����SڋX���n�*�,�ª�>VOw�ԛW�!��~m�37��:��j��0�M��sx%6���1��:�b�c��˽�[��<��d���(=Mni%�}0v���G���qBKD���2�r����*����M؛ِ=ny���=訐�BK+����}��OV�R5e�T ���^�#����"��j���}��U~O	��Y�(+���7)��@�R4/E�H�X�U���<�׷w���;������q�G�G�\�_��A���Y9D omݢO�����5]R���>��y�\��4�T	�Z�O8~Z�,�,PU�@�@������j����	>WI9�7�Y��l���#�(�"04��.����/<��Q�9��.�q��#�E�]R�D)0����X^C�^�����R��`D։�yH��
��3	s[�R��m�":Ю���?�H�Jh8��5f�����+����.���?#?n�n�+�|���Ow�ߡ'a�)��O�_HsU�E�7>��5�����1�t2y�xm�/u��qM��>2֥�T'�`f�>  ��IDAT�&�3+����u�)�Ƥq`�:��@B�-�C�6uM���}=!�i\�߽�WYY�HҶ2(��6��~�*N��о֥6*G��L��GN6��짛o��wf��zv�1+"7�� �u�{��Q��G͓�u�����]�zTb���:�9�8;k�S�G��tnG�N���֍��(��<�]�"&��^�;���{��9":�V�"�C�B�>�ﯪ
�?Q��L'�	=������u�I���J2�G%?����=Td!����&˵�5���$��X��Z@����,�H����������jr�:5��H�f�J�ֲQǑ
1�=>XG;�ю�glr���hG��Z��:�����0̥�§�ӧ+�a�ӈ����������m��;���Ф�h��� �-x$gܼ�l5�ǉdǲDzݸ���s��d��$�?�~�E��� �`i��������
R��� ϰ�T�)4�������q���Y� l(JYCgՐ��Cʩ��;���P�#H ZV��G�� �L��`}BOrx�,�m��k�{0@�`E��}"Bf:]�'��y�g=<4����<�B�b��_�?��o%�O�/f��n�<��U�%�L��[�Uc������k�J�8�,��n���/��+�U94Ya���7�G�gl4 C��hU�����RG��j�濄�O��6."��e1��o���x/"	w$L9�:g���懲w�������p>�4�#�㻂�A}�j�b��U��ܘ��qa�]y5��j���L�ݮʻ��>v��~��1�1C#W � K��H��0�=ק�\;P�.p��+��ؔ烌S����qES42o� )B��}~��=VP���ʣz�������rՑ��ٲlF#���������y�Bh95k]ǰ-;��Y�o3X�/TPa��������V?���b�	�[�������+�2l�h�fy->ܰ�m����*�ׂ`��i���3$���9�Y���Փo��C6r�Y��~�������[�jre��M!��G�8�0���\�ܠ�%�`-��>��5��v@���(筞K��Td��d��"�-�Zm�|\؇�6�̨-7�
�R�zs��וt���0�)�b%?S\��Ifw��'�1�Z|��d�O\�2���!Ū��r��;8%#Lx��>_�aȉ�� �Y�`�8�An�8w 4l*4�gw �]d���w�ח�J>u`vέ�s�?�U��9�8��A���E�<��mш
oP�xqć�zB���~�>��C�O�*j��OMᰯn�/�e�8z�G~ا����Ǻ�F���C=���a��0��79��AyC��n�u@}��ԓ v���Ϯ"���}ܧT���3��ӵ�H�Q�s|C��HC��H	�[���.���\���7^��V��x�{D��D뼉�-��~O�y���l�0W�~ڽ�����ׯS8�юv���	�A��hG;��~ʶl������8rקK}�A6�S
�>��������������Z�^m h�рh<\9׃(nu�դ��b�	W��E�%��±����P鑟_�"���z�qU� �mw�8��
�D���FK����2�r�� ���V4����X��$|)uʐ������pl
XY�� �&�uE�w`�9!�|�Ȉ���5�����2�e�ꕮ�Y(�ʝ�|)��B���@䃀�V��Gۗ�U�
��Jll[�l���2�1����K�h�~f1�ҩ��<#^�X��m��G�c�@ta��/��L�m@�b�h9�*��@H.(���?�|��:�y�*�݂ˏ=��`�۬��R[�R ��C�)�@���R��v�,� �*1�s8�e�d�v���m��|��1	�w�f�O��n�U}4� �f��4on����FMۮ�-�	n�̸��}3�[��[ݻ%�A1���C:,/y����f�@��h̠�I�I��q2M�-XM�}����9I�,���z�soIE���PH�@40^�ۃ��C%K�cd]���f�&[:�}�*�GA�}>�����@�����4����~�+6��o�A8��;)���;�Eϥ�2��ꜜ��#�[K���B���gWS.��u��V�/�P	ٗTx�D�T.m��r�C�}�k	 VUoR�h�~�6p�8"���:>�ߊu�S�xo�d�a�3[���܏9L��n��^��Iב8��YK����r��؟"�b=�����)7Ej�}�GS:�A�g�*M�kD.��o��jf��<���G����)���KS��z%�kȎ`ET��?�q	И�c��e2`msue��׼n��iwR���&+� ��G�.u y#n�d��}FGd��EV���d�"�>7 ��1�W,��;	�c4F�$�[4AEWV)g�JIM�}��Σ�&���dI����Q�JI�'��V�V��gkF0��;�j���˾�ۏE )�Ǿ��La"��q%S�\�{$\i�j����}��W�;���l-)�5�ݥ�oy"F�	d�*=L����f_-�-6&�jOfP��V��$o����v���h�]�A��hG;��~�v��x�Ƴ��:1�@�Eferrx:_��]�<�De@<xɌN� ��i���vΫW��*�#�k�3_7?v= ��Ƃ�,� ֪�HV�M���>�Mn#�s�F��`{wV�H{*�C��!���=�Ӊ�>���R��	�wWy�k���;WX��r=lJb�� ���Ŷ��Z���<xh�bʍ�=�
�3/�U �h���+�:
�4@R ��*X�l[����>����,ZX�<� [`���,�H1���ookW��lh����^:A&��m{���$��QR ��<�!t����b�AaUO{�8C�K��"<m|��T3k%,@F�P�P�6�q���>T�?�
50��NJ��5k)?��Z.H!�9E؆�nC�H��3���[_�=�����W0H�'7�u�[W%*��|�q�Z�}T�͖���� 7�3���&0'�|����9-E�*����
�&��kGS9y �.��^�>є`E�$�6حU���½m��
y0�tn���~��^J��@x�d������j�O$kK#�1�E�RT��v.�S<�'֐z�D�X ����
1gFJ���l���
�ݿg��A������;����AV�i
u.iM�7ۇ�okM��c}��oߏ�Z�U��<(Q����V���u�ֿ�̟�U�l�&1�L��Ɛ�_Y.�ؚL���֮�,��E����L�����7l�BS~�xl.iK�G�jcU���uMi7<(�z��h}�d���p^����On#�Ȏ4�5k�o�9B���I%ᰏ��n�7��?"�U8h�m$���,�P�v����ς4�ɳ�-e��>JV���G�3T+�\�!q+�y��f�-��]Yf'#��=�y}�|����S�{�����?��ǲ-��jHu��H�������؟i};,dw8����%�QϗYM�G���S�}V#Zz� u\���cP{}�G"!�K����! ��/��$S]����)�-q�*W�|d����?�|���ʔ��uu_#G�T�ݫa�O��oT�u�l�����lqoׯT �b�,e��Kw��<1[[�����r���/ʴ�*��G;�юv�?W;���hG;�O��P
vWT�`��]��e�X���/�G��[�����4
C�G?|�?�����*��s��%��J��Cp>'?�N����W>�$�V$��l�+�� % o _{�'zm'��` ��jW�}ջ r�2�`3uG�=,tdE�XI���?��F�es ��EDFz�Ҡ�xQoݦe�hs=��T$����Q�<$�:/�-�� ��>�'�T���B `�Pڑ@�;*��m�Ο���������U��L$� 0*�����t!��6��ѱ�sPq�W��8Rq��ޛz.E̙�oO�<�!���KO���R�' �Pu�X�plA� ���\�ڂ�16��?i���lv�گ� ����4�}P:U��a0Ri} v�|���<��ۘv����$|V�I�EO~���Y©By4ňW����-�l?J�A�}�|7>��ל���;�o�U��E|:�sD�#�cю�X��_	@����-�M�@w[)_��Q���S�c�ZU\��k�5��K�~jl7;/4���4�������Y�V0����OX/��f���d��*�k�Oh|�A��2�K��=��}�];N��R���l����Ri�&�}*�G�dR�6���H)hVpe�Ğ�e�R)w�Pdv�u������c��|��y�+D
�f�$�
�%V;�m>��Z��U'�^�Y%?bRn�8fS�����z�����R#u�)vV������9�$�#c�Z0X_�:�6e�;��>|��Ձ���x)�p�:�SFy�4��H��*�]�R�b��\7�����-�y%~��Xաx��}�Z�u�!d}�۸�W��ڮ2M 2��cۮ�XC`T5�����i�	K8��l5��r��m��:�]����r
2���)��J�N%�y\����Tɷ>���흢��.~ ��(�*����v1L�k�	�}�6�C�P�}����b�એG�G�@z��$)��Qf�鯳W=�?�俬v]�$
>�Z(:��j�߽��Sγ+hr;�ꎏ�9���ҜE�A�Q�CZ3cWHDb��EI F#�}�*�#rw��`��u�C�,��R��B�H՞�H�5�?1��TOF�0ˆ��,��|�hG;ڟ��юv���n�w�>=� ���,�~����{8������r%���K�����%�c����f%�T�Xe�Ӿ����Xy����@�id�w�d[���
v��aa1��j��`]T=���-��>�gyw�5L�,I���%��@n���F���$@��"�A9���P+��� #V=��N�@
O�V�H��� ��*� P����ՠJ�BPGU����~ U��`�$:h]Љm�gY� ��v����B��v�	L�k&���e����^�>V���2~�(;��o�_�g��c��w���""��
`����4����V�?����@�n�V��;��I���ɋƀ���R�&,w��U�i"pEB�Y'ԯ �dE�zK����nKs�tVC"]�ݓ�#e�xX�H�!�#Hj�K2+��)U��	}<qTC�I�4Ŋ+\��a��ϲ	���n�����m����n�#�O�y�X~�י� 	�E���c�j0����y9���,�8_.T> ��d�*����4	�5TYO�(����@�@����s�������U�,�`�퉀�$��O�!$�xf?����@1��$ڋH�%���	�[�BCC����H1�o��sl�A�/l��%� �?�_����Y�C�xÿa۷ ����$�_��5k]��f�| ��s����22��F�u�d��۫'7+�W־�X"�R�i�ii�%��@�����ߜ�c�n��1���p�b�VHXc��8Hy ϲ���4*���>�BM��X�͝����cU`_�*nPp��D"[�MΉ`�aGP�:�ĉY�M~����f��ʅ�V�}9&#�g@��\�V�7�U�\{$w}}��)��6�ܲ����s\9T��fŶ!��B��mx�enξ�8/����NFn�p���j��f
	]�����=��}�|�%�t�Z��#�2��0��;߯�{?J�6�O�u亃�<�c�,9������y���něX�p�=�~�q߯M//7�������_���Q��������WΣ'���j�l$�e;t{��ۺ(Wh�u �u��ϟRc����ڲ������症��5$�hc�+�oĮ�Q��V$>���d��g�xPy�8�xy��L���XП�އ�D�Vy�k���s	��0�<�u%�%�q���1s�����@�	C��#����l��FO�����/�{
?�R|�A�/��W����p���+�fy4��C���a�:I�������r�� �p�|C�Z<H	�B�Rt���̼�}������~!e���9�lf�d�U(Eiw�}w���Z��Le-Kb�q�v���h�v G;�юv�������U�:�ݟ�_��H�$�
�����8�����Nx ǿ������!G�
�}/�p�ݥ�/|��>�
��v������0g�ėKS+���T<��6^+����.�s?�j'!+����� Ekn��s{O)������ !�Q�B�������ٙ#T;�/`F���@)z;�9:�z������s�kD�AX�M����VϾ(���4_�R�.�bF�Ӱ%�p�H���g��bV�@K��7��b� T=�����j����^]\AGk޶٬o��1�l)?VA�6�)a@L�B��8|�CH�*˫�o<�����N�HMc��~L[#>*>z�ŭ� �%;��z-�����ap�.~v�]��l�wd�M*�؂�H�ھ����:��3�:"�m��?��p�k��qչ-�)W�x�-���_Fٿ$/iV].Pn���V|�*L#��0�;H�}@�w��X��֎%�f�9>`���s��墸�s�˘���hĬq���ͧ�D�6uj�S���� �e�#E����He
�dH6ޛݙ�)�dK��d�O$�;��ԩA4�[}��C���K����
��56?�>}fz�`h�E���
���H�J�Vd̈́�l�Z!E�*�fq�8~�����Jf5����=�{�Z����$�1�
��J��m�x
U���	:��UTX3.�����G�g���� ���]Rsh}#�h�H�m�忄�}t����<�R�%�Ҥ�;���GBr�;�F����Fa~�ҭMZ�W��>��B���FS����ۂ-m���u=��s�����72AR�k�0h�����:�B�_�sUg8�B���y����n�g�L'�`��-�}���������-~߾��鲯"���Ui��I��/�gqMu�O���pߥ���m���[��ui�#5x���^�}��۪����K����\U9�bK#��c�"��ך�F��\C�Q�@�C��4����a.AVD����}�1U�Rw%g��_�Z(w�V^]�z�*�V�ٶ��a~��~?t���W����\/4���ss�"�QL����Vj����2ܭ�h�j�K>�e��S0&�_ȥZ������w(��M�'u�[�V�v�m��,��B��85V(����G;�юv�?{;���hG;�O�����y���g�qh <dӣ��7Xxz:]�:MC�������Q���P⻬�X@�Cx���}�c :�����a���u��+����JՂ�
�-` �L��ݙ�˲��=<�eY�{:�O��凔�
�� p�sד���3�>����8OAvnoU����6�v�/���2w9���@��;�����%�=l��z�k��YI�)Fhrt����s�FU�����SǬ�p���`%,jX�Y��r�Zq ض=ш��@F��w{*Y�v#�	�Qn����+;YYe,}���
���}ޜ@aȳYʠ�[�Û5C�UFX��҅@h煭܍� R}n]�U���XGFnu��^�g*4�����c�����X��$utezN���I�e����ܔ�`�D����`��n��B7���mգ ���9���<G� ��q�����Y�8T.�m��u�fk��UFV��=��"����^A��M}��@T]����Pa���r�P!�1��u��ۺ��s���C�	P}8���v�G� ��)^�njߏ���+-�����)��T	(#��?UcL�I��$ؒ��m`����۸c���-�I3�?#�+bb�D[@�)��ͬ�J%P�s�a��o$��q<�o_[Z�P7-^��-P�;֠���}�v��pf^l�4���.t�'P*9��p�{�����z�/�㋲���C��iT�V���W�����-�yA�Ǧq�@�*��{f�H�uq����F�lZ�I�h⻆X3X@~�0�R1���~N���#����* ��-�ל3���т�a�;+$~����GA�kl�@� W�m�H�E���_�8V³�kD�����1bD-���R�j�k�<����yqT�
�h}F�mPqɚ�0���Aޱ{��OɈ�FD�o�oN�x�6���(�R1��Ѯ�~-��Y���7�#���3�DfT��W���CgY�7�H~8�#��TnKZP�`7z�D�]���+��K�:ü�j�5^Ux!ŹZOi�{�Z��0g��V�����#��t9S��]��١*�'���n$�Ne�`}s���̹B2{��5j����0IN����9�s���]�n�"-��>�G;�юv�?W;���hG;�O����PC�`������[xyy5�+�Tu��˗pN��믿���B2�D�3�1���ȮL���j�� �)1�<������n�.��	���Z���|��j��[C�@=}J�jV�δO1���qR媬Y�N�r�V8ʩ�oV�j�CV:l*\��^��v�	@�}	���������]	�ߡ	X+���Pk���"`����׷l�P�u �Ԁ�h����ɀ8>|O�0W�~SX���bd]����Fx�/KX��h����8?Z y���I8���*O������QW��H�5`���5@�TN̍�aZ8��Fī�8��顱�@�F�y�
#�L�:0)UB��c6�VC�}\'˃(�2�
~}�ǈ���כ�
��p�W�MS�؀Yز4���H7S�`�sm��%���m��b�Y���DT_<[E��A�t���"H=���Q
V�n��V:�$@��9�B�;G�ک��Z�/�6��A�>D�c�$�w�˽چA)�vh$'��E�R��H�Z7U�[�W�:g��JF�5�?��m��t�>ܪr�m�\����f������L��CP_�6�1���Y��$q^�@��6/D�v����s��
��ω)��?=`W��e�Y��C��̠��� A�4�^�]sr�s��	F�\�>��ɏf����u�e_�H���W=q�ﻓR��+>�]��R��2����h�������MA����'!8�ð,U�����#���y0w�@ߦ0qr�	�z����q�j�z��s������jW�^(}��bHv}��ڝ�CE�>?'[7Xj��O�(�����~��� K3Y1~���E%�4�o���,���X�� ��l���D�*�̵t�^��D[ｫ`Y����v��K#'�m���7J�  ��cmR���T���r&��Zqц��"@�k��]{�G_I�b�DI�^�BDC"U� ��=�Vh�%�Za5HS����a�Fl׉B�@�:�J���kȺ�od-��I��d�������{4ثa�f�۸Mfx�-VH�3��v�<.l\��y�"�9|��^��k7�t%0Ev�(�m���4H��{����t�ЁE+�ʱ����9�HMW���6E:�6kD�Cr���h�v G;�юv���ݙ��������+AXU�S_?	��O�z�������-��������z���}��T]9D������"֒��'
�o�%����_	h�����V������@�X`��$TiN t3�~�*��%@��v�A��q���d�=�@��Ie��\�3�>�-K6UI���Kȡ�����A��0�����������(݁�Dr2ŕ���C�*؋�(@� 3"T'4 n�L���M�/x7hH�x��V=:���t���,�2�j �?`����Pm�r�;��a�Z���g\���� �G;�U׊ck����e���	��2?�5W� �fj����lK��oSe�[ի�)�h���]U~���l4���=���PI�p|��J�]Ű�a`Ÿ,o�O�5υ02`Z2��æ9����PnV�sz�16�0"7yL����V5���A���D"20V@T.a	��A��H7rMr�f�걑$1r'<2�9s?�M�O���1��ɥ
�!�v/�O�� �v��9({$��df���,��ُ�2��p��)�6�iJ��~?����Ǝ�r�^�P�dS$��>M�6���"�
57Ѷ}���*!�����l��DR1p��/���hdUY�z
�Z�HJl%��e;?P�q�,��d� �q��"�SJ�Z��A6��Q䟎[_Ҕ�����e#�ć7�k'Y�}�/�^�������Յ%��[�)���Y��)�n��(�l%X���	���s��a�u�-�q�6\EM5��/�\����0�Z, 6a#?�Rm��ֿ�E�7S�]�l�|["�Ep�R^�A�@97�+�z������ֵ��_�F����S�FZ�"�Cd{���^�t����K����ZU5�h��м(���X7�L�F��@����ԑ$��۵Jӱ�A@:M���������ؿ�U}�<�Q�_�C���ݯ�R>��M����I�rZG�D�ꈕ���@���m'W0&���:E�(b�9_D����FT�w�d��!u[��k��[�=���Ȭ$�$�V�P�)�L8D���S�U����/����VH���(�[4�ؐD�Î�Ε��^�lޢ�K6cJ�[H骹��0t��OOUu	�c�ge�E'3K]7}$)'I��Wp]�	/5�hG;�ю�gor���hG���L��D`r��^��1<��T}yR,T>�.�{���XO����œ=(���Bb��@mP��Z��_~��U����]M {fNd�2I1�R!қ�>�E��|픚�yk@����44�ڇV^,O�,z�������������&��j�
�X©$��B���b�-��� ���D�ނ�	,w"ߪC�r����oo�
>��4�qMA��@�+����O���`�K���gx�j����+"@��e�ɲfZ,r���TH�h(��G �G�X(�Ε��>>��R����ú���/��c���X��h�����"��D������<�����m�<�Cj%lcl |.����������`�~?z �ǠWmS��v˦S#q0?�#�Fu��x�V�cN�[E��<S{IQ�����vhPu�����6:c��q�H0p[Vi��߻������\��n�M=�Z��R#�ײ��y(��38vW�̫Hz�c�b���G�[x��@4�Oh�A6k wl�}�͹�j��ɨ
�j�T:���H��MI�c�׷~n�l�5׬���T�����".���F�TU/�x|�{3�t6��e<U��� ��b�c���%���na�4v��)��%�XRTS��}����<��j*�)FnU�A��s�uk#%�� ��SO���q�4>T�7���['�,mb��Ѫ�������5���Iu��5�}��hW�����Gb�+�e��uT�yB��_S��|܎�Y���u�=ր>�d$���~��c�:�O���M��q���/TNŏ�*aB=���g6����f2�.WYR������y��B�ԫ$�P�]�D�`�+���t����t�n�
�@�p�*�:�{)���RD��Y�^&t�jcm�����v��sU+�[��zÞkJ���r�>��U�Eb͏��Ĉ̠(�	����?��v��8;�PU�ɬ)�e���9[�IQ�W���<���i��=����<��5�k���7S]�eys=��s�W��븩lBk<ٽ���a{�Kh0�hW��5�D����?�u-�M���V?��'�q�����A��~�U!���r4"+���wBem׬�v]d
I�2��rUG;�юv�?A;���hG;�O�{�X�]���z�|��zBx聯���s���+Ç3И)�ߞ-�`�� �s��{<���������P���@��C���fe���㚷Z�Lb s�|�c{�'h�_��j��H�bĵ>�[������׳��XhX)�b�a�Y��U���2����끵C4�x?޸�����`ھ�}��NY/��b�J�y�ͅ�Z᳓�p�!F�T���z�VI���Z�U���s��Z��}��ʰŪ�Z�O��Ɩ�9����e�^��oh��y� ��<��p˟aX*@���Db�+֕U	Z{�����gF�8)��Z����ш��|��ۭ_PS��T�,a��ϵ���*�>{��F� ��}����U�3��%��4VEN�6���T�g[662'RS�P���b �+� Ӛ@��F �v- Ly`�Tzu�E�X�C��j�kH+ׁa2�r�%�x��n��I��॑q�<\��-�p��նU)Ħ`U��X4?�u�1��� c�U���i0�e�7��* �>���������Ch�5U�+]R���T5Q���{�����v��q�`\)T{�*'��FM�eb�6\��Ӂ�V���I�m�t��g	��c��Vu_�'�y,����2D\������b#VZ�p-s^�ک�w���N1g�^��|�Y�RU��zŇ�3=���wBwI{ >*��x�YR}`D�.0���UI��c�/�_��QY}�2曪J�V�<[��|Y�}�����RJѳ*�Р�$y�����i$bc�}$�[��ͫHM�=H��D�&+����W�9�������	G��~��#�	�(P��'N�EA߹l`��ȶ/�f��o�]'̶��\�k������§�
B~�^�_�o�������N�W؏N��D�;c-`7��tֽ�t�w�ǋ�c �(��4��g�/�I¾6�w�����\��xA�3E
���\e�RI���Fn��H�0{��dUAI��Pu�'�X�D�Iyn�B�����2"�k�����0f����m�:���kT,e=q�!���ɬ#"�x����sԠV1C��[+m��^,�@���l���㛲7|�:���]3��b䓑&��v��Db���{rf����!�^���-�^E�q��w����1��'���{u����ǈ\K%�bU�n�+燋��w��?"��v���h�=�A��hG;��~�Ƈ�P���|��!�����ux�"��_����x/��� s��w@uL����9��C�g3m��XU-e칗Րq����V���?�)zp���C��iDM>V���B�\ܛ�Gt)��:���c}�' m^�VLY����'=DH������5)4���n���~� }�` t���~htز�e���yly�u�H�4���*�,�u ����9\�mĉ�5]A��eE젌��B2��/E!�F�"�B�s�`~����#�m�@�������
a�XE����ޭ�S ������U��;ѷ�67+���m��\�8��B+$�A ��b�͚y�=1&�nnS��p+���1t�Qe��vus�@�/���P�@X��Z8�� ¸����h{;����ܿ-��! �E�aj�^��V�sv�瑌j�L�v+/�S��x\��?Жu�*�е��n�e���T��%���G�<[��J�K��U`�>�1s�7;��2�v2�G�ֺQVXY�]�u��E6]�g�~�~���H��YV�PL	1��@���S�a����f#��b����AE����\?B��ո�/���Hq�]'�п���yY�)��l��N(w�oTB�RpH��+��~9X��8��<�_������)�ݡ�ߨ�qZ��q[%�t<�^{0�¬�D��^ي%�A�Q���R����J�S?鵦���1Ԭ!W�T����߈�}'Ep]��e�q"r�,nl�tR������'�Zj�x�؆:�=�k�>��~.. �J��-ɬ�\=�D�"3����f�3IJ�+�3'?s��m،T�,F ����6���O8Og*;V����L޷CXns%�����Q�S%t�z~��v�{�!c�qbߖ�w�LF@�!XMaL�u%������S���/��k������?��� o��k�>_���-�{#S;i��T\"RqO�	}�{��I�}��xe�E��A�W�U6�TT��nk[VF��^[�W������Ӕa���>k ��̴��I�u�zn)�YET����7ԝ���V(�`��w�
<�ˊ>xJV�~qnsNs1�oTh�.�I&����q���zbp]�u�D�j���D#�U������!����w	s�ϟ�%�Fh�D�������ܗ��
�,�}жe��p�X�C�%!�o�f��n�{�$���+#��]�c�~U�@�`����F�m��hG;���T� @�v���h?u[ �n��P�����Ƈ��}�=����%\?����5����C.���������nK���(,���ć�=�����p�잞� "x}F�[i͔����>]�<����bՀ� ��(��I�bUy��~l�̦�O�� F���5���W������~O�j�P���m_` ����e�?�����.St.���|ʇ
��`E�i��ـe*�d�$�����b%~�%-���}�*�6P�~�oa���f��BNlXAo�'y��,��46 �o�������~��<�B�s���}<��b����`l"3��h�yh�8�}"�-t�-�A��~|��-�/�}�><O��g�:Bf���}l���ׯ��t���z��ۻY�4E��}�3I��ȏl�TN�U��^����UN���c��P��8 a�Q���D$,���@��6l!�oR�E ~�{P�E0��z�zw�u�b�4Jm����;h�p� 4�� b��f!`l
V�Z�g�O�0�P��8Ȳ��25�}�_*	RI�9�@�%X.�kW����X-���B��B�I8�x�-� %4�F��CY�T����h��#+��,��~��oÁ*�ܳڵx�*c���3Upy�������}�M'UI;ɇ1�7���t�����Q���������!�ɬgL�4����N�¾8xo�a���O-�oE�-�*�������9�U	�����q��u�k��� �qжj��:14y�ss{�Y�4����Ü�Ic�䰫{�t�z!		 �>皏�� ��=�.b#�0����_���[X9_�`;�7Z��;8�l�lF4���E����؎�#7�	h�3���c ��t�*�rr�|��kC�3�����N���`65%��@��+�9���D���~������Ƀ����e�ޏ׫����q�c��ɠ}��Y���کV�5�6��u�g���2���)�!��a�q�ހj�}lC���z㚏�����k.&���2w}�����~���?��2�l���ؾNb�-�ZM񃆢�ol��:_�1����׏�p����k���������Ϝ�~}�ud�k�~�p�5a-��׻��"Y}8��?�|��������<IJ)f����^���X�u�L��)F����*���'~o��A2n����u�w��hVW}��>��ɷA���m�pNU����Y�a>І/bމ=O'S����~����&�9�u���O�o�]���,0�}N��YЕވ&:�{f��$yE�F��rq�p��4*��m, ���� �-���6D��k%?�]��f;�lN�{��������>QY3���\��~x�T����T`�u*M\���S	<�kg��u@}��,�8��;`��@��51<�̹���5��d)���@�5t#a����hG;ڟ��юv���k���Te�
��5 �%\���E.������_^h�5��������g ��+�-�е������YQ���ZuZ���*m��6�i!�]vD*��Ϫ���I�r�3A��ʟZ����Ў�ܳȎ��)|���9 �����'��T%��ri�Wn(0��
�y��s:��Dy�g��-<k���%k�e�}&I�
q�7>:�`W��q��Ը�N�d���`���Rs%d�1(��JC�P��7il�~n[:��U:xյJ�b�,6��H��"����o>>�﷫�+S|zo�`��1 qUg��|/��fK����ъ�;��h����H��i8UpN�W�D?�71.�Υ��&�����pa��^���qB>��9k���i;b�+*�I�>SE�f���AU��Z��-GdS���\�;N��V ^G���z͚?�@��ơVຕ�}B� �,�A�j�~�뛭���c�J
~��:�R�9!���O`	����eH�Zi�����B-���Ŗ:^ȷl�ڤ�}[ ��˙�H
N[Ⱥ,�e��l��edA1G�����j齯�r��^��+IJ������쒆��H��ߣ�F���H5D�#q��*yd�:N�~T2�E�H�s�8�TN��Kp���0<h}����g�MP���t5E��J�9�q"i��.$�6����ɭ� �c��l˱��p'��
-K�U~ ���̯/�>FO�T� `��
�ߨ0�un��vNJ��}YoJA��s�)����#ևfaW|>�5ƕ(����6n��y.5�=�g���	����2��t���(�J�%��u���y�� G�7!�%��Yݦ�ԵE��W$P,S�S�\����fd��Xɋ�LN.�k����	㍊�l�22��,M$�\�*@}������������H��Y�<����9�z�voD�",����r�4�}�U�?���-ԓIvS�m�k�9`o�W�'��u��?ٹ^kaB߼��e�� #�Z��PVY�4#�4$W��n[6^6U��N�P������ynm�Ӛ
��z���\\9ٶ��ѭC}�]����RܺTV���j�K�:���`�V{�8��|1�XU���r��_���P.Uҷj��UqJ��%�>�j-EE���O�<�x��M�mk׽m����&y<�Cݖ+˸>�_�w�9��RJ���s�9�w�K�Jt��c#9�^��{pG;�ю��nr���hG�iA�,p%��*A�u��Q�����(��P-��z0�v�<��<�?�V[U7��WU�����F��PwL�d��1UC����b��}��������~o�x$�,Tj��(m�4:C�[V������ �)��ލC���])�M@�֭��=LnV�{w��cB%����^駓�I��`? �I�%ɒU��#՞�<�&��s0�����iߴ�A J�}����T>jۍ�H��5��VUB]@�8<�77���U1�Y^����,�Q̪M-��"�A{��Ph���'����ۨ`�^���K8!O�ɪ��A�!�׀ͮv�n��0_J�c ]����;Y%}T@u4Ň� p��6F�� |�!�)�X�H��YE	�����)Mm7ٰ�dr�: f�t�,��2o�U~���yg76�K����BKl�_I<��1K����W�e����,C��c�q"Qhr�J1>�� iXod����B�Fl�|���q2���Q�SqfdT충0��4ۣ�@�8�u��v,f�"Eȳ1Y� ��mΤ�J�������Z��WV�q��
\'��y����`����A����G�-Z^�7R�Ji���9�����MEB�?�FZ)#x0�ºp������3+�U}N21��dC�LY���\��[���<��7��4��bkd�h,R��>#;�D-�dq��I�F|��.[�l$�¶���ƺ>/˿l����8*��8��8r�c'�InE�??Ҵ�1�4'?|��x���E�^�6o�/�H{9��c;��,9ޗ�~0bt^�
�sAc�@XO�
,Γ*�AR3[ê�OO�>Q�ֈ�Tm��m�O_�hb�GlC���S}���^��C�ͺ��Q9iU*�H����=Pȣ�@q�)\��qM�+�s����0^���K��?~o�o<G �/��-�@��wY�$LA`E�i�gZX��[��#����JZ��d�r ��G������_/!�ٵ�HQ�\5Z�e^�dAXLYT���r4tn�w֏шS_�;b��ŉ��{����d���1Ly��5������?��5�5�:��VǬm�M��XWL��*bW��zE�s��SFX�~楌�sn˥0w[����h�@d_G nKb�Ӫ㻨�X��f��c��7�k��[��(P"��v��E��"~_��5�bE7����!�������hD�̸߄�5Knw�5�a)����hG���� 9�юv���T� �4�RAU����ĪB8�G�Ysa�M��dx��o��>�;l
N������@$@O0�oѕ�怨j{�U�+8=�\hn��}��G>S�a��=�f�.H�z�����@��.��T��d<?���Y��he��\���J����0=L�b�9Һ��z����o)?����yUU�x�}@2x�Y�\ 
�R�[� ^���J�
a�jYj%z�:V`ED	�w��B�N"��-x��t��R�t5Oz�4��<�`�$�N�0��J�:�g�
��2 {�^A�������xe��|�ˆc��' ���S
pl���bxȘ�C̀u<]���S��~�����ZtN왿��m��H �{H�vΌ��X��xˣ���g����X�p�+����5@��
����sY%���`���P���|$���Ji�������S]��*"	�ru�f�Uk6V0&�����.[��w+���o��=������������*��I+O�-�JU���#�XO\��X�"�V!,��
t_�R�;a!�P�WvPm����
Q ��?�ױ������	(�&� ʍ���l��}�����Hxl y�Hd0G���R��9�f*CX�u�a�'�F��8�@�t�Ў� )�C�f}8�)���S��1�Ū�y-s�m�lM��7�}���"5{��ًyPq2��X�jq,�Vp�
ӗ=�C��T3��z���j��YOv�6��{շ�N�$;��)
Dn[�Rr�<���5m3ŗ�aX]�����"2�,��B�AYOR�nf�~Ff�����x�(��r��I;_�x���_�'����,E�&��/�I۶�jЧ�5�k�$df�)�x�L>�k��Χ�'.���u�}�<�_{�����}L]�J+�;fe��(�����:L9P�-�%��n�m�n6{��a��#�x�����������pA��_o�T|�.����d}UOM��s�kO��^0E׺�k����ٔd�j�ٔ&Xpͅ� ��h)��ع[q 	�d�b~�&� ��l�d䫯}�9�bc0�J��3��}���8�G��27���$"�=�\c1�?\˳^9�����2�J�P�[t_����\�V$z�J@�nP�Ώj3�s��WD��Uɶ;ȍ�R�b��f3�_V���$�r���h�v G;�юv����>U?z4������p�7�O����|	ۺ�_��W�\�����?�����������mi��J~�U&�Cy}'AB;�NF��i���A{����.f��ڨ���P�I����T ��*��g�f[��M�u	�SdU���{�o������M��"?{Z[H�����f� �ofXl�}���O��Xy6Ī�����r`��Q�qP�7�IV!|�Ȑh��X~+�⋁]�C���z����8�ƨ�� �(�r&�����q����(��@��~9Vq���5���l��2R24G���K�=I���9�\�����7V&�B<����ҡH��a��WK�A�9j/'T�ǫƂU%{��7f D��g�2CF�|��]d�Q�O��E�渝<`��lU�A7�^��
|OGxx�l�b���,�����h{��$�4`W7�	�:��0�CP��}d�V��M�xҦ�^k8jG|t��Y)���*�(�8�ѭk�*+�րj��> �	�Z%��6���V���B��C�޻�\�� ���ֶ�w{�b��[~�B��O�*h����r��t��8�<�~n��,�V����F�l�
�Jc�qQ��[�h̴�����ř@7Y���7��@S��)Ș*�jwR�F۬R9k�� An�z��#E�H���$c��ln !Ѫ��:Vч�L��ji3��Oғ�B���[c���m��y�5��ea�6Ŕ͐�4nq�_���+0xjJ4'��86!环ݕ,3�әW�8L�Ӯa�'Ehk�9~�T����������,58y�C1�D��D	Fq��k��U'3�� >�l0���ne�ċ	�*LF.�z�n�Jt89�}�l��ĵ���ݞmk��V�#�n�g'����Z�r����=GQ^�y���k���k�o���A*��w��k����:עYT.�>�������kn�r��G�9.
+��(��K��4u�~4'���15%���{ư�zTG�uV��,���^SԵ��.a|7���v'��`S �e6��9yP����|,(��Hd���hM5U���]=È�f�B���f�4܋A�1�U�,[�:�A��!q۾�T҄v�>UcU{���4+�x$��Z��s�o���,2k���T�~���˯��ؐ=�甩�����U�j�F�P��gګ�rU�+}�@��){8IF� ;�юv����or���hG�����"U�23e�n�����K����p�\�o�����W���;�����Pn�ekD��j{��6�����|��pp{�N4GڂI�	
��^B��^E�i}߾Ǜ f(�O���Z�@������zTU��(�w��3*��쟝�X-�z"&��du�6�?�V�翯y!A�W�{`:T8h�Nf�BEĪ�Q�٪�՜@j��ت�QQ��f����'����460,��Ud����`Y��B2�<X�dc� �����b+�{� ��&�*$�}9]*�� !��|`%�*�Dj�.�n������3T"9����zU��#�����X�8�����0k"#�&��f	4U+�*xY���}���K�|̓��%+�^�H�m��X��ե CQA< �D� �_�sJ*�0�G�XX���W�R��c�&�o;Ś!P���֯'FL�]�0��S#� <��@��
�QvQ�����t~25N�S��~��Hp����l��eO�q\��x��
�M�S��eu^r�@ؚ���@��N�W'hph�&�����2\�Z��vL���Y.E��9���Ǌu`++��7{o�$9�%�����Ȭ���Y���M�쎐stOwUe\�ÌP����!�5�k���? ����T5vm�v�Z�d
�h�UÇOm����҂s����2�4\G�nT�/�V�+]P0���J�d@�]��e�ւ�wɲG�=��$�����
]�>�u.�R�V~�۵��p�-�z���a�)36���@����,͊fߟ����5�l���H�%�z�>�=�NR?TUŶ�Ana���w�-4�+�������@����j�=�ل�8�W�����g޶�8Χ�g+vI�w^�!�W��r�����씌�[�9��d*����e>���-򦶹+��^�7�"�|`O�|�l�<���qU =��Y�.�W���w!���-�X�n���X�'�0qE�ؼ7w�u��ӴH}�m�w{�i����ݏ+<'t�T>��DY4=��fZFN*��s�٫��R8��v��f�D���a��&��l
���_��r6b!o���`5"�Ⱦn7�q�����族>3�f a/������65C2[�lVo3�:�^y���U��������ϯm�V���Ŭ�bjk��6��E�y�����{��f��AL��j�23xfW���{[G�Ǻ(E�+"��溷�Yw�紬����Q��F�6�E0���q�o��]L�Ɓ��L։�'�V�T�}?�hG;��~� @�v���h?LC`*�����;k��-@a����F�K�Ɂn����^^�
"O=��o�MU���a]���n����Fi�ܟ�|�?>D� ��7p_,w�X�6�"ZE>}�U�/�f��@����pdt#���ߛ%B<� �{;���	��.% $RW���۝Im�C{-����x�m�y�g��X��p:�g����Cl��,����
 t�[�eם���*��O�:%G�l����uLf� .���K��Y׃�;��m[dcA�TXu(��qN�e�X�HJ}P�̢
� ��U�ճ):��R��l�Ζ!�`��� NB�a��)����n�]×�gV�
8�{�ɪ+�F@ޤ%��T&�O"���@��Ɨ�@"�j`���R��l� ���g�O}�2Ĵ1�����ᙯ�6�uW.h��@6�<�w�]��}|9��t�����Q9-7$����rT��,"� �)>j�|�e�g�UW����jT5��g�Bʎ�n��V��V������Q�+�Q��1�V@��ԩ��F�o}n J~��#�*bKq;*��*
�qP��(���e�t�����+
�)R2����n�E���KT���bvf�8�'�y��L9��`�t�)7��@��C\)��1��M���S�x'�L���m�g����T�1J�#� ԩX�Y��Z��V} ��^	s8W����FV~�C~���-�� �x�X��G�l%��2{6e��I��:t��54˚Vy]�z�F4�����'�m~��Z��X���m|X�١8[��q�t=����5��߻�cW����Y<Y����HxU�8�8q�l}E��~��=��ׯ��X�)u��vҡ�L�����@�>��H�N�OW<�n �n,̠`1JsW��@�9~����y��ߏ<���v������H\<�0���Q�.ԢEycݩ�w��=�[$P�'�n��̕��eX�#C�wf���y��f�u�e��.!�K#@D�4�:Sy]+L�\��<��&՝>�P��OT�o'���]m��7"�D��Dh�Z�7;�β`�v�%q;M��p�6����T �j�ƓP�X����ڈF)�L*���+>V��4��}в��jJ�9�+��.�9/eE���u�������a��������n�_����	9�BYVgn�s�j�n#<i����C�9��l_��߃Л�,E�;�/�ڃ�Ա3׵Ŋ���7|���L��rG;�юv��Q;���hG;�٦u3.�bh� �A�`����U�����sx|����_������)\?FV�yV���=��!<a�?.䉴�����*S��[H���T�Y1)۫h��|����ќ|pB-[��~���!q*���W�)P �@V� ��|�E�,�G ^�������=���'��������*��}�J�)�)XU�̍9�y�� ���LA���S@@$���*�s±׎�P�]�6�6��I+��򀠥�f 5��P̓<gY��~U�X���L�r3X�9���㺙'��][�e���nV�}�- Z���<>so��?�y��|^��-������5�/�{P)�`����U8�B�3���č<��g8N>��۔8U�sk��Y�EU���ٵ�Z��F}��_��̑zʂȃ�� 4���n\Q!@�B�k�:�|��V��98��@, �j�N9,�I��
F(�вo��2B;7�+) uﭏ4�4n�M�z����m��Δa�$&7*��g� �.x݀|�HP�/-��_oW�E}�50.�f�=�������po����ٹ�|:�}�W��{As�C�2��O��:T�o�(>~��]��GV��s�����8$Q�+=�9ެ��?�{6f�m����Jˏ�k�����Z��P��θ7|g��ꊔ5昻�}eeGq=vT�e��  ܲ}�J����m�¥�t�y�:�$0K�3,���kS �h�����SP�Yy��:�����w��"��0���l*�d�-W�8��$r����͸��:�B۔����������*GY��5#&Wtm�<�W�"�bqs_�6C��L�}�8��*eh��H;1�[��y�.�\����yn������ņ�T|a�0��o��3��n�B�{���2`N�s��=������c@9�����?c	<��Ԇ��Hv��kx6%����wr�d�M*L�?����Nu��#H����b]#e�QŒg�K��U���PY\��y���䔍�(��`��g|/�hh#��ٝEpQq)��}X7�I��K��bLJ= ��2��X���Z�r��f���2�O<��8�uS/�-��8O��?��ʑ��`��Os���{��j��ik��]6��3<$�	�t���
4�����ݴl*�e��bqGS�Fk�$Q�w잝Рx�h���[f;<��[���?x+�,�"�@����N��`�Kx���˚~���hG�}�� 9�юv�������Xw_�%g�F���?��?���S����������	����"רhD�#A��|�Y~��ķ@oTہlXV�M?,(`+$�DJ`��ɞ�@��̂	�L�4 m���{,�D��r߬2X�n,���=�$E�_�d [��~��⠍�� �إ�,e��pI��t�����85B�@�t�g�)6���yc
�̷�w��!�} ���������<���p>�?f������U����kν6� C����J�:+;`�����7������0��zH���}���*dM�I ��^ս�@'4���=�o8+�����������E	_�	�nw�k��a?�'���#�6 ���������>>hL3� ��#<�އ�G��p�c�4�ݮa^7�=	�������B�U���M�_qp
���V��~�9��x�O[�uL\_?�ҥk^�c#^X��Α��u;P!o�A�fe�2�=�j���b4���f1���u�%���L�B�	d �c�j��H^�(�mX�^�?����i]+�6��#և�n���ֲ^�Z65
��Ҫy�b���-�,`v��M��e��= A������d=��,�PE�~�����e]�����1?}����o7�\6%�<ڍ@t�i���\���:���fs� q���Ivz 6���0��'1_A���\ ̹at+����g�ļ�j$|4��Ϗ\{������
R\ �'���u�\��p%WP��~����r^&Yۤ�yi��^�����A���N���E$����B�$���
�3��xo(�� р�( rV5�����P���o��� <�#�_fEL#��U�ԽϷ�9N�`m���+���
"� b�#æ���,�ǹ҃��RL}�x���;��)��6G�}(*��iT{�(f#9��̦,p{(����q~�֋����ރ�\l,uF�r�۵q����k�w��iW�^�mX�>�@�-�~V�[��"}��|&Hfy�R���ݲ3�û]���"I:�/��Ù�\������u"���B���P_����Nf5D�}� ��j�Ö+o�~1+7�uֱ�g��FH�<�?=_؏{�i��
k�;,@{�Xo��d��m���n�RXa���u"i���gi�*(T���^Tt�D����Sgd�B���T����\B��vF��%!�r2b��τ�֫�Y��F�{�L1��m[9�w�?MR�<=<7�!�dA��˝�
�E���DJ�YuX�w�&�|6��H8��v�=st�>R/\�b�ˇ��[��X$3�6��hi��P��]<
5]��8w\���ٮw�]��4�y�i�{H�;�d�3��L�3�2�XŔ�q����x�����юv�����A��hG;��~��`T�x�}��BU�������x	���^���_������ny����>P}��$2��F��g���u�w�<�O�X�)�n{Uȱ�7+�3 �Z.�<�� ܺ�[�N~���lI�P����v|U�nC�0�|W��%8G ������	�ܢ���֙`6@�|x R�c�[X ��x�T��&�P�;�c�r��y�f!r>*W���Ԫ�	p�ά���X��U�����|�*� hp�1�n���%�Ǔ�S-PI�@��߭B}���
vnȭB۫R�3$P��,����{�l���QH�X�h�O��T��N`+� �R$��l��iܬ�����tK�Ȱ�m�[�G�C\��O7�b�=D1[���q�-��af6��ؔ7�Bp�%8�����p\������j�ɪ�=��8��� "P[n��	3J,8���yT�oq \�ﻦ:�)5� �)i����= ���
ƪ^[���`�mi�!�Ԁ/z�,�$X��� �]#��q� Rt��LePo�G�c��e�zY��.�$#�Tm��6$�1�4��W͹�w�_���RSp,���~��6��2aO���@r���9���
0�ͥ����I����^O��J�{�mc&�,�b^�ַȶ����;�NT(���+�<C��U4�@qO�j�8g�Gk��T.��EL�������=�����smΩ�C�iG �M���U�����������U���6���[��zCĊ�O,�E6\ш 1;N��+��;ę�3�]V�m�uT<t�@���W�WW"�O��T{q;H���b�����T���MUȹt{#�lj�'Q�hM) ge`��/�h��[�"�	T��z\�X�ҏ�d��%��-�ܮ��+�}�fs')�ٲ�@G��^�H�*ڙ%�s���yhx."����z�YjES3�{��W`���s�g�)#b��R��m���''xn��sN��2�I���k���a�?*NH�o��^Eƹ��80�T٨�1�Χ�9u��x�sӹS����b�y�o���ݩ�0>���ϫ�lsG�0z~��ӳ(��;oF�yK�Pk�+��<-���u���R�1���Gl�B2����0��Iޣ��	�{��h*��ѕ�X��R�F�oܯ0&E�����α�� �k�D2��S�#Z�JSvx��^}�d|�˛]3���p�����hG���� 9�юv�������kjC��ۆ���Sx����sx������#�˿�_���
��� E�\�\N��(P��as�n����f�4<Ӫ����uC�Zm��X �q��Men�������PT�g' �u�-l@�l9n=��1&x����V� �F����?=�­�|���du|��Q�Ԇ+���KT
��W=���c ��v_��ѥ!wR/�V�a�dg�n���"�q
��� Y�� G��u��}�ʒ)� A������cS<M��GI��^�'�U�^-��熗�Ѩ����a��fqPIb��jr�Z�~�� A�V����Y�!���+U�nW���F����]��@�L�(��/�J��æ��^a*U�b�.N�mv=�
�}��N�Y�\o��`�j���ý�O��xP�,Ψ�S��l�5\VD�-��`>��^��$����:h&���fp�12��Q��iX&y�mI����
��V]�y�|�a���jF�Y8W.��2����Ν��f]���m�#�i����xT]�hs% .r%�v��Xi9d��Q˾���)E�K�S�}�^���y%��`��l����X��f"[?�!�<�uE��3�)W�w��*�u>Ë�DO�� �h�VIl1����h�W��Rm˭������[��Jm��hA& �U�%�Hj�o7���,�'x���-}}����!�K���뚧�~���DJ�y���.+��b9�v�Rd�7�p��)ʡ��n���Ȝ����L~��
pv�3���8�;��Zk���[�ji���q�uf�6�
��P�a���j���1�y���"TXa�o�d�\]�;���@sȽ��>ؙ r�,��صq[��9A��ي*�j��	�ѥܙm�) [J	�� �.f�~�Z�{M��Ѳ�E�|4�aK�L�B~�L��[aA!! 5"�
-b5�:����YM�K �@�-RL,S�����M��������>uE6H󲍛d�Mq#
d�Wd�g�Z�yf
փ����4��`c �|?2�-s>���]v�C\B����0�-_W�H�n����5�u��z���$����{k��눎��v�	�2<��`6�;�ɤ��9��~�N0U�9�
�>�T�z=�]S�D�C�x����T�����Y{k��ǶN�ˋ1��"�F��Me���p,�����L4ݛ'�=#�6E�?SL�#;If��*"��~�+c��5x�ol�����T$G;�юv��_;���hG;ڏ�F�"� {J ܝ���憺��C�a���������������n���N��A�8B���dVW*r�r>o��`�y�|}��ݝ{��Y É@�{�w���j�`�Y�DU5�͙������	���j$Q�P�a=�K��#����l$JH�:	��36�x�̐�4� �Ơ��Nw
�����D@G��=�ICM+��0����2"�t�7>,"�EU��P@���ڰ�˲��V���,���v��({���"c����X����6#�`�4���ׯ_�;-C�� �+I<�  ?C[�UEz��z.P/ F��R#�D�8�;2.�X!�3���Qcd�U���;+|�e+��]nu��mKn�������t6�P�80�H>�	���Hi �z�7�� �*ӽ)'��Pq*f �Cœ6p�������a��jUS��̭�5���l%X�m��[u�B�+��<���I�Sf�8V'xAe���9�r2�y����T�̍|Ę���4��
�J�s�5��u\� . ����U޸ʨ���	�A�XB�L)`��Ɉ���<W1e�e�_<2
��O�B,���v\;004�1�5��%1ڥfFbVsN0<Z���d\ٝ#sQ�k�68>X�����ViA W����ֹE�TJ����Z/+�!Lo�)4�S���� ����x��Ζ���j������\�b���AnU�g���j���!h�UX�a�t��q�csx�k�-M����2�rA�R�6$o����;pu���t�=*?ܫR�l�0M<3�3˸4�f]8� �J"�Q�NRE� f�|���W- �J��7��?��9��L����ʜ�R���ѩl3P0�pf{�~׼+r��ň�r��>ǫ��Ø3�ɬ�ϧ2�eEAGw��F]�����$�궭Q�38�y3����g��1DX9�lj����5��K�����p��'����z�crEO2R�	'�d����lK�1��A��Fǈ{)�;�6g�R�����s[̦1�����)~JSLh�S���j1�:l�IV��������9!��o�1H� �c�g&�j�����Ǎ���T1��*奩vx����쳿�^�8�hC*��s��7�r\�v�suh�,�}g�Mw@!��0����X���Z��k�^ߓ�o�����7����⤣��6�܂�����D�g\W�aln�On��+�U'�lc���H�kP�b#������hG;�ю��~;���hG;���!hf����}���%ܧ9���-|{�F ��9��jF����_7B�/�n��N0b�h�������������%l�h�CoJ5���}�)LV�8}��&�� �rn&	> l��������V�>ϷVً"�s�70���%��g/���;UZ�-��� i� ���랦p�ܘY�)(�#���|V�GN}��m� ��qQE)����#�}�V 8A�P1r>9�k �w�h�z����'�p�Z�Ro��&u�Pq�7��nݴB����?�?��O-����>��z�[��"UO�ŀ�j�C��|�����~=�.���dO� [�Q��PX���cx���$3�!�f��̝�D]pXO<�)��*RSP�:�"��>��>���F	@)n��i
F&V�,=10 ����*ʐ��
݂k/0�(O/RC�T2op����m�LS_���4���X�^8���P�	�#�a���$�x(L-d)V}�y�Hy����Ȕɬ�*��N�9
� 	�O��7�K;",�lA�p�FF0?�^�C�iU��RPM��VMk2N��Y�0pv6P\ Cj'Ӭ�5�B��	�ڀ~��5��R4�I�D@?*��S�*��)��]�4�ss$x.�z�vw�R�G\S�17�0g��O�n�N]�@_l�~�A��@�RMR�,c����"� ڪX��k�kX���Y�q.�?c#�8DɨUf.pMk e2;�@b�
E32m�b�,�(%�E�)*�,�Ytk)#9��:�����ޭ�4��P��McV�K��#V�6������|��!'k�$o��鐂��|��)Ȃ���R���C��e��ܘ��~�<�g]���1��c]䝐��vJRK�w���sq᎚'���',��3RW�ܯq�l�L�DT��\�F�@c���P�5&��yP��]��^ld�܊���a9/@�eYj#ɕaf�/�e&8)�h��#V�o$B������-R=�[�@����c��A��H�:>�3�se�%+�y>7�:u�~������{Nl.��'��j�hf��\'Qy|fC��g�MXk7R�Z�Ȧ,Mկy4��	��v�t�d�k"���,�ȳQ�T�0(�?cD@.��W�p�N����ߴ:�d;�,M��E^��ȾFٚe�wok���WS��{�*��' \�X���*��s�XԐ�����+ ��x���ZUf=ɾ�'��3S�uT 㾄{��~�} �9�z����X<��b Z�ES�κo�8�럷rkJ!� �iŕ���
vqG;�юv��O;���hG;�ٖIU�B�.��x�v�����5ܑSe1u7��&
ne�{���"��OnK�p^�?�u�~Be���#7R���3�<`w��.@?��2pf�7w8�탔>2�ÃϹ�R�( m�X�>g���Hn��7Z��9�������Tu������ϫU�H�00�������4�;׳A�6s'XYh�A��t��J�~� ���q,a���
r����i}T�e��_}��o���:�?M	�(�JU��t�2��Ң���:7ڽ¥�]^9����++�i5�jo^�� 4����}���p:�0�7�ˌ q\�����+��Y>�O��O_	�������q���W������܇���uܾ+O�"U���B�����$&�?�u*HH2%�tc�<�ch�d�6/wV��:-��8W� r�f��^!ٲ�H�F̞��@�*�,k����M�!�*�^��`�۵�z�3 Z�A���	+Q3�7�B\�|c%t�@w "��*v|�{qk���N22��0�Ϲ��f���d�Ad �D!��o�isr��>?=�#�f�s� s���E ��d���8 A0/-G@�յ*Zs%�@3t���,~��t�����ǿ���45=�����#C�En<��2z7B�X�D�!@�*����*sa_S����@g�2�RY����}�i����D��b�D�)��3+�7�)��W]��[e�by���,�7��$%#M��	��ޯ��E�>��u�%�9�4NdC� �>wa�!�Qu�[�`����).R�ݚ}ڪ�pV��� �Yf��ނ+����;��u�+�56���d�wiF �¾�����P�]NE���e#u<g�U� U/%n�������cj�ފ	�� P��CͪI�����u;�؊pr�.��F���]����z��JՅV�{�킶,]ps.Y7z�N�%O��#�UTߏ�����U����`�z�V[��f��o�;]6%�e��"|���O���KZl|N��P���*|�t��o�m{S�4%��O(f�q�qc�F;��'RS�\����c�<�]#S+�nl1���<P+2diʵ{��Jv�y�4�%�O<���������Ә��'����rg����n��g������
>�.���S�#B���;������HOd��
uO���ʍ@�3�۽�X�H�ŊM�凨�������e�dS��z�~�::�x������V�[�}�2�L1��E<԰F�#��0�P*V܃0��L�������юv����v G;�юv���R�m��q㺑AV���{x���6����e ooo�6����b�)
I;�8�@��o��0��\T#t��pE�R&x�A�0�A��J9Ak'<��B�s0�J�!�4p)?7հn����D�&6�"{6���3��ȕ4Yh1��9�&3�+U����)<_��Z?�Th5�j�� b�j�6��t�C��U�1!( e��R* �Q@;lZX��^�:+�#`<F�!����z��,Ǧu=�����٨L7*� X04�;�e�퐼���~�m/���'���4���U7OO�@��y�Qe���S��s�f��x2B��V%�}�[����� w����K8?�C�x��˱��)��Z�k���������L?�����s!8�� �p�O���n�2�/�׎~NȦ�m�L�N��Z�n�w����H�B��%�[ltT�J ߓ-�O�C�=˶qK.I�<�3dz������!�i��	 M83[& 59���^�+�&�0��	��.�� �0�ޣތԐb�s<�D ���ٻuHT�8�8�?$h�S�-`�����$~\���t�X�O�t K��79��b`|��ـ�ήC����ac5t�Ǻ6G��cŀ?Wf� ��~�� ;�����x�kD%��N�#�s�e�qj��KI�h��`6�-�rI"H:���è"�E��f��C�sU�M£�O ���*iw�����%-p��bk���(Xm͢:�m/ �b� �h7� u'cY�8�wY.���3 1��t�E�e��N�
f�u�I��3�;Z�y�7�m��k�hD����b���)v*O-���`yG���(�����;0%۸�Y !� ���5���zȹu�-�&U�Si�j��Q�{���F��.��3�(�y�NVs�rG��q���Ѳ��z� �5@�Xz6�M��=���ǡڟ'����o ,����Ţ��f	˴�2�]˳]w#����d'�-�&�fW椙W�;�o��w���M��s-g�Ȥ\�l�'�f���-�jvIPSe���
�LMc�N�QfQظ�l��=�M!�1l@8�>g�&���F#�*�P��o貙�vD,��;�%j>O�k�e�$U����#⥺�$�9޻����)�9���V	������y9�|�J�?����	�VH ��e��QX�g�BX�6r�H�=��9�d�9�\���N��@����yR�d*WY�����]Y����q\��ɦ¢�Y;��ҦX���p�Z�l$Z�Zn��f
3I��Bϐ�!vlRq�$MT$dNy|Ƌ,��� �2�#=g%* u���%q|Iy(@�v������hG;�ю�ô�[�ȰfT�����t_hA���`{o�T� ����
��u�js���zCU���NA�C�gV�-K�<������뀊8�|��� ��9o��V8��$�G�^7�us>(��+�b��~ݼ���������/��޿�o���q��[ 8N#�Qn	��`��1���D�c��������(�
Un�{뿅�� ml��7nH�[	_�Bb��u�Ǉ>|���������ub�JH��O]60U�.�k��9����w�f�t��	��������� r�sDE9� �a���*�lh[����L�g�X�^��H���GU�2�4��DU%i/�ۃџ��	J��R� ���&�V�����{������������瞬*�{M5��ӳT6U��ixb��rR���K8������X?���D�?�������=�����H����K40��U���]!�'������sxB���I� i�8Sf����>��l��J�Aa���n�
�U�:�&Ux�ڂ:��& �3�_�d�ိL�����'n��iPe7B@z1�#6+�Ώg�����;�i�
bl`��	��
/��y�b�r+�dP��%6%? |NX|�����C�S#DH� �����j�QY�U�f�eV>�$�,�c�R��2E@\2�1��с���[�q���g'l��5<<>�u G��]����_���㈋4��*Ϡ���0�qn3�~w�L��,�0�iݖEJ�v�: ;#��,�A���L�����,�ee���{�å�	�{��bD�@��x(< R�����ro�YVP�Ӳ��"��"{B#�hQ՛oq���	v�|������$B"f�o��< ���0�4-�pn�6��i��SB`����.pD���\">��5 "��"!�~�b�<�S�#+ET`��67�g_3#6�Uݮ���y����S�#bI�HE(�<�9���S��j��޿�j�z��ln��(F�w]g�F1� �xWnǽ��β�� }1eD���s�4F���h���
����Ҳ\���ٵ�0B�Q����]vUZ�ʙ����ccl�����-�~Қ�c/�u#g�8��7�z@[�j����Ta�?�5��Б�Igf`l�Cn	ER�/m�¼ur	�">�r�։����@���H�$T�vl���-����#G=+���$l�d+�� vyG�k��+���eK��9O��?H?'	��QU ��*�U�$z�/� �	S%k�g�$���'0؄ի�F>�f#mH�Ox&���)��DA�<N\;I�{?ٹ1���[��<�-��v��F<g�n;��A��J����φA�<-���-�i�C�P�LjVa��т+�} l>�T�}t�T��و������f~vn$�
<�? �κ�A�������pX�-��hG;�ю�;jr���hG��������ۺ�z��3����"��~��������=}y�����O?�����5*9������	)+������r�����j��nH���\� +r +�y"�ba�����v���
��9���EV'>>��O���q.���J��yx�y= o/o���H��D���ﺁ;�&��Z;�r9�B�Kf�R	�e�1�OWV�a/�>�P���+�	a� Z�e�Ҁ!��C�w�%��wX�z��F.�}�AMX��|{x�����?�o��.�*1����B�|�B����CQq�-`U�<~���9���. �n�����ˉJ���_�g��������~+3�ʑ5��9�I�Â����o���3�`�!T	łJi� g헏�~?�֞�s��ϸ7�O��a�M�bBz��1_�l�0��ʭ}��X�	X���W�W�������ǟ	d��k�����$���\J�~�hw��U�{�G�?�����z'.K3a|u1Ġ���"��|zd��<�J���B~�}�m h��A� ��|?T�;���:G
U7R
��q՚ 0����eu�3��`)�6������D�΋U���z �_�Ó��	������4���9wY��|���oڠe���6 (bRuf͑-������6 �k�Ğ9���2��D���I]V���6獜�u�a3T1�� Ԡ
�`J&����6�?����������u��:O&�>���m�����$u��`�����\���W�~�>>���$��u�El�c < �w����Οֹ�ex�5�]ϐ�cp]��	��z�P�dE�p�� *A��V�g��S�	�-�d��ױp�x���vał�G���_[V1^�y�X�/�5�4��cAϰݪ� <op�fh  )TcU�@h�P({%lYu��.�s!}��g����
҅ǚU!oa�g�%��|$� �qq�,�` w�A����	D�D �:�{�ܽ�a�����|�����Z��Bf?C�0��M!��<�-��U[1����,"k�S�W�#�'џȣ��G;������ܨ߃(�!�82W�âl�V��"ȈS��q1�[�<�J�W�.��l�`���
*�6tf���K���c`~�J���
�)�:4�:
��V8��i�;I��y���<��x*�ȋ��$�Qq?d�;���X��L��,?q��;��^�>����N%����YD���bP
Rf��b�vh��G� ��(�F>��s����X�B��)
CxKCf�:O�g�����c�L� "'�� �1�Q�H]#�|=G?�x"�ܯ�~G�C5�{Ig?ǺB�*`Qj��n}��Y�i=d�N/�'���y�d?�yb?���cgj���I����_�,�x/�3QN�2k �L9w���V���Q�#S	�,�k˩A_�f-�t}�e=>��-�����y]�T*�,�Jk�<t�M�?�%�A�3��T���[���펹�D�s#բ\�;�:I\v�<�юv���N�A��hG;��~�����|
3@�u���^����O��J7��x�����矨�8_��|�Pb��OX7@gV��x�~l��iOt�_��>,1��Z��dg���q����H]��aID  ��YPH6���*�E�_���iT��I 6�?}��N�VŖ�τ���	�X�d�X+��� ���_��b���Ī�3�&�k��^�y��v7�K/��@��c�ܕ��lAlh�ZЉ�)��ș����N���?=pQ��Xu_�ζ� ����S����	b?}{����6�!鳎*f�>�� ��iY�&������XX)�Δ���L�gQ�U%#�U�^7�6�A���a�|6��Z-T{���߉볾�y2K��g�{�W���/�ԧ�O�y�����ޯ�un�����|9�����jf�xO(�c��*} +gV�K�4��R0+T�g⦪�����>���l>첯�Jb��Y�T$�Z���?{�v��
Jf9$�^G��=�jU����ֺa���T�m�%�?�j�kHL��)U�Ss�j��%_X����czy��л�G`ld��z�sz4K�`l)�V˭�hw�wmdE�����-b"CkE�	�."+Ub��'K�.[�}U�C6�b <���S��E�T\�T"���4�$����dk�p]0O-�~�0�6c� B��f�
wSA}ԥVq�i���T!?��|�L�#U�^_�����@d��J�� \���1�,��d���c�
i���s��%lYQ �1n�eu�z~ �I��v���|����C�=a�x�@�1��q*�&y�Bg�� 8���檂��#I���՗r(U��+��[P��`vt��uN� ��d�A�&�o�[ChѕD�t�q��ިFp_�Ki;�p���$F���ϙ�n�)����,�5h�뒢�2�J���ɋj��]$ç��ϕU�fM�?'�W}�T�Q�b�,�=�P� ����/����r�����k�N�v��/N(��JǤ�ܫ�n�0����0��9h�\C�-��đ�Z����\���A^%��T��b�ę�l�0�jdS��1�x։rP�B���2*�|��>w]�{����G���^m$��FT^J���g����!-ܬ5[���6��Y�l�]��r.p<���T�tR�L9E�;��:����?���gM�o�~�א��YJո�dy�
�^(��6vjڔSP`%Su���ye�N�ؿ�y6��Űz��o�"o٭G��K����ZNJ]���<X��pͷgZ��?���?������ �9�9*P�����<XC����iI�g�����hG;���юv���j�6�|X��6�k� �����ŷ�����M=������7�#�z�ޥ�X7=��������h �Q=0��o#���A�E���0�f;���U��%��q�B���JSUJvfG0qs�P�F�j�>�r(���x�����$�����Lr�iRs�|����P�|�ΰf�`'��Y� ���A/�C��qQ���G���8���h�#̕ ��b���vP�@(Xn�'yey;{�������v&�N�l��/���z��.<O�X�@�� < /#J� B&�SI�`�φ���!��Y�����;Ke	~���뫔P䁶Ⲭ�p�����t�͗��߰ݺ�:'�6�W ���>���3���e��Lk���g�@�Iկo�oT�{�"#�ݣl�0Ǌ����i�*�1�1. ��P��E���Av�&@�o������`,m^��m 1U-�;K�e��B��q�|C�׊l���{Q� ��%��WU*�D�R�������b��v}�W [q�<�
���׏��(�N|�:f�5$��l�\Y�q��Y��3(n��8g��$��/X3f�����Q��Z�s�ڑ���/�T<�#x�#��[�E݁Z��Ho�(�m	`'��r_���&�5�����j���fm��d���_���M�C���FF���k[4%�fE?zS5 c亿����N}ܬ��R�8�ذoiY)cA<X���,%Z��$k%o�)�
�ڬ����f��l��ȟj�>Ŭ_�$���~�h�߁xD�t��n1�2'�gΓb~��WHf%�]�,�Υ)�x��,�<W�,Ǡ��UY�9r:uvoTp0�-׳�5�Yw�dhU)��XY�ވ�j`�����[�7�$��׽�4z��d�2�?Ϙ yh߽��h�2�����H�Te��4�u�i��4�"�+�S�2_f#�����$���,�kGT��O�B���s���+σй'��\׸ޛ�I�s^��wL�,��Ԍ �s��xvꘑ�{���cB�0�Py=L)�9�B?y����'�S��c"�m�\���=�-k#��y����R�V`��^�$�ȶd}�����]��3��=�%� )�~�J�P�=�0�i]k&�;�X:�����x1?U;f��k��f}V��5|�c�w߬�jn� ̃�֬y��������a㰘\62"�����M���ch���HT����q�{xI����G�fZ� �kN�Mf*H�C�k�����n�'k4����{��ng�̮9t6�P���k6�W�e�
p�=@L��-�&s�����hG;���юv���i��h�h�e��zx��ÿ�ǟ�/�}�f�v���󺱌�����*(�������Ǜl<�y��[7~T|��M�[> ���ȋ�ȏ��̫;볯WZyt�*Ft����=$Ky}5�oZ.UU�SnŘ� ��+l� ܗ�B�#?����&��B�� ���8�6({��c��E0;C���0�B�g�����1I/�keU,��M�,P�+�U6���ח�VN'�[7����)PΊ�E�B){K��@R�+6#���x|�
_�k_��`e'<�Y���������^`�O����w��XZ�b�W�0�� }V1��;��36a��<��+�n\�"�6��������/��
XX�̬�����i���$U��Oc�������w��`9�?��FU�.�=,V�K��:� #;%��+u�n#�`� 39 ��~�~��X"9� |�PRz��[p�>L\�.��S��b�{����lU��[���!@�S�reWAM0���u}�p̒ /�_i�Ki����@�Y��X�9b\~�������F��0�̃��A���nMY唺�� &F��. 2=���D�y���K�4'���$��^�:e�\�nM�3U�g�Pq ��B�c�g8B����S��a���^ͺIn6,�^D�z��׭/Z��.�pg�o��\�*g�v[`�<L���z�&al�dr=���#��'l�CŲ��^F��Y ��)L(�ll�L��%D0'���؝���@�f�E �D�뾂_��9m����
u̱��um �D_�\�XE�����X�jq��~Y�'eϬL�?�N�!���cWEB]h{/"@md<���u�$�D�S���@w�;���5NV�m*�����d,�X�ȡL/��[�[�D#��6HP���b!���?�>�U���k;�Q�rk'�9���;���\c��.����&5��]i�!�D�����v<�jz��*@��~��6c;���qUV��`�8*�"�<d�!;m���A�ɷ`�>,ԘA��UM�7�"�# �(�7�9�g"�s_����l
*T,���O�b�
N���@�%��k�K�c����ň���,���R�!u�Ƀ@�F�e_����O!�ݷ��࠹X�`��q��fi�9O"d�۽�rF�q7�E6��R��Zf�ےhT�T�M�mn��M�2������H5HG����e�0fFi58�OQe�b{��MTa���m�\p��S�4�gq����.~�ʢgm���m�M
�������q�5�qZs��9mugKx���hG���� 9�юv���p��vo�p�]X���_~��_X������뿁�����)����C��������죅�U�c#4N�0�Fn� J @��7���L �@*&�ֿ�Z��띕g� ���vp\nwD�n��.�I���u��+Ț��RT�#cd��l7 �/tPe�|!�G�y��J��@VU<�RT�6��A*4#g�Gzj�G�}N��y!#�s=�6ZYa�� G�o
-���Q�T: �Q)
p�j�<��T��Z�8O'n�ieϴ"�����������7��K8?\B��yZX�vݒ�u��Rx��{g��?�����V�^i;Eb"� � �jB؁�V
&EX�	!P�nO�h�����|��P��*��R����&?w'�����NgXO���e�X�&�l��g�f]���&P(� �H� 0}�`ൃ1�2*z-b��])yhY�	��9g��Y 5�+���[*�F`l';�E��Ed���,w0_��3�̤Ea� 4��w�H̊ea�s	J��%�[�Sp����d�L똈Kjāu �@�0�Ǚ�
s&2�M�,[�� v�s tn��$`* ��SU�Hœ#L>�� A�Y���*�O� ����U�w�2g5/澩�8*���I^+[�"@��G.�M��Vh������[_4-�9� g�H啬hXQ�j�a���V� �Q�=NLsS�ȧ����#��\�I��#Un}w��N6��EFōj*d��j�.Y����N&я>���-�h�e��FN�,��7k�RÎ��8E��l6p$��Yш�SV�m�����F	ǃg��V7��@�"�$�����:���a��>�L����g�2�T*�់T�<�-/(q�'ee��J�,��P�M��X�yo�| ��A�n�Ə�����[)�TQ�V��9X�� �(r+�M�"U��Ј�7��ǔ�ae4 k���
x1��U�l�������>:�Ɍ@rDQ��`���n��q�Q�1G~fa�~ae?����Z����~��`�;l2�Yq��a��9���ެ�c�BR�:�z)lp|#H䬬�]wJ���F���p��G��w��³g1�I��l�ZRyGf�8��1r��ָ��.����H���I������s�ETdd�u<Ra�_q��m�;iB��l�xo�xQ��J�?  ���H�3��j�V���'�_�`1*묞k�
~�v���*�M��S��6�T'�ޞ�d��wX��T��72G� (�(6�ٟ����r������ОOtM+I��� ��m�J��e�gaCnַg�o�|�brُ�Y�F�U�ckoҞpĺ2_����4T�꛸�5���	���qG;�юv��W;���hG;�����   �uݏ ��������?��7��H��~3����/�f#	d�������F������BZ�ჽ�,�������*OV_/��&��ť#�� ���@ћeuX@e�����i��z"�_�J�!��;���cΧ�I;�]ö�T �$k���l��!úу"�V?�4�UA̬ʃ ��`�d6 �A6�wPb h�<�i�Ċ��;_�7f�8��:o!�̇0�f32N��X���S���__ÿ-��s8�O����rA ��.��Y�<�d;���^�U�;�w�
J�j0�4��t�p#��eKc�@�߲�41�o���by�W�d�wo��>��ǆ.:�p�»�׼��,ˊ�J�y�	'�i��E���� �"UN#���:�gއok_\�A�C��#�UR���X5�$���^uk>� ��qP�!�V%N�����>T�@�,D$Ƚ�����!ʰ�B�>,�2�/K\�p��f���{��1�؀Wgೇ���

a��h�"1��C5�_��N\0~���SB���,���*�p���=�k_���z�~D8,�եY��X��ͺ(Y3 JW�x+f�6d��fV�N�$��l������H�s� �l��� ���8 �c��O6 6�-@�yW��Jy��ۿm����,;@��i��w��ހ���N$,�kS"�8�����N}�챲�4���`$H;ڊ�RS~�.����>�R!�^C�^ӝ:S���ֈ�I�&��zwi����*��7��	x���}d0@#���I�*�$j�RS�tF�s��Yc�d�)�F��*r��a�_W�@�R}b��:��Pf+>��v;I�!֨\>e���蔤.2ID�-�UĶW#x�- 4I�ei�.�Rt���,�W����������ap����#D\M�s�f�$;��d��`e���=�Ն����O�0a|'���9GC�dau���T~�$D1E���|�s@��� ���3ַj8�+X�X���H򠋃٫uf3��紀�^,�"&��y��'���^L���������O&XϰƂ8�<t�W�﯍��f��)�Hl��Z>_{����0��C�*���ئN��s@2�)�i����z���Y�Y�8�a�(�ڧy{�p[,,Ѽ_3�̈m�E�S�Ub��K���(lr%5ua��g �*�C���Wu����m��$�:_��6�_P�*�<��D�UX
�|���/�I��������!��9h��1���U+�᚝�<���C3m\� Ҭ�}�����H�yP��|G;�ю���v G;�юv��-hcs��/�������A=T2���W �����m}�De���L֦Vؼ�j�B��)[�>���4-�%��=��5�����l?�-��-V}v7�|Ba��)�t�^�7ԗ�E/O�a������կ��@��]U���(��6� �n��ϸ�[{�̸0 �̕�q4��fyЇ` º�N�Ї?�L���@rTT��+T���1H��6��9 H`����.��t[����3��V�k�{�h��^�@A��eV�lE�3A���J@$���wJ��1��ƽ��p��Ԭ$T�[�M���|�}U�*�I0L�^���cL!��~�� ~���C?t��?�!��>;}}�����q#����E����������n���!�A��/9���$�-0����N����w�1 Us�I��|\��2-F�Ȟ��f�rW�35 �X28DB� sT}.&�ۉ�����m b��x(D�o�W�E��>�����Re�B���$����vօV���,�u��cZP�c�AaI�c_6�|��A���U�P��^sf�7�n�-:G��)����ҥF���q&�_��Z-[(��Z lR��e���i/T����/� ��Bm�)�,���S����ݾ��q�����yWB��ɖ7������[��TނD��fy��Lꡰ	�,�Ec*Ж�� ]�SD����h�2 � �u���'a�*i� �Lte���0��vR���!5@]�VI�6������eGvl�`�eI8 �q
k:VNwF�b�d�I�Rj�I�.�*���b�z���>7��ɼ��=  K��jqE� �ɲ?���Ⱀ�� $�1��w
��ӳO;��� ʎ\x̼�>����S�Lݲ�]8��1�ӎ��>�Z>����3��r��߮����?�����v������d��&3�%�
��j��~݂��O�-Q2���qr��r�A���+b��g#`k&�~��Zۡ��v�3�L�d�2�VFk�Z+p,�[A�?�;ȍ��I��F��ڜI��N�W�,�Pp�J����MN�p���&~o���>[nPfQAa����Jv���>��ǁt�Ný֘S���?�hc9�"��'2mo��f��T�uTX�|̆O�w;eBk�k�.�Ǝ/ɶʎ�K�K���ZG�,�
W<O��T�X��wo��>#u&e2~�kn�3�9Y�y�=#ҡ(��+�+�A@���A�n�ٔ���	J庈P##K�W��b7�� V}��S�$E�q�gY呤Y�)�i��]���;���z[�V{���hG��� 9�юv���Pm@���y��+T1�n�~����¡�[<��u=�Q!� �����
3"�VJ�b`8�J��qe ���l��%����Ue�m��&��yІ����q�ڀ�@��@�ͧ��������M(7�7���U�ȿx� ��׳:o�Mˊy7�|麁����{Ho�r`1&�
��FZe�*	��[%/+�-T�A۰7�)<<�����r������ �.�E��ķݨ�f �Y+}���_~�-���pG~]?�ط�Z�����cݔf�G��`���N��ԫ�@�����>o��E�m0b�[2@�0�\�� c�����a���!P"os�V�j��<�9ql,f9�`����}Y�����H�Ý��M�CػQ=êי�y��:�xb55�Ǒ5�ߨ������)<}�"��]d��A���J�]c]�.ɫd��,�&��Y���n
���w#�b<�呩dƽe}`�B�@�Y��]�(��_��J�$�m��w=�����@�K���Z�D:6 ׫�bG$�8\����! ��|�m��ͮ+�å��`,��ׁ�t$��T�$��a�D@1�by�+�MUf�_���8�Ւ����Ϭ�`��b�ł��s:C����fD�+�B��¬J;�CI�#�@���ẁ�'��aN�| v�:�Y��#���*��Y<;���θ402��Hy���IP��Ͳ�i�"�i}���FU��"bP����ػ��g ��"��fN���*$BwN#Fh#�x�U�cl�*ĵU�{v��<�ABl��j��0�^=`;���	Զ~���/��)��TW��c��z�P�1��J�����V�����A��i7���I�����߃�&�2�1V~Ԛr`6O��AU�7;�%(s���\�3��TnITۼ�kϴ�S�+�F#ŲY�yPS�@z���e��I�����:����g���I�UN"��c)�6uUJ۟v,��-�S�:n�]q��?+�[<7�qc�J�)�����r�Ee�&$���0gefɂkn���2[��{��3h?鯁�b�̎/7k&)�*	�����|����(� i��|�q�p>�۽���Ǉ���5~�L�-����V��I6M��ѽ$5B��E�M1��L-e䯈��P����P�F���*�ܬq��,�Y��ADPL����Ww�����~�UƗ�3vn�3�����`T����u�lEGx���|ϼ����E�Un^
�#B�5@�\�*q]gPȲt!O�=@U�Ȫ+����B�:~E�m]������lWS0"DD�`�?�]`y��ma��U���D�uT�!�hG;�ю�;lr���hG�������7��`3�1�C�$���6��^>Hv �
߲�>{Y!�oᷗ7U��oj �o5�8���B����6S�f#�����9��>��Ъ�r�l<����U�L!��������~gUv�4��g�H���u����s^^_n���.��� ٨��r U���8��y�� |���y2�U���6{ T�?�R\�m��8�7�g�0���}�M���c�n�	ZϷ1��n�ܧ���f�}�u3��f��jҵ���>�M�8����>>p���^����@c�`# ^ ��˯��8������r'	�	X�� �;�TC`g ���PF�� ���~�Ģ���>�_�/��eP[@A����U Ɉ(��#W ����BG�"R���o$��<����I�z���:�( h�
�'A�u��8꼩P�����S�;�L�u��9؃���*���*�-$���� � ���!+��\ɂ��b�I�,���O�a������]T%���}�z��b����+FV $C5:����UpB}�J�Y�n�z6��' 'V�&Ju~N�y`{1�ث��ܡ�H̞�u��d���I����s�>������+T�09	�Q r1�9�� MY�X��B;��[UVC�@�	@c�����cA�k��R�4����n��-��8�J(Eں��P@��x||b�_:�Tso�@��0{��:N���p��<A/MZ��;��Og���Y� �8NZ�eﳮ��HM'Cd�7�k���"��%(�G�W@&�ˠ`�d��2�Z�c��ܪ�ayp���ÄA���C g /���9# �֗�Ը<<�$��@*P�$�*+��"Y�x��h%��.P��/��]���΀��@\ڨ������]�u�\�,1輪m�6oG!̣��(�UqT�� n�̏�B���gA��4��+��YND��1?VKX���BP7��s;C���RZaI�����r7*?�8֬�<����Cm 5���*p���5g��i�߸m��\��Fj�5�������f �Um�s�<�ň��J��e9>>7�'�AVS���Y 2x�|�)+��un�^�"ӈ???�IS��LD�R �K_SN$w�21��c��{�ڧRT>�Pݑ���»٧dN�x�T+]Yר+�v���S��I���������|�0s]�:tf�u"�O��f}��'�*K[vS�,�����T�3��=�����rj�����nS�k�Vd���("����9̻r�^hK#\H:Ͳ�Z�������(UY���;fsQ���s�w�nt}��C�+89�������[�m��0�g�.c���K&ۢEV2�L���S�[x�Eh�a	��}m�M��u�3�l��0��S���cH(۳m)dHi�\�;�}V��Q%慱;9�юv���w��hG;�ю�C6�T�m�zlJh�	؇����b�2�ez�YP^�;cf$�h�\�	T�vny���RJ�}Qx,L��D���ڻ��,� �*��J6�s Ѕ��l����*M�H�[Q��eQ���6b#8���*x�c
�9�|�g��æSUqg��F�N��;��󊞥�e!�=fW�����+^�M`�,>�B�v]i�4�5x���]t��7�p�~������@����l���11P[���>��ά^�-���7������ ��.4,c%����BM;PH�u���*I2����PQ���x�"7D8�nvmz�͠o�:iL65�]��@�e�Y�BK
�'0E �Ae�����9�^�; w�f�f���߮�.`�
"�%�g6�j�ai@:�����B�Q��~�'�n�lv��V}�KU�
��+N��r�������9$g����S����%1/������Bӗ~���~�k�Vu�U^p��V�Y�1K(�uJ浮>��#�f�t�c��VQ'�B�9��U�\���eiP�Tu�r�g�ږ�4eU(������y�I*6?UHW��ܝ �a�X�v 6�u����rlB
(�۬iL	" O�b�J����IA�2�e(����ؓ"1�%�j	 �}�L�c����ԬpZhu�]T�#���m��&#N2-����=��<�v\n��뷩B�B�c�R�bH{б2��)5|���M������#UI��0��cl�����HSֵ�o�1��d���P{�7L��{�Y6����?��I��KqE�����/#�D�ny(���� ���@�tA�qō������EU�l���葉�hO���k�[��^1"�-�Z֍�R���PhY������3�W�x��gd&{����,��P�UnC�T_J#\IE^��]?��}�~�>�;��"��Z>Y˵�a����¾�Eu��L�y�Jǡ?5�۝f��T{`7��%�m�j�a}��O�Z��"UyQ���/<m�j��1m��x.����b����q��D��@}��ORW�T�v;�����8�!���L�����{�>��c��]N��QF`���t��9Z�|9�� �L��_�o������/E�4�?>��b�;�풴1��G&�N���P��q�=�s���hG���� 9�юv���0mx|
� 2x���,���a��83EB�������N ���ټ�����L�t��]7�� 3%Ⱥ��$wB������<�'4���n2[
e4D�.�`Fm
�m&�$���6��7{�$��%��BFDf���Ȥ���옞���[Γ>E��ޕ$ ���Y�g�X�"ڪwUf/ ���ݭ��9��{��`F2��Zb<���zu�_2v�Y�2�����g�dQ4T����De=./z�e�f`�/_~�j�8�O�Z vAV������[xC����\	�ow�� ��T��p�$P��e��WYdyOㅺY�y!���b���<d[��M$�"	��@o�u�?�ߛ�L{H'�d��Y�d#���l��B��$��{�=�Џ`��w#P�a��M����ݢ"3�sode](���,`��]`��N���FK�҂��.�S���QDI4p�nR��6[�\d=#��s��Cu���]A@����:����c�̭?��<ؕ�K�K���W�;�;���:+F�H�	hI BG��%�%�C6��b���z]�[���u��)��,�� ��RX��������"e"9���2�M�2�a�۫� k����Ș�g��sм=Q���TPͿdS%���ӿ��5�a\�S�D����m�vHk^��c�i�xǟH��Hpu�b�]K�X�O��
��������<�vf� �}"�g��^����4��a���۳
�����&9��.�N�o�YcVlM�2P�9�����5.�Z
V�ĸ=�]�����"ui����Q�e�E��j��Vo�'D֍�a����ad�w�UW �������)G�b��
+vBvn�����a�SE����]O'��,���x�NF�NǕ��#�1�&��9DkJ3�֚���uo�=�+��A�����M"?F���>u�ʅ�����u�U�wIʅ��)z�
���pK���"�;+E�$ɍ4��ă�&�Am�gR&��r��A��X�ZF���;��s_��sB�E҉X���k.BK\L=S���Y6ޟ\ݓx,�[��{V����	X��?��M�'�ٞ�0޻TP~}3��5�7�m}�}��{'upP�`�5�'��}�hkdp�b ��ֱ���3A1�LЏ�21�"5���?�p��J���g(n��0t<� ��s�EI0�*$3 	n�0quIR�	�Z�題��w��͟1��|���R��$�5�)Z�^�nOd=�º��v����l�v g;���v�_��ozQ���G[�*���������Z`��a���j��^�@,������,����|A��J� ���,%,E�,H����|>����
�w�,ssǋ/^*�M�t|�4s�蕎��˨�[�;U=-�fE	�{quK��CH�"�
�~�����[5\�K��S继s4�U�C�U�fS`�g�9�*1
U8�HDx�6����7�"��,7��2TxX���\y�����f?f��!R��܀��x6%nyF�皨�ѱ/��V	��(�\@�%��s�F���&�
-w'V�ݍ������6�-�L�5�O�Ȃj�/^���U�������a���	p���SU�g��K���ݛ��1�Bg��n�6~��_+�	�0���b������2M.�L�nS"��,���>,��b�b%���+0�y� ��R]�<-�pj�*R�x2u�b;F� T{>�N&YUy�k�B"F���Y�p��	��_/��u�X���UdEfP��Tʿ����%�t�ɉ�>;<ԑC�$���V8�����Ϗ�'�m�\�����)�9V�9��O��',Z�`����oSer0��V�P��::<q�?�9iU�TC��u9+cHH�H�*�A��I�d�4]q�v��ͽc�O��H�yn�Ͻ��>�yL�A0�F*�<�D���r_�s���hddS2%���U��gR��J��{�G��j'��)��q&�\��ౚ-��5�w�|�)�G�3�p�=�� �0�׮V
��޿�\�y�?u���
zG���c��3X.���6;�������*pkW1��6�N.8����؉X�3욙4�d�.M��WeI��pL!�{����c��9`χ�We�P����C�o��^�+��eT���T]��ܺ��W4N����bd�����"��W���׹�]��g�:��5p���w�k�[�}�����6~��?g}���9�v6Z�Y%�)�<���>�3�\�{o5��օ�xp]��s���g���#�����s@��x��������+I�p�_s���ǽ`���6�>T0�2>�{�ҁ!����T/i�t�@т�o���?�0LT��� $GQ m�����fŚ�m���@���D}t�9u"����u�eD���7P��^B��P�?v>��$��%p�lg;�����i'r����lg���w���y�k�G0A�(oy �|G\�X����jy��Nz�ٟ�v�� ِ$�of�� ����h�f.���جJ���H�楲�r���X<`��Ť�����@�m��=ąU�������cXA8�Vi��� T�r�y�>^����_-�N��*U*�F.���3z�}Jq��0�/��l�Z����e���|���	|ٝ+8�ͪ:�fUh��h�����8M��t�@�/�[��m�;oH@�fcAr��2ɣ�cZew�폮.����E�����s7����:0�T�B��"��ΪJ ;�lU���m��tB�-ί�5�&�,uY�7�k�ޏ�j@@u>�~l��q���ʲ8Z�g�uEH���!���^-��d\��� �]�X_:�T:��k�f�q����}���;����&�ѲAZ��֡�uu��@����/lr��F:����w�L��U^&��&攍H� ���>>��Z*y`;��f���Ie�\/E�^N$?�(�@#3׋/"*D�@�v�=y}I��%8�<�Z�U������h:�7 ۃA����g�g��+�u��X���<'ov�B��pr��T_��/�ˎ�Y�ŉc�9Z�:[�>���>6�J͗IbV�_�~6?S�䑓R)����x�c��֍����Yk�m�H���k/��)2�\���n��*!fG�[��89� ت� ��s��^�}Ka��Z���*�[~��/8~To�y�-��l�:��S���+����=�,��١i��1Pud�j/�'m�<ODvVX�\-(br��Z#j'/�6l՜��ү�lK�vg£~!Bc�H���Cb��%�V#�g@�m&���W�.�y�����X�D�})��i��$݌�U=}��Y=��,���;�ݤ�Z��~��{�wui���������{.�zq�d_W�Tנ/0�Ag�q���f��)K�� �ԹZǩ#0qk�b�ט]rv[NH �{L�_�N�㹮)�I�E#��6�6�����,N���t�<��!Z!��#Շ��F��s(fk�FP�8���K��¯V���1_ve��X�#�g�i�s�+�o���s��2��8_S��n�ۢ��sQ�\w���$Z��z�wxOB��s�.X5���v����l�v g;���v�_�=������5l [W���^QŹ�T�m���vc�ܝyD�MMq�ĥ���&���Z�ȗ)�/�z�gH,B��qk���(?d5e _޲�<���I�����C0�m&D�����Y��s{��K*�@�%� ���A�\�.����>~(4��l0� ��Z5<,���x�M?��z��7�a��Z���U�^A�*�KF?��$��B
��p��dV/�]���-������U��v��	@Wu;��%X%�����\ŋ�	ŀO�aD�/���½�)8�@r�A�f1Վť���
��w�m��F/*�b�i��L���,��+
*G��IQ��
$��"TXv��ܬe��|�E��6�`�	<�׏B�Cp:#]"U�Y�x�[4���i7k�gYe�nOR����Y ��B2 �O��n	�v0�{���z^��a�N�i?��0�Te��@B'R�	��r�Y>5��s%���bO�W�@iZ�<{B6.އV����ʆ�_w|�:��?�_�l��²4\u�߿1ցE�f���-���I�&���cW`�}�w��m�� ob�q]߫�}��i^�<p���7�닕Q(��1�!�u��[s��A6P��k�tr/Y�<�'�PVO��"�TIL�)J8g.�X�l�uiS��G���zp��u��30�Kd�Q�zߔ%�20܊����6;#��v��N��;Y3����_T�='�1MDps`?�0��7zQ����{l�/@�;A���T$�9��_�t��?�I��
�ߵ�M�+U����Z8H+W/�`x]繄�?O��c�T���I4���/:�h�\C�9�X󦕱�;1^�)B������ʛ�<A���QV����Z%L�� J�އ<?�󄊊c�y�kMT`x<֧����a�,\��oϥ�*m���/^F"���B�s�nC�
��s�AV#~t������~��[�m��a��u����9Q�P���,�`�y�)�d�^^-�t�y$G���CD���2�L�ў��K^K*������u(�q��5u<[vb�	Y.q�<������=l�L_ר
��d+�"�?`+�O�gK'Q�<��w݋�M��nA��?���d/ȍyg;���v�?w;	����lg;�/Ӟ��i+� s��jd�@WU��H�ﮨ\�K؏]�U��E�>Udȣ�;`�2{��x5��%�( 3������&0�AQ��vp.�h~�q��Jg�����g���0ῗH�Y|5��7h�׿���I��u�*��I��`-'}�,���պA!���U+A���SU��e7tg^<lr7`x�q��=�ֽ�/�����g �|ٮ���#�B�)� 䱋,:���dX�x�1s9��d�TZ��|! ���n�����r�VPn��Ö��
��jHU��+
��n���r���K@�%tM$Ɋ� W�Kia�f<,�
O��|<� �pMK�u��^��҅���gVع\T��mf�f��fV9���,Y�����]�-(�^�_�vaǂ�`� ��<����F�]��nf��t�9��
�L0˫�c�\QH��E�ݙ�oUf��k��a�U�
�p�J��mg�d��l�pN�N��A*l��.��E�G��C�o`vS�,�G8' �� CS	�aZh��zkW(P�R��)�뽙d(�����+���F�T�@5#��kj�O�����qo����yr#��d�� ثIq^�o�<�}�D�]�s\;�O��X����s���M6I�7���Q�Q�U1;٧" ����a�D�1z��5j^�>�OZ������X8�Z��5"Ҳ�ٍ��Q�?28��fu����|a�Bk]eFԳt�x��������9��iHc]��byl9�K�D��j�`N7�v��
��@��u��Nb �D�?#�`5Ih����n�g��|��� �����r)�<�ϸB��A9W��@ �' ���O
���m75�-�ڭ�\��s�`�����Os`���b�~�R<��<�+���P �y#_�N�J�ߨ�jf����BW6NmY�a�����Ґw�{_)��y�,���r��7˵�&k�aa獄R0z�	�>�1���i����	*b͖u�+�	�,m����q�ԕ� �y,L�~�����X>E����T��{9��`	�]ٜٽԊZx��$W�Rl�g)$^��g��iƈ��g\�r�z�f��>~N�U�N+�X�~.��-���0a��@â��I5�Jefk�,��L�5xZWP�y`.�p�vx��rrc�Q[�5���^4՞����7���F��,>=��lq�ea�	w7R�9\+	�c"�sYd�����/��=|~>���v������N�lg;����˵��}T&�e`�^C���5�GP��s���x��v���c�C;^���%��ٻ|��L�^I����|�D�v�����/���`k����W�4~�b�#�$S��ق��~������U�"  N'fGd"+������<��T��⸃�n+w ֏�Y�Y$��?X��j؝/���D^���� �H�x?>���7Y�Y�8&�X:�ɲA��7�6&��-&�ڑ9)���FP�j�,@Ace-�[��M�,�ZAԭB1{�~"�b���]jP�Ub�&�	z�0Q��
��)9��'��]��?0�����1f�M��0�EJ�(˰���ã��mfx`F�P��U��q����C���X�
�'���卪���$b�8�&�	��Xi�  �
�{y����A��ۍ��� �Ӷ%��Q~�Ȥf��z��U?�F�%�+]v��֝��ꤞR&�O��T6Ѯg���1v�A�F�
1��W�j�e���2�T��;�p�E�S�	�B�i_%�sđF��c̪��h��r
�b�zE1�7xj��\M{;�D��1t�n{�6D粫�[�fA�N�gN2`��84����S9C�ò�!�e�r4�'��F~��Q��.AĊ�- �&V<���)1�U��˺~H ���Fն�R�*[�#�,�v	f�lnM���  W�VV��l7��S1�6���:Q�*>�-XW);<x�%���~?��f����Y�� �z�<�^1 ��Av��I \n
济kl3r/�����d4���ʭ��6��o���l�u��A6��*�َ��ڹv��n�����Xd�ɨ���M��m��x~�+���&���`~�t%�T���R�M�ٯ*)���*�U�ύn���0��נ�fJT���=t�f�)5�Uʻ5ۤ�c=AW�����Q'm���YTt?/SC"����j�>�z����!LZ�ך�*�qP!N�#�WP��^��'�1������C�X��eRw����~�˵��!)GE!��"u*�"�<�sԵx}|?_Ã���C�!γ�_��U���?5��F�h~՗�*���|��z�Be��{�����ث��ǴZ�M'<��;����D�[^2�f
��س�����&�!��.8AԭE��EF*j̍ب#�N���B'ߏ=��r�TfD[-/>���i��%�ߋ\��<�.�����q��"g�?l<���OB��v����l��m'r����lg�%[q;�_x��9�����|��]��>?�ě���#�i���*O�Ͽ]F.���ׅ/���3<A6/GO�pp��v����slj�ڗ.�G��x��\��,H� ��
�.���b���	x���W~?�y�`�>���rp�����H�]��I
=g�q�o߃�������6�'Ç�������x������y�|���̊���WfyȂ��y�ZVb|��\�X�^���kU����N�
���x��`�X���%;� uY��71L ��v! ^����@8��Vg�<��%[@�UN�1������I�/��q^ �����`!I���,�����I�۷�O��t8���S��ǹ�`1,�cߤ1A+����A�W���R-� ��l��E�k�(p�����Of��$밪� "$;�,Ӣ�U��h##Px9Ɣ��Q��~�:4X�2�/ �A���-�CuESN��>~|r>u[�,��cI5�1Y?�?8�8���=,Fd<�ղm��_� �9r|Y1�,fUf@���_t�I�c#�I{��u#�'�ǵ������ �������H2?��?��r{���%�$��
Wl}���n�1) �:1"�.��1�ѫe�c�qc��s ��E�"s̍�?���q-&�?��Ǳ���'	-���x�u$���iΪd�$`�uB�>�Qf`�D������Jy�I�a
Vy-Ŋ�*�WP���ztO`�	�uK�N����O ����Y��g��vV��k+�ZV��Ɔ�j���$��(�j&*C�_;���h[����yc�����[�t�ҩDUq���Z�2A�L3��÷�Ud���p�PNj�.Z�y�O5e!�@��.φk����N�r̅ٮ��Vb���'ylT�d��>7�����YͬF��0 ~��8����osܳHcɫ+_��]l����r��Q6� �J��1����?�� w�?�/�Rs O����
����ݭ��\���%���aD��g�C�8A�s�X�!��*ۜȼ��z@��l�%u�H�ŕ6X+A���?c,Q0 ��n��{a!x��O��Z��j�|����X�ST��A���u�	L�x�-��7�g���F��^˦�tB�'�u�k��VEz�ʯT]��6+�+��B�w�C������|�3!��v��1�pL�[��cַ\c�eBA���E�UCS�\/�ᤙ(��z��6��aW�K񈹗[��u�D��w�γP��T�V���=RR=�a� x���B��Go����K��C���w�s<3�j�|�5-�.�Ea�>[��� ��2�a�ߨ���^n[���� 1+-�q5��{�Plp@`��s�2�\��32����(4j�>���ǚ��>Y��v�5��o�aKv����lg�s�� 9���v���:�W6����J�0K,��@^v�{[ţ@�Jp�J�f�Gx߂eO�@���q.|�IA+ Ԛ^�>��������n�"_��Ǩ߃)FB���ނ�y���?;x� wT�gS�$���-<� U2�� [�D�V�3���T-�KЃ��9��3k�)���B�%LD=�1�:�*�Gxo$P9���g{{��B)��)�HҘ=C�"��N��l\`��l�^�+�^r�� R�=����� ��H�)�E��cĈSΊWTz~�@�^��0��B�0��Pک��O��j�H���췛Ȱ��	TL���|o ����6fY*$�ʱC �m��T�l �n�}Tm�xɞ���D����@���~ٷG�����bVR�4���A�A����0��_����<�nI����sO��Gu3��yy)��+PL��A62��;t3vW {��,HF���m�8ͮ��~XEs�Pi��9N���܎d�
U��色j��gV��C��%�e-�b̓��x��w��W�����%�`�J��~/W}�`U?sh��vr���[sx�ÒPvT�G�l�|�侒�� �dd�4�����/b����m}�Z�m7@�9[���F9��M^��5#R^��?��r$��W[������MIe��yiʕ��MR�SH�ƽ��N�$�j�,��fP�vc
�̈H2JzQ)l��.�`���Q���qic�>�Um>�G��+joT��^��M9R�bJ#�DSIy@z�kU`�־��/ܛ�HpP�C��su�L�""N}F��b��)SN=�?�c��LB؎��=�ޭ��+IB�횝���n7���r~>�����ͼo'"�G#%wB��9��?����yXn�\�:	����t|ɮ%���&q��>YnTp��sb��kvN1r.��r�YN��S��i�}_���I�\�b�ğ����4ǜ��fl������l*��O�-��a�XM�򲝨�Ϝ5����K�K0E�o��D2K����2����9阶���XV�lnU�K��h5�9���P���$G܆*�>G����~=�%��d����f&�ϸ���>������������&?���nW���$�f+�L�Q=Ptut�В���lg;۟�����v����ln����j �^{?���
ƞ}��bi�����U�����]���UT��K �`�9��l����o��Ĭ�`@����q�E�E@ұ�0�2p�uS�Bv*���/�Î���u�CF���B}��� ��MU%=6҅�WU�'R�q�<�A/�[������g�=N�g�C��mP�x��5w2�C���H���
NV�#�"��@p�,�:/���I@���+�3�������gH�DS�H	��yģ���
�z�8� ��MՄ���N��)+�Q�x��#3F�� x6V�{�j*�	y��V�J��:�/�>��jcg���\���>�����]�i���P�1*\.>q	@E��~n�����.�C`\�9+�c��a�/��m��"i6;�A��Fg���Ќ��vMв'F�x; $�2 �~&B��m�h�Wu�$G��r�O���9W��\�m��,n)��Y��
kN/"�@�hcIB��(�ܿ$��T��C�J�8�� ��nLv|f�-mX���9�Wy"N��y/��������{�<+c�c�w�b eL��12[�|�^�)����`K�᷂T˶G�2"0Ǳ7���2,y�m�Ŝe>$S����6�`Y ��()rX���z������y��
b��)�ٮ���ڸ��Ы�K ��A�2��f�dYG���ە$��=�|�����c&\������������*����ޟ���gx�X�x��I_)����F��f���W�x[�l[�[;��Y1n
�}́گ������(qb�1�^I;�N�R���מgx|{�6X�w7PX�G~�{j;��
|s�WR��?�y_�w��f��C�� ���,��D_z����eXnA�B��r�rh�r��R`d帍��MvP��Xb/��燲Ӫ�E>;|�����i���q�Rۜ�����Z���!WK_[�x��$_����y����H �n}��1����~���3���k���z���`O�5�����(�?����Tq9Ǿ�:�,���_���m���@������yъ�������کb�y���
�VD��:��	�C�P�c��=��W�lg;�����k'r����lg�%��V0�|��̍t	(�g�<���^&{2�_���gQ^� �� �=/fe�
 ���C0�~Ru��������������}�K�=Ŗ��B2�<���_�f�B��������&���b@�����o��T,d����/&�|LX����P^�P���O�P��w0B����m��JM|���v�����M���..�щ��E�*݊���3�!t=ݤ8��`���`�[5lv���V���ʃ�/e�d��N>a��V�������e�~z<�
q��I��N ��X�������x������⾌���xax�Y9���~�b�����2}�U��R�$/�:8-u� -p��]d}t{��X���?w5����іc�8�1�:���t�z?��S'(АBk�e��n�.x\���d�2��j�|Su�lq^���������[_k�Z��(���GN�5܌�m:Ij��=����U�l	�g�U�>��Y�m�y���h�t���D8�ꙶdǶė�~��V[�k|7K/�ޛZ�3UT��*�2���Ν�X��C�#�.�N�a=U�s�8�?�?�+	�K��7�9[�x>g�Z�C�r��� ;���������+x�=�㵓Ya����"	<]j;i���	2mKj
Ǿ��մ��5K;\.��b�IK=WDa�
�LA�T�������:��氐�탄�S%�\u���L4��v����M��ٹ�F����{��%��'W����&~�ئԄ��ַ;�B�$C� I���F�~'�P\P˸�L��*�m�,��C��*%�Ô3F�I���/D��﮴��k��Z�1����3��Q�FS-�<o��D�9"uB�<U�p�,VP��璴EP���1�-#\9�12�|�$��}�����v��5χ�
2�ʇ�����3���W�<�8�QEt2�	9SDN�B�0É5xGsw�פaIڏM=f�~v^i<GW���U*)�y����]��+m�6e<��VX�g�U#��K�rw�cBۤT�Vl��/^�`s��Wp|��K���z����,��)?�L�ВM�S������S,�I9E��o��h��sE�>)kj"��N�:Fϑ-����lg;����$@�v����l�NCQ}��>��B7ب@�+`qjY� xy'�Ik��B$4l�/{�P���
KC�g����F�FP������`����$��]$�׵-�.�g����Lm`�)�2�%�֪�rfYU��p�2��m��i����B0�b��ǟ�C��Վ��O��E��1Q�2��\��a[�={V
$_��ɼ�ч�|ǉh��Z͒C�*�3,Z�w����xS�U�Y$��;s���v{�cǗkTM'X
-��f�30�G'�I�h�-K�<�I���x��VJ���L�?:����'-"�u 8��lu�Tݙ� �)[��s �@xW��J��cǗgϗa��)z�����MV�3���l��X�CY$ �*��H*��X�.�Ų�և�/��h�i���8n���úca���1F���q��uP����G�n��/�jY	�i �g��	ɪuyS�c���[rBB`��@�l��'A���ʮNhf�4�8j4�ɪ}' �$S�����Pf�{�P�s �����;p4,Z�y�����B�@wL�J�n�~^������P�� x���3s�ro����!^}>+�:xZ[W��*h�WndY��������A�Qq.�o���#�0�Vٜ�tU��[���F�R���J$U1�����w�*�7���z%r޺��vJ��ͽ��޳Z� �d� }5/'P�'!N�U�ry���\�p����t�%��<�u�55�!��I�R^z��߉���Z�Z {����jQ�IkBJ</X���0y.�T�)t�l*P�2���5M�����׸�j�ݫ�@u��3HXl��<j')~4O���0����w&
�����S�+�]1�5t����x�,�=!ΣF������t�>$/`�|-?G#?�z��#ZaF���<�5N��r>��N��N"��W_�'���Tׁ'vo`�w���<�qmF�}~T+Z��	�5�'�#2�M�Q'�}>��堆A���R�u|�U=W�\�����pnr��¤�L9�����exM���A6V'K�YAa��X�-�Ɵ�qo�c�g��>����q+d���G(P���y(�9B��N\y�us�5������_�A8���������=��lg;���\�$@�v����l�T��Ù���PsT���`�*��>�;a��ի� J �٫���K*������$�_���RRQp[ ��%Z��.�WU�Ό��8ޥ�4X����B��23;��cY�a;��_�g9_-\<*���^1�x�n��k�]Um^���Nہ����a��&�Ie����j�P��ߡ<�i�-8h�
�o"p~�H`��"�[�Y��[���˰�*�w����tt�jM��k�^��I@�'�st{ �i���<s
,��{'�@,5B�b6kS.��S52
��|1+���ɒ��\�t�E#��$vX�([��rÕ�����ύ��y7�B�\셾�:���|	,��c7P<ٱ�2���}�Zh��S~FSw$���c;�Z�ɐ�D/���Wo�c�K�A�y=��mED ��� ��6��v����
쫙@�6$?�ZK��٬bh�R7#/�Ϭ�*�G�0���z�5�?Ȃ�q\������L%P������6�	��K�y& �r	���լ�6r�呧���r����;U�cP~Эǂ�YndNW|���H��R����࠯E�gJf�����4�P��Z�a���=��֡��x�Tt\'��o�R�����z&
8��qj"}��{Z�t_� �1��l��{�L��$�� ��y
�9 ��'�����:O��en�������>���݉�vx-@����*c�%}�L����*T�.��\����g�>&K���y�{��Ŷ{�u{QIhNYU��א֛��*��;F�e���?��X��q~me���n�c.h���Id�
�ۛ��<���L���#�N"��3h�媤��2�?�6��+8�Y�&��Ί���`��N���{Q�U�Hd�Q�Y�?��%�zY�����g��2g��2�1�{mC��+>����(Ń����?��H�>��~!p	�O��q��+�&f�cMC.y��x���G�3>�������i$`-/&�Lp?I��{�ԡ���L�P��T(��n�:������c�$�EL��ׇ��h�u<�-��3�nYt�*9gt��H(Y�Qa��\s��*lF_�@��^t�x^EV�l���~ެ<�)��Y����!�r%^EX�f�K~M����lg;۟�����v����i���p�Zc����;AHz)���,J������&b�K���h��U/i�՗�D����*Zs� �����g.V9���gy3���K-@�aQ�~�)���8�*�%����6U*?�=��P��c&�0�������8��"���)�򋸘ANw�sX�(HW�o���l�	9Q4^�����B(��C��G��j@p���G��Ʉ ��2vH@�d�@H�����E`��t-:�c{�T���3,�� (
g�h��P;�l�"�`Y�َ��6����X����!��@�1�+БK��d���
Vm[�1�>昂 7�^�+����������n)S��Ȁ �����8���@rn3e�NX*�,�*���s�I��u���/�P<�8��ǶS�"�/�&4�5o1�
�X֎�0�χ u,����qBD��gF�*R ʪ��x�����+�S 0~/w�X���7NX����Q%�bٰ�R��,�t���j��w@5v5��ܶ*X����ؙ��O���bUǋ��e{p�??�g�d��gE(��w��^�M�;}F� �Sj�RK r��b���l��Pn\T�m~jn�p[�/C	�L�����&��Wj��������(�VK�ے�>E�p�J|؇\V�7����m������iy���n��F��k��xk�*��2,|�9 H�T�5L's�v�6W���d�C�}>Ք��<Gƃ�F9a�U�kc�ζe�� ��"��q�2���c���@n$6֮"�Nu���?������<7�G��$�B���D(��
�r	�z�u��	v}�i�a5�,�׭Ͼ��4;a"��~�ީ̌I#pzV���[�*����k�I	}�
4���m�~8�x�2B����!�M<se#?斌l�Ǉ�0]��H�xý�'��3�b�� ���e��$�h'���a��R�ľ.���~�_H)x�8��ٵ�y�=V��ÿj�*6��J�;فg��pO�"#�N��6��_���7�=��际��)��sS:{?���!c�Q��
+[��ېA�K��d��\e��d���'*3]��gd{������99�����v��rQ����o��0nR��d��%T$P��w��y$������-|��;���v���9�I���lg;��~�� n7y�\��?�:Uh�>2  8��ۛ��� �р�_��
T%�Ъ]6B�J�_0{�?�\gw]/]"+�n
f-��r�d�*��t��[^�n� ?��_.=���y7e��e�6$Zk�l�ڡe�|r���8h�� �g؟OCy�cXr��U����=�Qk���t�G5��/$H[��D�VW�����bA�ǲ�e��":�녨����9=�{'�:I�@�#�1X���a u�� 4ۯ ��/Ź�.0K%���c{�����j�����yǹ�i8m�����n���꟔9A���5� *@�@�(���8nY_�F�Q�؞E�����c`�M���܋Y	d��ǔ��>�
]�?�H��<KX��`,�,��U�j��  ��IDAT.�� ���v3+�4�%H�rAvX��<� o���Q9�}7J4�taʫ�Â�Y!tR�����V���@ꀊ+��mRl�s{��ʼ�Z�Jb��*��e���+��PB�U�J%����O�c����nW�!��lD�z	��6;!l[3X�sM���c%a����_� 4޻M��%uH-�Oq��ξ�����w�"M`�{�?����漗�u"��+�$̜Y��Pk�n>�}$ȼ�%�9T��N�`�Pr�4�u3N�5��㿾v`�໮"���B_�kW^���"a��ԩO���8��>";,f����>*_�c�Dv _��LS�hι�ë���S� ��8@��E !\���a��k��K����6k�Jؾ,�}ї��������f�����!1ꚨ�P��m�A�=�]��q�e���/�]�T�<�1w�}�Z�7C���=���? �]A�	���G=�Ǜ�^�|��b ޳=��d��&e�X$���d�_s�	
{(r����P$�Q�Id�۰�;iS�tg���t��Ǳ��VȂ�������p�����������g��ӵ�H,��d���_ ��^0�Dw������P~賙���y�]�[;&ZhYw�l[W��{�j����S�|���G '��k'@\����	z��ceV^q�x^����}~pV����HS��M��͎�&�xҐ��U���//RgY�6�5wQ�R��D��������֟3˔����-��lg;�����$@�v����l�L����8x9������������7���;�a/�xEf@m��x�K�ŲA ���@�
/�Dp9��`Uf����xI������7 8b܏������_� sp�}����@0��T��67����0{$�L	��9v����7H�t��-|�yC ���;��j�͒�Tx��� ����я���L����.7��x�����	A����\��A� �����]]��O���s�\2�0"B��r*�|�C���
Y�1SĪ	��!�*�=[e�8؟�[�$h�b�A��x's��:�7ig�6���
 +���D��������VQ^�>�[�~z{wX������s#����7�O���'��C�͓>qCk7��U��T�<7���I��������mgU�������0bm�l��D8G�/��ղ��1/��z�x
��(�i�OZ�\�����N����~�v  ����lE�>��n7�g_�e��ȯ�7�_�Pi8A��-�Q��|��n�:�:8�?���
�����u-�-�[���p����`��?�Jf�umϭ�� ��QU��{Q���o��"?�e�rLv���;X)2��c�v/]A@�I��+�m���X���{��������ۡ
�]��W���?�ˋ��ѧPO��`��9#�_d�jU������X��/�[*C���"�)�	�>��>���c���xoo��p=�f�&"��۱��?����^����M�4)x�O� IՁcE(=�YJk���ޏ��X�K��-|~|��߿���o�{�ӳG�]�����_,#��n�ۿ�m���0^�C�d�����c���z�#�,�Dǻ�bA�	�2s����YZ:���">اT�����4���d��U?n�� � X#�\D�~~$#���7����lK�:窳v��Ȕٲp��0vo}�b;��yd$���# Y��s��=$���#W������IwؘG�FB�m�1~��v��%���*�Uv��E���������m�b�{�y�Ė�/�?�/��4H�Ue0��e�v�\^T:��zD.
�ȼ��q�����6Y��
s[y��X�o �ME��]Z8N����ސ�F^����D�m��Wstￗ��L�%�+����}������q50��2���|W���1רr��}�W�F(�εj�Ϲ(RJ�aA�T�=�e��g���*؄�D���.�b�xI�J?&�E�<��z��'Y�B��z.���&\+|ޮ�����x���r{��~�(�'�W����qo�%��	��Щ}�xި��+����	,ѱ�Q��o�3�z����G��������	����3<���v���i�I���lg;��~��4	+_p"�i�[�h����=%���e0/JRa�2?ǋ��:�!?����RV���h��$+ ���z?���ߣ# pX?=��ie�BW���S!_�U@&H_k�/��j˪�}����W:h��x�-���A��*�G�{?�w��=��+++��W9Z�;�n��WDn������ڡG�9������v;r�4ޗ�[`�y�#5��y�G��?��17U�w�n�J�2�:j���8�'��Ľ��Z���I:�E<�V���-Vs�h�e�fu�&���k��T���Y yǙ�U'�:�U�!׼a�&���<�O�P��n&�w���,Ĺ��>gY5�$	R�$��)1�9P����p��ƣZL��Y��T�C6k�b���>^i���z���J���.�4{�l�_���\��� �A8�����1�;��CJ�jV<�	ѱzx�+4*�a3כn�d��ʠH���Dɣ�,p���BE ' -�\T��"�j'zZ�\�����_H(<5N������q�e��mԼ*�� A*�l�BAޞ/!u����(�j�vDb/�^�9ze��y�2B'��]����!ﶃ9o@�q�X^�ژ�s�ѓ~�X}>�Hb��)�ež��
J`u���Ǐ޷�V� Ɍ���r2c�v�3����Qt�a��-��+����Z�)�������uP�=Z_+}>�<ќ٭|�  	df� ��8^M���?�O��N���\i��,�x��ŀ�*$�� �d�6����vl%s#�2gh�g����V$@�3<�
wZ����=[p��e��6�/�u82t0���"�,���`��>��Q�4��,�����f��1Y��~��O�ՀF��:e��y]r;��)4p�e������VZ_���ߢ�{h���j
)�f��{�~�ܯ9���$Zs��8)��<bk��������|��������-�$s��EPep�x%�|x���s>��U͚L�d��3�U$J��{��*s{��e~W{�f�z�uY۸�S��.���Ş_H/�_���U]ﲺ���%U+6���J�~߂�U}\��[2IE���Xk��׿���K8���v�����I���lg;��~��v  #�$�nU���`�5��f�a }���X]�=��6��	U� Y; e@EЋ+&Qu[��T�B���6�����|�_[�@WeLYh�Oߑ� m�P-}7� wPҎ�r/��P����|_P�_�)2��X�ɞ��� ���LXY-�J�O���3���(����ȷ��������?l���X�'�0�S
^ܗd@������@�T�N�Q�^��S���_����߻6id�@�1۟�o�Ρ�=�Q(��.���F�UZ �>Y�j��-t ��uD?ϲ�+�����y�YO x2l���;����+lu��2[F�o1�|���@_�yI��T-�mg�?��A3�:��m��`��:�{7�o���
\%Z���y܋��	XtK'?'Y��߮��eWfTV�����A�{a�B	R� ����X><�͊�Q҃�	�-����C�n��V]�W>�D����;��jU�ɀE����� ��������V��5�>������{6�g,x���1N`�#DJr`�����g��h�^���ER(���1�����1*���xPm���1��*uI�,� �re@�قk@d���|�HK���G��(_7�i&���
@���ccǬו�,�k뤆�h�{ q�xX�e�����ܤ�H}�|[X׼<�d
���
�|S'����꺶���}�5�:�9��7�\r��w�����;�,=96q�) [����W�v����6B��_���WĮK^��g��Gj���gk��H	0Sƌ"<x� 	�3{�ߐ�uCǝ�c�#�����={G� �O_g�t}z��΁f^��Hq*����l?�"B ��ĕg��1�lO�[���?�Gh�9)$���K�K�����qN$�gl��oi$7��͑/�oC'������Ӵ��gsW?�8��hJ�Rǳ"l��f#Ac�S�
�fqs��	m�.�R�m��}���PU�bSRT{�g6N�!4��-��]̣"���k��^��yw<�22W��a��.T�ֲ�����Z��j<<���<ѹ_OH�u�hZ���܎�%8��j��X� �$e��{��[�������������x����lg���� 9���v���R��x9��@ #�_X�Ue�[��}��{�Z��54��e����xъ"@�� D)9�u�)q�
��6��ܫ�D�P���$���v)C�c���
7��-��#�
��+��dE�߾���Dxu�+�?�D�o���Oq�����:�Of�|�Ny�#���iY�W��� rߗ��vۧ�V#�#�/|�^v�$#'Н�f��ۭ�x,A��@)Gm�Dj� A�D��g[�0k��$���a�s����2'|Ζ�$�F^K0U��<��aM�J{�S��12��	$#���)��$
T�ץ�wҎ�rŃ���n1� ��@*�M��jJR�>�;�T�S~9"��}Qt���5ܘ����Y"a i�<�@ �&2#�u느�keh00&i;��o:�*𲔻����'����s��Hh�c��Z�%�m�:^�F$� SQwPu��̧p+*���	�9��� lSL}���D��;��R�x�Y�>�/��Ms��u>n�e�R���iWt�_Ѫ��8�jp����Ƕc�;��'"�H�$�v`͕�jT��wwS~0lw�}�g��/k���u���1�N��9{���'HXE�Lt��^Z_��eu�3�O����Fs��~���-]i�����_�L�a�ue]�,�k�ǻ�{�S�+`6.R ��g�,,���[$�� ��.^�����7[����߭���$)��u�͘�#Wkd|������u�+ʋ��j"�l�P�P�a��/� )c$����P_�Q��:� 8r2�����c�0�1�`Dƌ9h�YSWVҎǠcr{MW)uE��)XKni��#�b�\^����n�c�b��<퉠.�Jk��� MD���b��jOw�+ e_�u�� ��y �Z�_3y ����Ӝ��[䙃�N�h��[6�Aj�c���<D։�I��ױ}'��|��$#IR�r=�997��H����s'���M.d!1es���j��di<�/�O�5�g Y�ESq�p(���j�$��w}/�]F�?���ο��b�Wɰ��T3���������yR�o�=s�g�`�>G�M�n�K�'üZوq���n��5��x��c.X6�޳�DnE�߈g�k����~��7��۷o���>���v���Y�I���lg;��~����%p/�����/��.u���/���Qys�� ^n��Ѓ�d.7@
+� v��t�/;�[���;(�����.�{����*���R�0��ظY�Ҫ '+$&1Շ�lr_��f* lPP}@�!�,*����i�2M*Zp>�@:�H�k�1)Y��8���,8����{w''u�3z� �_�ix<�]�*�ϰB�+�u��.���j�Ѩ0D����s$+�����@�`!�dD��2�k_�>�RMԇ)f�X Q`�0C�5��Ge+l���܁C�寧s6@������
��E@���0���Q(�$�����:�@>̀Oe����꽚���<[%i�Eu�4͊󋄐ٖ���mQ�p����rn����X��ߔ9��P�XdQ��%l�Abv����	�l��^&P��
fU��>fn1%ņ��7���D��-�����m�x@�_��o�J�2@�m[:��<>@N���G 8@;nS�߫���N��Rzp�r̗5�f�dIb�P38���5���5���H�	��ݷ�z^��p\�̔Ap�6 �0AH3��s'���c�C��V�3N���sy�?�߰���9�d�UR'z�*��Eўg�vb����Z�.�6�q�"d(I|���t�.��by+��O���k��α����s��6
���.�\=�F2S��%�ܕ"C���p�{Vt��5w���9x�l�V��8�@n�kW8�%����^g���R�n'@ZI��@��*~(HD~�<�>�GJ꤈��s3�bŕ	�=�~
��Qc��^�F���P���&�r6��Q�:=;�y¬�8Ok���A�(�]�N��ve��U���vV32Ta~M�=��	��̎pU_M
.}w��+0���3+<o}�,MGq�<��2N��`���2�j45p$��������1���^�>^�[^Ԕ�������9�f[�����3I���1�e
�A����h�O_O���p�*r��Y15�:�ԋk�ue�zN����= ��\��|/����<�-�jx�=���I�ƽp�u���s? )�@�w�|c=��P�>�)�`A��1���o᯿}��?x�����[x��=��lg;�����$@�v����l�L�+�\�:����ͺ�e��v�G����T�����ցj��͠$����i_�*(���A��;�������?�%"�
���?�^���r%��R�B3�	ʆ��^xgUly�
R����R[�0��uXI��O5��lIf;�`� �/�	�
˫Eꇲ7~|�<~8��#ˮ��|f��>��T-�v)Z��G�2@�GR]^P�ǥ����pa��C`�� r�l�0�����l�Nd @\6K��XF��<����=+z$!��g@���*�`�3Pu��bY$�.Cڭ�1�������v������j��	FF� ���>��Had����]GD�g��VEn�C,r~���^�u ރ��[G�,�R�������UU݁a��� Тj|����{U����B�^J���ݚ$�)ū�E* \���8�";�n��f ��?m;�e�jE�)9�8�')���0d۷�x!o��ϑ�����rD�vɖb���� �R����K��9 ݫ��'=Cz�����]x�
y�/c4�-f�6�j'"���"�\j�k_�A~8���q�c���y�8�|�����`/�k�~�J��T8��4��ٟÂ�3C持�O10��E�:/� Z9�%���J�������9w����q����p3%2T`󆮻��F	7�Ϩ��&����=��xZ 4�W !X��m��7�d��48>��[34?�\	���|��ϕϱ�4����m&!���u�o��d��Y��Ք�N�T˧��A߯�)U�c�JN:�a'e�D'�x����m��q1d� ^���8�:4�H���DM�eP�N�̊���7�1ϱv��G�����~VO�kT�sܶ��ɴ���9Q;0�6U_��P����{Q��|��Jk�q�d*�:1M$�Z����m��_��2(��[�\�g������i�	�;)�c�8�q�2�I���>�����1W���ﹾ��(�MB8�o߾�9yC�O���s�}gV1�2n'��^z��[��8�rH_�ڠ�`�$c�UC������d9����m9Ox���<���XC����B;�g;�����n'r����lg�u��x1Z,�x����Z76�~����1�,l����i�PE�o"͗.��!1��,�e�� /`n�0�����m�����B5E�޺Oz�`�s��E������eFT�5��"E������,� y/G?&�ϝ���x����B��a <r>��$��p�4�����n��	&w4V����� �3�����b FP������	� ��7f�����>�Es
v
��8��r#�����C� �e��-:4�j�6�§vR?�P�����d<C�!���,)׋��������o�&tESq���\|CvA�`�8`�d���j��6:7'B�D�c.9YfU�)���w?@ڠX�==ϳ<��:l#%�o��L��"�耫�#�_��o}�U��W������OΣ���*��^��HCUBs�����nT�^���� ���I���*g��w� ���X�s����s�<�'R���T�6�@m�w�����Vqm�jC�hf�Uh5��i��R�0�h�Ҵ,����Ky-��}x :�W�C�X�N.�dP]�mZT=�,��j+Mj�9��-�D���xm�V�Xr-���!�3x�A��ð����_��~���B"ف�lkj���s���������4�"r? ��!��M�]1R.QWS,T�q� ��J�����N2z�4���-�x�p��+XO�}�B�U����$[J�+�E��f(��;��8+��U�I��͋�=��o]�U��?��H�A"�^0�|�h�~����~��(��0�l]��X����2�L4�8��ooo'�cqB`؆�U�(|��r.�K�ʏn���z
�E��?�|{�?V\?K݋C:�@�~t��Ϸ��D�vbԬ��u� �^T������+|�t�R��8��ů䇓N6`��[��m����w���>��4 ݥ^�y�S@�`���W2���i=�߭���Kj!'r1|��}��g�c7�Ij�8�
@aU��a�c�a)��~*ؽыsFa�޳@^�=�U@b{/�}��8��[������y�D�bjo_C���,jc���>�0�=�[���ͭ?���8���v��?�� 9���v������0P��`�E�ď�8^bd9������gA��MU�j�/>a����İ������p���\��ђ;�
�j>�c���el�/�h��X���E���uP�m1��T�GO��
_2�˲ �v� QS'@d�@������>YY�r 

�1++�r�f��c5��;<�ݬ���X�,�`���h�EpN����b ��{��Kv�L 1�����P�8R�K4T�*�VBG�Ĳ���,��d�u+Ə�(9��|��;蠁�r�oVt����E�72kv�o����s��S��=��Ȣ'"�IlN�JR/4�\	���0�YA�s5��&Z�͢�ꊱ��vuM�
PV�j�h���޷gX[�`�:z%ɪ�2L�.�P�(C�Uя���fά�7��׉4<��B�j��.��ٺ}���W��,H���o�F�~�ZF�
'���~�+�/k��oG�@(��3��R���D�E0/�~��-"���B��B`������7N�f#F���?����+T��:!��$�c���5�����Y�v���s��+\ȣ���Ǧ��u'D{Ye�����ϖ?"�E��z��l��J��<'pJ�d�
�cp� tb| �:���� �7M�����>USkQAx����<���D��a?�Ⱦr,��!�x=y}6�%�ƙ+�}������*/�ʨ5��ｿ#��{�f������ۺ�1���	�X�1GsW����f�/����~|`>h��X �V
ר�a�� ��r�"��%�;Th��=�D��-Â��zZ��MZ�Ǵm�q�����U#R���*��B��\sR�),:)G����Rj��X׾�uO���_����Ee�~��J��kaֺ�J�ǡ��J�J���q��N�)w���E���-}mёLم�^���i#(�j�g��$%�w�]Y7T<�Bi1�T��l�����C�{a��=&z$��1@����p�.]��}�E����cb���rl�m�a�:o�$��R��XR'��֕�}3N浞A���g�$�8�s�ڪ��T p;���<���r�WP�MI�y��,�yO�Zh�l�O>�]o�d L�����:�j�P�1Jڀ�<����*R�
��h���ɞ�9p�X�����k:mUa7��S*ˊ�8[@�:A��nq���z˜�s���SJ-}�w�;a���r<�ύ��>?>�r�5g�lg;�����l'r����lg�e�@2e3�	�㟟F������Ǐ�m��O��<aY����*� �2P���� H� ��?iS�������	��x��� A�˷����<^�3�&�}�-��<����?�V)��
�|Un��<^,���%/h����[؏�G �����Nۓ��Z����M>�$�V�A/��Fpƒ��@6^����dZvE���B>���G�jb ���G\�"�@E�;�����~G�:^�/� 9�'�`��􀲗s'*T�*�*�n��?Ɔ�^h����}Wh�z���sc�D��971���TgS�=(d���i�g%�s ��q.
�/v�9& �Hmp`/���
Չ��m
FG_���8`��w��b�}|�	��:6���?�r�����_8��>��OK�s��5r�`ҤR�Jd#;k�Ul��,�.R<�=�R<�v+4��,AA� ��q��s�������N���|DQ�ή�-��d(�A`��qW��6j1"�սV������~V��XץWFǨ�sWc\.�}�Z@p4)ӧ0�$�l����8^xg;ZgY��N��D�= _�!�u�� ��+;F��8�o�ޭ�T����#�P�e[��^LV{H��z�����On���>�����y"���0��Wf���[�����Dbe��QY`-�sVj����CɃ�" SAb U2RD�����\�gq~�V�sJ�G�c��#�!__7�j�������o'H�5v�6� O0V�dc����+��`��1�Y��^ޮfÇ�{W��	���p�r$0�k��'�M�*�@AI��RU�܎�3)R�?t5�GU���n�2;�9~����#|�����۱N�8.����1G|,@���-�����+���%����\<��*Cd�U�m9�2���,�h$W`���s6�F����[k��c�N:�?��<Ƅ"�V�>�c�?��Be�Ȅ�E0��{��v���c��!���К	 =���� �6dA���c�k���|�5��dᜬ��l��"���i�8i-�̬@(zN�=��sV�]1P�J���<�����8E_'%C��W��s�^$2�$}_6K��n��DTtֽ�/����|�p�>YXX��
nC�7%��r�XP9�"�gVs�zk����)���(�b�#�ඥ=�m����ׯb*�a���2��AW YnG��*v�/Y��d���:���)�'���|���J�qT�aYYHj�8�QyoްTHuR\C�y���='"����Fc�v�ix�D��Rۉ�Y����q/�uW��
W�M���V�q�~˴:�����`�����zܳ�ߎc_9�$��sxs��?�Ϩ(�"��<6W})����yW9�&�����쏵�/�x��������?~����/�lg;�����o'r����lg�e� tQe[��9Xl��r�V���%	��,\�	$�:�_�A%��B՗|�o�5X��7�b�y�%@1?^� �?�\ Pў��Xw�;*{*D��������/�"S2�:*?��}0P�62�^��1�V�QQ���vU�M��V=����x�nˋ_<���\ә�2_�ԭ�߽���r��������7���a����)l�u��޷���&�|�'�侻�dT��0�>	
�T�}��:<����@R����gy��^��b ��+[�/��ݤDhY@��������w�K� �~��!.VfG_x��{��PtR�����~��﬎�R��n
/�|�͔��l�vd]?���<�,�g	���$�+�A򜏛*��ǹ����^��jm]��9�`ޏW�WSZ$�Z&��i��R��l��s*b�VT�ԝ
�^%^zU<�%8�e5X�1�L!�60���^�`���n��uu�H]K |=�ȁE�	>��X�"��m{�z$�>�G�8��}��sn���K_�\!�F.��C���>e.������C�5���pk@˳1�k�y����>c=nP:��}dYt+���L�:����>�C�7:�h9�N�vxm��)�<%#�F൬�H0����+/
���۵�h��]\�$�/e"��;�R l��s��g"�������~���@�l�kߺ*��G�r\\�ʨ�kp1�;�����q��s�#X�� ��6k�;A�c�'$��u����]�z�$;>(;�?b�Bɔ��A���Yp9	I��//>'7�TC������euP_׹l�p>����jcR���P+4�W���^2����>�W�����j��
fc�k��F���ίT�ؤIe�N��rY�t���3l���v��[m�$���|7�������X͒*Fe?�r�J&�=�kK$�$~��%O�e0VE�_x=f|`�m��(�j�J�FPL���bV�"���j5���w)^���� "�Z�~}+��,�8�f��E��]��d���CZ�-�LdY_hRoV����g����y������q,G��"�̪�ٳ���s��Ҏ��
����3{�oN�;�v|胢(	� ���+��ԇ�d�,��r������믿�?$^���8Mq��%�	;W6�\Kq���䅖�P����??"���g��ծv�����E�\�jW���~�FuDC�����j  �q� �@�͞sD$������Jp~cu\<�c� � t$�A�Ϋ���	�/V��|����jQ����;����:ֵ��I� �`g�_�H� ۀ,b�3
�U�C	���1��f��.�w��7Z�l��^�z�������`��<�23	��~J�Y��,��+P~x߉��Y1�����:�_�O	�%y�V�E
��kGV���#x��G��]�S�����R���k�l��,x�뜻u��
J�,(���
I뿔��Ӷ������c@�W��~Q��Um
 U*Y����AKV��6y1M�q��b�`d����дo��`e�D�}��}C��6������ -V"����8���@���Ŭ�#PX`i2�)U{U�'zM��|�M��ط���!��#��z��r���4�60�M�஫;*J��m�t�&�%�­2����!d��Vx,�(�s����Pi��[���~KpGs[�lv>�W�0��1n$�/��Z"S�}|�eژA�}����[W�$S�`��J6%R�����l ��ϐ$�e�Dr�2��gŏ��Z�k/������B���=+a2�Wn;A�6\ٲ�@��ch}���<�w���lyP���0Ɠ�h�X3��{\�<Z��Ze�""��[�P`2.\~��>�g���W��!H����X�~��.�
��9�}刺A�M����3��g��U>Q�m����DV�C!���?�F�eS�MɃӛ��x@#њO�4Q�C5���W�mZ��6���f�&��	�)�����,ʰ�t�͏�O���{��������W�%Y=�<���|:>ٔ�6r��᪔T|�c��
S_��R��\���K���.>^���S����A��ªq,�iyfuՌ���O��گ��ҽl�X��B(	=�Z�IϖS֍���yj��z�YR2��d)�-�kqE	H�dۏ�K�b�����8o���$�4��zs2�1�h����~`�P���E(��j���ާ���*,\?W��C���g�$��Y�b�a��쥪�� N�lze�ұ_��׼���C�!��S^�ծv��]���.�jW��ծ�۶��R5mf����#��j^��J~lD5�j@���������d59i�pQdj7�e�)S��(�	 �%�tk��nʁx��G|mRi0��N����J/ۇ^�H�8>��������i �=\</&�J��Z�SZ�f�i@��<����Nz� I��Z��m��W?��ρ�蛔̒�$k�%+����J�0�.�t/8���(H��1C3�c?��͗8vk;W&3�"9�������T�-PmL�*���J�5�N�6S] � 9�j& vu�f�����W����A���oR |��n��C��#-��dA�$Tn�����-���V�?B̱Z�q�`�|��I�b9�d[������T�MO��T
�x�gi@�"���A�b�J�-Q֗��9�sr{#rG���ܠϧa?Uu/e��U�)��w)D��1ɯ\*��	�����@�����i�"�{2�0�"k�l�RʭȦT���*���ey�+V�I��	us�u��8�&2
���8�_/@�-c���k�� Wm\�b�
��3���!ZWQ��I��R��Z�� �R�2�\���4Bβnq U����[����/P����i���ɔ9"7'�E;�������["���,N��:��S��Rp�A��IVO33I�V��Pj��s����8��;� �}l��@)�ZXa�._ oU�����`=U�w0�ہ9�ʍ >�}S��E�N�pmn���iYN��c�X��"���ڌsϲ.���ds���b�A(zߒe�xp�,���C���Ua�Mf��a�K��c�1�	NO����q��z�^��rU\�Bֽ_?4g���Hb�ޏׯ�~M�N"�_�-^��0"���4�s��)���uT����r'/��8������n;�bY��A'���BX/�A$e���x8GG�M
��+��h$�N�H��B�8�η���vW�NM��r�t�䖇���.��I�~t%�?m[."�`�Z8��4$5�oc�;$V&��c�č�Mp����~i
�i��l���Ŕ|���5�6z��)��>��ɚ)�����g$�f^gJQ���2��e�c!�B�s�OݒUET��fؔ���G���%ex�s?��G��ծv�����E�\�jW���~��Z�Jm��8�Tx2*��H�%��������>��/�@�j���|�
~{`�g�ߨʠ��]���~�� �A��V2��m��(��\f���ɪ��{=��n���w��Yn3�ڙWb�9�t,���|e��L���J<��*;&'��5�6�j?6>D�C�m]�A{���@:[ą��s���G_=�u���>���o�$Q�a{���O9��<�K5�� L�B�*P�|�{i�g˟(���]��ظϯ��m��W���� �uϡ���oy$'H��y  6����ϰ� ����%�֩Jt'�V̞�6@�U�k��L��
˼wP'��__ 7�n��K���u%U�S5c6/�o����q��2���"�9�d�5�Rt���?e��Y�[q���=�}-�A��/�s��O@����_�CHx�]�夀ۈe?I�HW�&�M1�ۍ,'K�S�U���R]i�:a�${*Qm�e����d�o�n�͓��^�:������]�/n��L��u��C��O}Lt�5�yN��T��]��J�*K7&	H�s�+g<����a������dH1,�b��lպm��������=(٪�S	�P��*�,���$��UeYD	�BБ����5�r\�>�N��Q�굕
�Ɥ��vs~<���}����dY�̉7�px�&+�i��b~Õ@�Xe��nQ�#�`�s�l��)>�&�y�y"!�5�W�;�>���1{+7�K2�Ne��a���}UH�-�0f�9�m>T�C�gl$T:��In��N���\t%�W�+�������kcV�w[���I���)g!��R�3��,�4Z2�cf��T�?~�㳭�x�F�d<�]����+a�I��m���J����9#]!�}R��t*V n�o$�����}#1��
��bw+�xiN�O?�M}7�78?6��/�b��o��8�����X�2�|=@ޯC9��mܒۀjT"�����y��̇�Aͮ�|�m�\����%�1�^l�+��,jP����X�Q-���s�����I	����(H�FTP}<�PC�j99�X^�gz�ߵo�E�m@N�X�PE�� c*s=��}�9�9#s�q?���D����{���]EX�ֿ�������>���������]�jW��߯]�ծv��]�k��N���O�������"=�7�1I�.�2���l�X�! ix�aY��[,�?l�}��b}5������H���S�[h9!� �H=@:@�[�<���i�4	|����� 顢x2k����O�ռ�Ia���{�^ۋ`�+�4����R >Ͼ�
���[ ��i��pp�B�y��Տ�3�@��6��n�y�2�2�~S���HyUe��_�� ��79�;AR��A�+	�Y��H!����*�@g ��ސ���jH��IFԔ9�4���T��X�� Wx1�$v4����M���@^�<��1���7�����|%��y
���������m��x	�T��u{ P�T]�Pzn���f��9���MI�4'Ϛp������J�y�*%�Y�X�b_d�f��+����@b������پ�> �ª�Y`������y��!�\�yJnO�-�p{`�f�.�+M�٬����
&��� ��M� 5N�����\E�zyI0�L50V��V���a�����<,�l��R�!�#��RXs� R�ApM��؁�9UR}R���2�#R��g�&�A4f�U[�w�F���ݎ����X���=�qR�xu��F$�G?�EF.'`�{�}�����fS?�x�οQ,��ǹ�M��,�˵`���VU��ɫW����9����8��m|T��_Dt8��|�����}��\n']v���Ӟ�#�7@�m�yE6I��L}�SM����s_tME!@�~� uy��s�зs2U�VT��b�J9�K,�ǍrZv��"f�/�A����=[Y}������ۗ�Ί�_YR9�q���#�JM�ZK���9H.R��6�+��e��>�C�����*��޶�F!���M��㚌D�1$�L��D����"�Z��qLe�Q���ny�e�I0�T��:�N,a^!����D�P���;�2*���`t�����˄Ƣ��{ܫlCq�w:dZN,L[([����hh�G��0���l�x�&��VV�`��c��^�=Y��q�0��T�Z�SS�%�ލ*(��F�{K��{��~�3���'����{CD�ծv��]�o�.�jW��ծ��4zC��<��@���x������@so��G0���n�b�g����ڀX;^�̊ �}_G�̰�ɲB^�L�^RJ �A%��u�CP8֗L��I9��%�u<_a�%��n��vӛ�Mp�u�X�]=��N�ܧ�}n��?=��6�/C�����6#z���s�R���T�[�4��FA�R�息��Fy��&I�>�'�\l�a���1V�:�EJ��Ҍ\s5�ƇE
�!��A����jW���[����T핞�A�υp��UOe��Vi ���8���٢�������lC`�T{5z,����\d�d�[�k�TJU>l�)�:�����y�7Q��O�.� ����շ�?�4��P����R3*��ȁ�BL��$L'_�Y7��D�U|���1�YꌰY"�  �6*�gT5��Pt���:v�w)]� �)�C��#ΑnsC�ٛLͩ�)�1��U
IO����0���[9����^%�=�����l���������dƠ076�}�3�6(P5@�`$�l�T1��~�8�N.s,��Fp��S�n�2���9� �AU���O�='@<�a]Z(.0F�Q���<#���&�\�m�q�1�� �)��	"�g�<���[�����|,��L��P�N{�S*�,�V�2E@��/�7���+��v  ���Ǽ�NNfV�/�Pnu��f��}��s"R��K}�F���1��LQ-ϯ�ڤpp�B�we��V̛F渺el�@�e	�
���6�̪<�ݝ+dI�L�}��	�[��#��1�4ޥ�;��?�Y:��':������q�`2�k��1���',�}��� tW�h��r���A]fו^`��"�$�ʫ�hn�և���d2�`�b�p�8��#��sn���瀏�)��s&��������G�Xv�;��O�-���/��:o�J�=�	�u�<C�G@�F~���͓)��_������Z��B�=���4����s
|L�8[.6�"��(�������A����ۛHS2O��r�WN(/YH�
3=�mx+v��c�����Id����~��/ΟP��������ծv����or��]�jW���;�h|ؙf�ݦC���V:m�i�%��h��e���������c��8�-��]	��
V 
���	$�A,7#?*�F	t�*�$�'�`�H�ؗ,�+�v﷛T���S8��?�����-������SA���o!��1x�H��*>�Cs���T�(�+�$8�nH����a�vP�}�h���{)Ȋ�ºalͭ�|#s'A��UV�.H��0� ����l��[_yJ#�ā �� �@�血M%��e-9G��@�����v�Xw u�d�� tT�z=(mЊ�ӝ X�F�؊}|<b�`�6��	� � �[�h�@�q�|��3hN�]����S�Pʍ�����qf�:u�D���6���v��Pհ@j)d�����2>��с��K`M6��.͋����3���P��8���I���敦�F#0���Ƣ�}O89)�J� .,$\���)l/���m��UWS�D�,R�tB^,�G 2�ue_��/�=*��j���f����]n_v��$��@>M����O�Nz� r�Ī�����Vi��'���faڝDr��T���j~̱�c�7~b�ެ�~������l�e�$#��E*Q�b(��`PN	�����\���t4T�ok���[�����mb.��\ђ�sa@���ge��_�g�ى�l����}u`�[*a��b3%�����/�W���{����(���f!�1T�Q�}���-��[B5�^�6[����rkS����/x�L�R���6�x���t�@��ڎ���>�
||>t�m�@Q	���\��;��^nѧ�u�z�d���9�g���E99�U99�t�DGX4Y*W�l��T"�z~��a�e��"z��ԭÜd(\_3+�fa�\o���۝}l�d��z$S�Կ�ĵi\�q�~��8Yf9SS�_'�pY̦�٘E��j���x{���Ѻ*�5�q$2�)��1�W���Y�G|�'p�v�L���
ߚq=�2m&S-������x/lJ:;N��T.����(td��撽8NV�z]�T�T_��s�ĝ)py�%]��n�i�M�I�b��L��1��Y-P�ڐ��Z�
�DH3���U�J���%4��כ��{�G�t7������v��]�j�v W��ծv�ߪU��6�������2��U=[�c�L����c�; b��Okz�"D ���։�cQ�����~�x>� >z���U�H�����S�,��-�R��*��4SzlIʓll,2�A��F@`3�1t���-��fVn�E�,ScDu].���r;�`)"HZ��g�9�a����m��ܩ��H�O�`L�b�vV���{�ф}X��~ 싩D�n�l	�폿>�G�/��U2$�&�Ri8��lD	2`VZ�s��}#O3�h˜قK9���@nep���E��� p�/G_�M�=@��)S���;��J+0a��lʤ����3$ ��ê���3,��������WZ�(/�P(�xZϯcC��{��훀���kk>� OA�Q��JY���c�c|>�#��oi�c�9�0h d\��\��G ��Q��:�* ��� `�>�G'��"_�W�l$>��[�$��[�N=)�Nl���mU5t�J�ms��Y02r@�� �O��yX��I�aӶ��s�v9��������g�dr��G���jd�U���! �{���yѳ1���N� �)��u�M�aۻ�cOPw���d���1��N�)k���Y����:�c�G:^��Yw�����H��k���=�� #Q%�����Y����������=�ܛ#Ӿ�9�r���/$�D�g���w�G�g�9����G��fGj����:B~1O@��j'�{^�l�L���n$H$���>��({9���#���vj�V#�gζ��U�7l��٤4Ә��x&�`E6sǼ���ɠo�wW}���=B�IF>�Z���Pm-T]ߌ�v���(����_�H����R(�$h9��c�4�����>�y!
`V8��(5�a� �p�����Ī�_�	ޭ���][��s���8�`�����g@ya�Sǀx�$��*S� C��>W�b�ǐ��!��Lp���o�m���
�� h�e:!QMa�<��l=��`��њ*�j��K�߸0g�#sRFے<H��}�c��(B�ٳ���8��A$�#J2;́\�w�ŏ�����þ϶���z���7������
��2[�L�{>�b{zF�Y���mN.�+������qo��2o��rYcR�"�c�jJ�d�hY���d��Z�*j��c=����dN����IPV�J:�=�q?U���������2.S�|g�E)'����cnُ{��,�֔n��M�>ݟ^�jW����.�"@�v��]�j�U��&����hV��i=�r�)4z�/{��VUvV���Tn����*L{�?>�n���������nf��#���j<��ZOC&y4)%�i���D���"�� ��`�
����V�D��`۾<��c�=Q��L����>����7��{�Ghg��j��~�j9��M��������ї*�˖S�Zy��z�D�K4,/��Z�}��=iK��mt��1"bk�g�LE��G�����1n�Aރ���=*?���3�����i��a�+���ZsX�p�l��Pzep<�u�H6���-��S��n��}(�������s <��bqL� ��=��������|ɾ?�P`�����u��#��T��59Ʀ��X�8�,�l�l��%T� ~m8О�4��{y��8%������K9�]�nUs����`�T S�jw���N2���|Ӷ�Y7w�*�^=��ǈ&��x6�T6F��<2/ٲ
,\���<���k���Ѷn�ݽ�I!�������-w8�a�d��̗qE��N�4{8l������ܗ�|�,#%���06��N����.���k�Bϵ���g�WZ��4�I#��@�md^\M`�j��:��܃ۡ��u��j
����7YrE�7��٬�V7��b����;ᘯ�Y������['�[5�S�I�xHQ����XaM� s���mq��>?�EU��H��t"S4�8H?�qث��:���>�G���1�R�߾=� :�uQ^���,꠴S?<AP��:��'졲�����`��a�{_z�H�f( ,����Ӯ�?�G�*ߏ����y�S���TZ:�f��D�"�׼�~F&�)o�����@�|�!���Eq$Xv#�dm��)҆}�L�w��$�\1X�D׾��۠���$~�H��ag;=����wg���C���sKH�i�9��<��`\��"`��Љ�������8;㖡'�=�,�T��Qq�%ܺl&���B�1H�b��B�a����{���������	1�����ؿ�z�tmE����i����ۚ�⪳�ƛT���!a?���k��{<�eR)n��ٹ�ծv����or��]�jW�m�[��*���bU����
ν��Z���C��Q48�y�W�Bu��:��z" ���MF>Ȟ�mT]a����<!`�/[՚���uf��U����\��$�y
!{�~y��5�����;��3�U���ޥ>Pd�*����@�`O5v@�+ԃ��+�͝�N�4���Z�9G�;�\�x�G�cȷ�r3���QXHU���H��[e��j��,<��Ve�Y7�鸥$Y]͊�%�A�J�VY|;��܏���H~`�H�	@ l��@��*X��U���z����y��	�!��E栂��W�'�����\���Q.X�	 T��c��~â���2*�~�Q���*�u<�Y�X�P 
�\)>T�`��ZJ��yy�
� �q��a�4{+M�qWo��� w�$�Ϝ �O�6���e�*d|v65O10Ϋ��K�
m؎v��h76�ml�+ آ����s��l�|_P�̪ڵ+ �O<Y�6�i����e �CJ���n/��O��������ұ>W;���� �wu�HG���=28 ��S,C�L���*���`屟�Iab
�U�!K��i{r%��6*�v����0��0�ʈB��v��k��Kq��n�'��x��q,^��>�b��U�+g��~�/FPx4,wS
���N���1���o<ղ�4�
�M�ע1� ��c6����(YhiȬ$S�����~���Y~mru���y�9{�K-ȼ%'��Sշ�|��*Km��q�!�~�l8X�u�:>�s�����L(tfSV(�Ɏ��s�d6��#<����P�B�� �e(_@���v��2��R�ԭǔס+��[RN}�P���c���_���e�.~nD��G5�o��5$�����~ ����Me�9�s̵��f�OT?���!�{��n̩���9�u��y�W�1�2��=�˅�ϘZ��י�2��y�+?^w���Z��/|Qx�u��w�j�}d$����9��.�9�YA����={�3�0�sϡ����]�j��=��L۱)?�g�u�y���):lgx]�l<n�Y?b�o�[Z_�,*6� #�f:��*�	�,T��z�������|��d�z���5�w��]�jW�{�� ��ծv���֍կfwA¤XYi������¦�=�Þg��b����~�NO����"˕�V�{��F��W��s����5:'Ѓ��6�~^yK�g���7Z�P��߫�V��/'l��	�@��3�=wc��w�����l�\��m�m6�ֆ�/��[�@�r��V��;
���;��.����r����6 �c�8^��~�%ׄP�_��A9P� �Ed��@�n�����ڌ����B����-�nX���{�-
�PsIX��[3��ʲ܎2��[w������K���LtȗjA�Nf8X;�\&�r�u ��w���P������I`�۟�b|m��2s7����u��1|i�"%lgt�0��9:��F��l���~���;�=y)2B��Anc5#.{Eq�n��5Su̦ P6�25樶u�4�4���8W�_A�0#'�t0�k5���SR���S�@)DvםT�ky2��-wvد\�f���aڷz"X<ˤ�^uL�@ �]��� |VB���J_pe���" ���[ا�6�Y�X�r�"-h�rˡ��=��!����Jb��nD�I��<�k�(����"�'#7�<�)>���}�}�1�f��M�Z��rSr�� �����2 yt�|�F�ZҏI){qiFO���
b[y# �[��H�k:tm�L�TL��#�";��jp|�p�\��FU�*�������66G0�5:VfCg6U>׌��H�-�%U���}�"�y6�>������=F�h�k,t3��B�\���`I�Wm ���E�r+ �ԭ5ǡ�F%��_s':���>�=�~�}~�B�qn��I")�!wFj���������~��ye�
�s	�6#��JM�T6���P_i����SW`��r��+%2(�9`��C�~������(���.cs�Ԙ��'�tS��s�� �F�I)s����Q��6�q�x��/C^XAR�C��d7��e��և]܌�L��`���C���J�7.o,��%�|�i:���b�C�p���v����۪��$�J{>�0�sq�~�+)��q�6���dحDP."�� )B��-_�jW����&�"@�v��]�j�]#ؐR�4��D�e|�f��W�D7e�����4u�~ K�C�5��Aψ�5��a�|�Ci�䊒�H���ʱ�������/f��� nA^�Js������:��֌q��?�(c_L˒ ��)^�וUۖ�n��*�#�p���l{����d@� �jiT4���QJ�D��T��Lȸ�N{�f���O�#��Y}�"�d� �O�����^a-k�[�Q��$.��q��J��x8��+�g��vK)vϾ��{Eq`蕪|6JS3��8�ȝ1$
�9��0ϪVWXR5��~��]����P�*��W�X�|W��������庪�	�#�Ɯê�[� �����<��g���u�'Y��Lb8�8@�@�yq,:h�`�sP5�o����5,�����f1�[_�D�G�7"F�9�7� T[�D����lY2u���93"�\=2iE�] ��Е�!`ֳ/<V��k�f"w�h�j�;��&��T��W�[��PM���c);0�'1r�f��jޖ�O6  f'���l}g��I�짲�oy�h�'d���R���@Y��`�h��@���S ��Ґ}���3�=�C};K�a�1��Yn�֤�1b'ӒG�i8�a���f�O��\���u�eV�5�'^s\���U��OqvS�|=�xVy��^f�LS����5�'�{M��7{� 36�������ɏ��s��'z�	L�Yf�w����N�Uu��YQAri�U�yɡ��sr���J���1D�Aָii�D3�*ט<��f�A�����C!��2�m�\�2�_����?e����{lk�TR9�$+�:��N�ױ�v�K,W׉xete*9�\z��[��ڕw��fs�[D�CRDnmQ���M$kW�x�:���Xޗ�I�.!%�w����jc.M'��ͯ�=8��}<��#Z��*9u��}���t������Ͳ����7#��yS�Z��jY�4+v�Xx�[Qa�1?,ǽ�'����ܷ�{�?�^�֗����a�B�:`�11�C���)/���Q��L$���f�����yNF��~��W��ծv��o���]�jW��o֬:�|�x�! }��
�S>>_?�+���ٮ�U.ST�z�C3�� ?��AUEz<|p�����z��G���rxVL� ?N�[P:+�6>$��I��H�j#�����aY= s$?���������9B#�c��6,����ۉ��뭜	�a�v+$��a���r��Z�����í+E�~ۥ1�U��T\�Yky�*8w��<�����m�t���A��C6 �a��R�7�4>��
�7�K1EL5�V5������I0�@��� ^�~�5���M ���B2�:B*�l���E��W���U��U����V��2FR(@��Y�������ߺ�8�����e�=�kP�Оg�_�D�$�@d,'}@� �uȽ2ߛ+&<k�<�v���w�i���4������g�s�(��f�.���� 1};ܮ�A������!^e�1����-n��H
h��:��y�6v{Zc��l9����n̉��B� ������VX��̙�����bj��`�zU�x�Ұ�d��>����ܽ�����@�縌�#$�L����Z����k�y�?��7�.���8�a^p���1(����?M�ӽ襈�%��]����f��K!����t�f����0���y8{���)�`o�EY; T�F��?�s��8��N߻�j�g>I�vL��;�����cH�N�>jP�x.�����h�88�fȔc�>f� J)ƃ*�5O�{�/U��"p��KĂ�a���_�:�8��V��i*"��4��C�J����=G�+�4oLm��w�	�-��\��u�b�|���_F�Ny���=E��\�/���v�y�ɚLR���Ȧ��=��\���S'R�8�V-@�E �6dgٞc;@�Z���I�&���������p,�)�=�_�wc"p{?�����s�*���W�x�����O/��Я���Wm}�qS�W����m�3�M�m�la�O�J����������{�IU�ֶ�D�̙�Zg�1����m���"?�vhE��VT�vtX�B;+��˚�x��c̅�eb}�
��Z��߿_�jW����w�� ��ծv���6��?w�����χ,$&���)�<���m��`�QT_�Էnk��dm"VbL��U� h�N/xT���h�%Ya�x;�~z�+?=@ydwJxnT}�w4Kzћ�H�x��@~l݃���'E��2���o �#O/�2-Rxp�cU@�=ȷUx[�b�mQ�|`��!�,w˨�*%%��Vr�	#�ͪ�����(/ 
�����c"�)��;)S�|[�ZM�桒 HS�4��c���g�� O���6�Y�=���,�ù:�٠��ҭ�t��EX�ý��Ɏ������n� v�+^�bf1�U�n���l��q0 �|�$@�x �[L��?�J���!��Y)�9���mc�XӘg���q��J�ԟS>��]n�>�U�
��s����w�-@!�9�y'fյm5��+9�,`��lZ���-�j���U�)�.h�c�ޭ]J�c��yH)y��Y�LFڈ0PE�1�f-�m�❓g�p]��sJ����fǻF�:�$Oa���i34��VA>�{�Gk�jǨ��>�3UF��Ρ��:���i�7�+�*c2�O�@Kc0��x�����C��ɔ�ӲU'*��^:�{"�m3��h�� ���A�o^j!�3�b����Ʊ5u�o_�C������~,�r�덪�<�Տ,�ߓ��p��o���	M�v�U��y��oy!Ө��@���ܢ�N�Mc&Eݾ����`u�����ɬ�4v���*���9��*�w\� N>-$e�`?p��(:�������P�����Q���wS�lF�n���FK%S������"u+���iY#���;��=����-�Rk�J}^o��OR8���׭�9��<d�{��Y�����q"�ۻ�1ϲ~�{ ��nF���F����l�1�W�v\�Y�=�}��l�0/�~"�$���	�PלI<͉��~ˉұ}pvB�_�]�ۜwxn{5�;Y��d�dMWWj����}d5�*.���
V���W�眠�g�.m3-��}T
1��M)}��MR��1^y�2�)�oִ�l���w����r�(>Uw�ש�`�@�q7K�( ���]�jW��߰]�ծv��]�k����
�i���, �ҺB�(�a�Ù��w�_F|��K�	��ۊ��yy?�k�S0��n9<���z����S���o'� ~���!hP�)����K���#��rݰ���B� �{o�K���'��w�mS�dJ�����Hp�䏭R��6�� ����Yu`�0vۢ�L��U�UHZ��1�8$��>7�~�Px �}|�z'
X4F�L���C:}���Y|آs����ll��G� �D���n�.9�eAU���� �5�*E�" ��*'��H��H0���EV���X���{rk�;����Tmd
*\�2��<��E�r��v��ӚO�ȵXn������e�'YC�Ma�D
���w���� !�Y a10L���@��_�f��
���W��"A9�[��������,��Vcª���<�j��n)4�]��AK ?�{�)U�o���v�߹-P���l5*�LU�5rV����-s��1d��
�^��!�D�04>���d6�	�N(�����+!Ү�#���R�q�m���F1K=�ט%�<�$Z�Pw$�r�٥!7!��X
��U(_T� Ժߥ�20�*���T��X�r:� 3I��=$5lk�b6F����q&9>�U���ɖ�ծ�1�L�/kTs� �,�6U��Ra��8~��8�����*��=���Ϊx���9o
T_����OX�����?���:��Bٍ4�y�܌�u�Y��ʚ�7�⠠��F��f��*&ΏF-ia撓�����"����f�����-}�9:�[��
B�fUwk,�J��J�8�W�{�/?���L�;W)�}�b�m3K��g�x-T#~�e��ϔ��� q�J}�� ���^��:X>�qx��ZC�6��
0\�V\!׏eo�N���n��GX<�f���?7nۨ����X�9*O)��2�}�CE(�Y1]D���χ�f^��|��m�8w;�iꖂ��Hl�<s�\�.K�����ITV���s��t���Yg��׬���MZ2EG��g���7�?c��A\�i�f^�{���y���̈#?z�[���"�j���q�����X�B�G�^Ff)t�YX����zk��?)~SX㽞6 �z4x$���wpn`J���X+����-˿��N�}!�v��]�j�v W��ծv�ߧ��z��B���Gz�n�� Ћ�inӖ^���g9�BLc6���U��".^�ؔ�`��.��s{F�s��\�o]lb��++��h�B���U�.yh��򭤷���5#g�N)����&֫B�WT�X!�$�G���(*s�������mi�?�]pp6H�T" NŇ&�c7�Yf)�<��6���a��~�*�����y��/퓸	)3��`�2�>���9>�Jm����b�a`���O� �����W��u5U���h�p��|p�Z<�����,��I2A:�L��� dx{��<���H�b`��[p��{���#սߪA2[Ų*�w�h'a[��iD	,��)M�[��t1�md�<Y�ix�/�2Y!�R��</�Hڪ�m���!ݍ*�
�����&Vp�V�~�|�����'������26�Q�"�46�t���R��[�����\�2���&���+l��XRd^<�����޹ll@`xy&���	Y�=�M�����X�-U�j`�T&���jζ���JǦE�����b���B��<���~�u�_�ohWr`�rJ4�q���1�V��Ͳ(�XY��mT%kJ-��bcLX�&��z�1���;�'H�� ��4W�$�zr0X�t>����W��Z�6�Y����'�>�x��������mR輇=+����c�q����%Rd�uՎ�AXf��}�ɺ>H<8.�&��y���1p��^+�O�qX=8z&Q��y0v�HAP8/�;?>����w�R�LKw���X��;��5_f?��zm���
aƳ���������/�/2�ȫ��,�٬�\I�'W�`��
����?LuS�s���c�9�fM�L����G��>�x�O\�bX��]y�&U�r鸒���͑�C��`��5Q�KX��1}>6f� _�W��'��[��J������]�Yͣ�m�*秧x�kP�	�z�׺�([�J�y�D�+�\ɡ��dcj�ՉDaΖ��Z�e�n^��*�;��D�kj�_"^��[����%��wf��c�M�0*���'b���'�$�寏Fz������֣?طfmj��fR/.uI?���9��'�If�==>�$R���e�	u0V[L��q2����e��a9u94�����D<HfV�x���;�Q#��]�s�p>��?���ZM�Z��us�n6�ȵ��x/h�68��s�*,��>#I�����v;��E7����I��n�A�ܠ���q�cN�Ђ�)��q�^�÷�|�Y�ϷTU�t��w@ B���cM]]-���x�C�Z3E����*<B6�1	Q���-]�jW������"@�v��]�j�u���,�U�&��I�$RU�=g�(�ؿ@d(*�_�x>_U>�q�\��FP �"2��:U	���a{�:��0|���U��[躾:�k ?�}t�,��x���m��e��KD������x�$�f���Q��iݷx�ϽBݷ1%4V�ߌ�t#&�}WH8�s3�É��m�6 R�o3k%��U��F+=�=� ��f[V=�O\��+�s�B�'y(��{��2P���Pw�FVRx(]`%�[�~0O�t1�� � q,tݬ�~oH���D�ڜN�  C�g��OQ�Y����+|���++�a�b��^�n4V�V�+TU�C��^�}R�|u��5��v��Xu��,�fS,x�oST� �zU6���+��-[��Z�1��a���� >�o�� ���d��@V��:Cu �{euN6�M��Q��t�"h]H`�L���d�7������q |,p��a m�ܧ��nA�VY<����j�@b�f�41�囎�ծ�J��1o��fK&[�^��^�}D�Â��e0Y��Ψ~��R�e�)8gK�8q�:��cS��n����KV�MkaY���� ��i:ק����O��������s� A#H��y3>�l�w�9t������3���ƱBs�29��խ�z+R��m$@z�<���}b�J��}�')},`;�1�^k���dW;�ěg��%��%s!B��N��Q�ݳ�&�k��9��\m[��r�@��7ρ9�?�=�D�"F,XQ�BC���R�� c���������u\y��ט�R
���nW�� ����*�u8���l�!6�cJ}|~]L�c}=�f._�Mز=�$J"H ������-A��~>g�H�,s����d3%d�y6����J��9?-��u�z `McS�;h,�_�O����(Ӧ��R�"<�k��P\q��"ѧ��㲞�?[�{���ydSŹ�r��M%BҕΓ�>JM�i��j����M��߽�#��3]���Ŭ�V��2����l�^9�?q_��s�NW���Į�nE���l�l���6�&��w�/$�hM�Fs�/��W��ծv��Y���]�jW��oݖ�Z�FQw{�y~&��x�+8�T	�*���V����1;x�,?�|�xxă*<�Fz3��K�wī)���+��+5���4�U��y1�[�|=�9	�كa%q�ۇ���X�D~ 0�ؗ�����kk�7=H>6�7���p�ͷw ?|�����mD^)�e}�1oz���@�59-� x�@��K'A�C�Z�&ݮ�a��*�+�;�g�o��w?@af�ǃ��#c���ky@�dU��ޓ��4i��n�R�+�Iː6њ�Wc�����ܒe,f���Wy�X�j��a�>FrQU%��7S y�d����(nj�;� ����U�W�L�8Yuv;3Ȗ�p�����U���"��qi��d��U�$DY��@�v+n��{�t �6�S�Vn�&���v
�f��.['�6�R�LslC�"W��cOv6)jY	��f����U�Nn�l����2�L�*Sr�1�xׇ{��'�/����`���И&�q���=�@D��(����;��G�9 T�"0Zw'����j}V-��.���2cX��+�4����l��BSv�O{��v������i$�� ��tRf�}�a�,?$��� ����s�����cw�e*˥J,��H��dW��s٘� �lh���]V]Cڹ�c�犈������h_풺Ӹͣ��n�"�k�����eCy%{���l���q�l�I�C���k������.y!�mj�e���h[G���F��l����ꊱ2X;ɾR {���vkLSzH��G��h�+��l����s�����o�8h~�>�F����9�k7����|Sڍ����~ҪkO�cܹ����M=n1�nOFd+/���$�����6|��7޾}�}Pz��8�]��䇿&��O#<$¬i�1H��S��`��[�5hU�B%���Tf:�_���i����vj�)'��d����jsPL:��l� ~���ONT�|K��e���p-/�;t;.yE��(�r�o�P �R���j��(�J��tq�^"˃c���*8��:�\ �NV�b1>��7���"�Ͳ�t|x����@�p2�'�?ẗ́����[�R?�*��jW��ծ���]�ծv��]�kK��ꚶA{�R��	�/�㍏�zN����� ��^N��ʊ��}<��	�_�=um��+�^�`�����������SH����b�����^�R����P��'=,&Ub9�#*�I*�[���kFlx����bn2���� 4V��fNߎN��G������Ys�1  C'e�Pd��q?�����*��+Y&mnQ��NV��|1��ʝQ�����y���-�f� �ȠY��ٱ[��U�3H4m�Z���m���6���f"�9 a_��Ǒ�ze� �ݎÌJ��su:mU��y�yn�������@��k�}n&!B ��׋�Ӳh��M)9T=�Vֱ���a� �/���@L�NtR�C��9�'A��88�L3��m���R�Vq��@ޱ�Ow�#� � ��6�`�`\��e
��+V����*�	p�F��G,Ϩ@ޕi@q�s)�ͮ��n�j��4Z�x%��n�r/���ȕ�a��9}6�^^���5���Yn����q�}0���*��,�XY?�����`��/+���g庈��y��q#@&Sek>��<2I6�;,������Ϩ���S��H�]���[��� �$�P��|/�kl�B��e)��U ��z����r�g pI�'��B�@`x�N�9���0��4ɓ�ˋ��j�=�yl�g���T��rPD�q#I�k;�[�8��ޠ2�EU?��g�.+e�:��!����s~$ze���&Bu7��ğ��rRu7�_�����3�09�(�4|���v�X�B6�\͢sw]]	VB�"��߄�9��1ϵAͣ�yUP��솥 �S�Y�&T�6�yW���? �yTO6�vr��g}R�q��T⚗h�ZH>9���� �%�)�4���k l�CA懔����2f�^L�	����կ�J�1��:�{���F��2`�V&'gm��gNjR�4��XNV��+q�|*D�,���5�g��/Z^}|>zN6���a�^L�P�ht��>� i^t�א��<����f���Z3�����m^��BS����~K��Iv�˔���w/����{߽�fug&�1����+$v��_�jW��߱]�ծv��]�ix�h����ff���vg�@�ǋ�^��V��� ��a�0<����z8gU���	[ۋC.�O���0�T�0�|�a�b$@-m�g���r.�~�˃��H�ad����uSL�w<�B0� 5^��y��@��������*I[������z�>��^��;�&�qCd��9�֚n��6�}�Фd}]N�N�gX�L@�@Dz��jz�em�)�|���8����cj��e�j�Ͳ`̿�@��m�!��Y #��H��+���Qƃ�RY�7����λ<�ay�JEZh�����n���V�͊�*˜�YC�f3⃶^��j���M� +�j .�(�Eߣ�v��N Y��$k�>�#P�d��ӄ)�Q��QM6^= \��}��BH݂*F�Ug�� ��S%�qʧ�g'/ �)����r�B�;�*!qq+?}߷ǁX�B} EKZ�[�i,����$��w��e6S�8��X�߃C�ez�˩�5��1j�R����F�F@�KV�M�S�z�5�a��/"�@��#Uh@%>_v�E'B��X�o����7������W��N��YK�1��;�T�ƀj���|�F�1P�l����V{X���6�m��8NNTqu��/ � +U��SZ0N$2<���������%�%��ۋy�=ޯSK��q�Ϸ���*�t��L�y2��,��ǵ��N:OV���?+:��Q�N�M��u���D�M�5�`��q�sVI� �2�^�gdI�sV��S^��4fAdj�i�'ew�w�'N|���s�����͖�?����]
eot%��yH��G>W��W|?���$� �c�Fn�J���N�}��M*��8���+��n�5u����*��ڒ�<�;ϥϏ�?|{��m~��e����~i��H�x��8�>LS2k�l�c,�RU6{>���0rsD�J�3���x5�����4�t���gBގ����H�F[H_�gzPa�k�^����Q�R��R3,*�ux2J�G1��8NX��{��c��J%1���`#7�����d��.B?���j���{ ���Z��tVHQ���=�vQ$�V�Vʦ�³B�L�� ��vS��>��c��J�ky����������r��]�j�v W��ծv�߮��L�h9��KO�!����G��$�O����+}>>-�Z�? �!�B��\�Z>~������䅁2Q���H��?~-��ۿ�I�����r��;�#H ���:��xʖ�@��x(����m)a��
���f�����Pw<�F�dJ�y�KZi�;\��O��ǃT 8�bՆx�v��[O��2��"�܉'d<���fd��K"�� ���z�kQ��U-Vm�l��[����o���݃NAl0�b7�yv��
��\��l�[ S7x���*̓)B��۾��Xz5�u?�ZE�
j���!�-����>ю��?��� �r�n�}t�
��� �tH���t�Z*Uw�~}83t\ߨ2,���n�ӂX�0�m��KʌU���6�FϏAx�U���X�%�*�E ��������W^�_(�:��=)���.D,�F������zJ�����@:�S�Ul��ەS �����Ȣ�<;[����ju(<`�5�B��������D�D~��u��i��H�7����ǋ*�8��s �"d2 ��~�f��ZF;U_�1�:���Uվvp����+�I��������s)g��1u�#[��\������=�����6��
9;Pݷ[�E�P�H�����w�*���s͏ᙈL�8���g'z��Hr=�H���av���l���r�:���8^�N�Q��y�>O�Z^I��a���9/�[~AI�N.���"�gA[6d� [a��C�fd�~ZƸ^��?�C���+6�R䢃�㿐P�:��+���E�!���7V�sL�X?C���ꄱ���Y��I*�����N$�Q����f�2��m
	s�,J+�[p+O�!K����߿)����i:[~i���k�1!�`*+`�;+��;�oo���+(vS�(۫��gIAnu����8Mۆ�yT�>��o��M��9�$���n�����S�p�N�2�B��{������O)���$��������^���"��[���i���{.�o)�\��S�-1���1R�v�]a[���n7�i7��9v]�5��,ɋ��J�,c]��׽7Y;� #lٮv��]�j�v W��ծv�߲�!��BT�R��2��XE(i�$�l�F�m�$��'$���A��fA	�`���|��! �*��bs_2�Ŭ��L��P����������J#P '{ox&����~V�*�j�-�x|U�HS��7��##��U����vʖ��ID�|�ú�2 �?z ����Zݻd R��r|�F��j$IV�)fI��ʲ-�d8c��V���Oq|�W��܇��[Z_����l�Z����������aO5��{쏩TXA���2Q�vA� ^pܪ�[#&�=�!�
�2Ɩ�����&���	ZF�P���L��f�CEG9�==�3�ѝ\��, =s��Ͽ�n�^��fU�v~�oV�W�:n�H��Ϯ�A@�`���<LX�Iᒢb_@��VY8��b�*��T�|f�ڹ��,�*A��>�)����	,�|{=�B��f���+�@��#��-��I���ٺ��D�a�%[H}����Sx,F�����eA�y0:�s���l��BpߟzM6���=`�$-j����3̸��"sXU��}��[kc���/]���b���į��4��9��)Z���zض)u�
�P[����]`
#Ch��j�)���@���}�MM�I���mVT�ʆ	�5�T	�B	0���4�0N���<��y��8��������Κ�w/*�q���[ئb1�C�yɦV�yV�S�a܊҃Ɲ��{�l#5f�H�61d�-�,`=�~LqN��^
��]�'���ؔ��m�|\T�$�|�5\�:oۉ�9�>���n}w,qv�D?κ�x��[;�\���Ө��l�1W�I}7'�缙�ګ�Lx��B��c�NT�׷j�+�`��y~��9Y<����B-dA� ��fh�ԳQ�Fx<�l�p���=s,�������Zژm�8��=�M[��#YGP��4�����C8_y����U%c����T�$�j��Nj4#?�ѵ�~ɾZ�ᘹ�q:]C�F�>��/�첹��y�,��^�H'��C$��{�=K��cn�y��ܽ`ɍ{"���u?\��h͊@`g֌�G����{��c���l�������z�����-��m��=0ڜ��u�٬?Y��r?J��gW]ʹ�{;���g�q����+�jW������"@�v��]�j�U��P}�j�������Ak�������%�����Ί���<9+#��WY��X��~6U�2${P&0�"�Ƶ<��S���oP+1�?��T�mG':���I�Qɔ$����v�I�úb�C2�� �(�S�3P��P%7t��� k�|>v�h��6#9hT`Y����4�]BN�ZS�XCd߿�� 'Q�v0�E ,��h V��jL�?� ÒoT� �
�x~��La��^(1�k�5��l�0�Hă:�sN�i ��A��;u%�63}ͫ�I�~��8���,��(����Z�W x�UV����l����p,ݾ�i 'H���'��3�b3���e�dۂu)���������7��ɀ�#��</�.R�2�_c=#���#�J-�+rP���Ɯ"*�*�	�}M=4��G �[eSO����d v	�,<�(���勍���S�Nl�}=�]��`k^ٿ s ��I�8��&pߕi�s�$M&8N��8޷EA�ڎ�+����T��j��./~�.�,�^�n܎��ۍU�;�/��R�v\���u׹+����f7�zh�"+"�!x�8�߿O��5 v&=wvq���[|�-W�|����M}%����1����L}�1p�W��F�d۬�M�<��˿{��iR�u��Q)��3M��ٯS�l��1]?gX�.B�@\]R2��e�8n�Yj~�XZ�<Zf'��:I^���-����>Z>v��c��_fA�b�G{��n���_#�X1��i >�u����YAK'�[��}��P	2��ͺu
}3�ň֞7��0q�[�+�R�=��h�ϐc��㼇l�I��3'�G҅ ��*L/��^���ɏ�H�
��/w�u��f`��8w>>>��PV��:���9�A"�H�P��~�Q8����U���������۝�p/�
|;,X4Ϡ�ч8מ�ؘ[�U��)N^�?�y���>�0��������_E,�P�h�v�I#����;	E�m�L�7RT��~U;UZ�a,�4u2lT��}]�ׇq���s<�������!H dS��~�"/�+��3�+Bd�3�bJsݬ{����������_�I)yvG����a�#Mm �®��ٱ�*�-�xΡ��1H2����؈ ��`��"v_s<P	h�"��ZId�`��=���>v��]�jW���� ��ծv���V 2' ��a���S��P��[ Nxhg���������퍥`�X�˪=o���x�iF* `�AS
d~XǷ]�%I�D  cD!�zH%�����{ �ݲ�� �&F� �<�����{3�H�ϷĠI��̔����������nS��H�tWU!��o7�����#�����\�g�9�^����"��[����k��"i�ˢg���"\z���>��ӎ1 ���fU�Z6l?�@�o����� oV;�9���.2D�|�F/�I���o���R� K�Q/�CcJXU}�߬�^@���#��2�y��X!��Ab<��"cdƤ�W�'�)'n��(���8�G̓o;���6�8���  H 8���ql��,����� �Q�e �ȧ�����u�B��{�S�9��
hX�xe=�*�S�I�n�3��c�����V�1���U��R��A����@����|n$i�mX6����K ��Ŀ�}$�hߢ0w�>N�������Y���x&�V�S���7.���q���ˁ�>������m�+� ���ÒI�\bSg �%K����Ɯ��������,i@H�,0����H���{5�q����*�@Z��g�\���c,Ѧ�H�s�k�Be���~rOy�.��i+�׉s�f������n�,��c�6�_�+���c@y?>y=`6E���{w�H�$�4N�9�_��x�Ϯ�;{��	R2�%w�O�Lc_��<i���q�|(�@V%�a�cnz�w��� 8#�tn��?���dǞ��R�����jr+�M�*��&���<h�1E�*[)G��Ĕg@��[&C� ���>W�w��Ѧ��5����M}���$(��Uu�|.@?�P�g�@,��͂�yl�vǉ��L�W���
��e<����[��!s��Yd<�A��i�1��C�;�'~�8��+����^�l�zu˨fL��Ö�HTl��q,��z�1���g���d0O>m��slog�	�}���)ۨ�5�L�R*�pM�x<��P2`��l�� �����ꉤ���au|����=��T��5�F�;��%��#vd�Ttw�|���0WI��-_w5����B�h!�� �!�ݫٽ��y"50O��������n�"M�f�q\x|���ղ��f�s#qc��y�{�y~;��"���aF��jBWMp{@@��h�B%�c���-��0?B��v�/����G^NX���a��n� �0@z/|��FK���Og����#U�͚t�d��p�����,�FR�����ܥ �9Q��o�ۈ�o;��fcz�菫]�jW�۷� ��ծv�����0$@���Vin6
��z&�� �Bh5����FD������L`[a�[T��/� ���F�&�p��I����g���m$� �O��� �rƓf�#���"?NʊTb9n�T��[��{1+& ��޻���-+�\U[C��
�����n�1.Y%�)w<;�L�� L->�sQ��j�

�"<�=O��ɑ�I��,��A�yQ+ _�eP`���2�9��|���2�)6	`C�f�5�lk�V�d�. �Aϭ����^\�|�{s��hTڃ[�?��*ś�p� ?�C�YyU�pQ�.��8fy! �Y��^d�-w�K�� k���$Y!����@�8i�~h+�d��r|��d��jpel(�@\5�!}�źd�5��{�q6C�f�FX�d�� ���g<��c�nFʠ�jT�+�Ŀ�p���I��"�����:�J���z��=-Ȋ��y����,�R��va��m!�[����R�m,OQ��1���6�(�ʞU�CF����c-���J*UDj�Ϫ�,6!�N��{?ٲ�tW�� ����W�O�#�M�ذ,ڥUS(�a.W��>�PVN� �\������:@�}Je2	c�*�eq�L���A3=c!}YmϦZp6P�:ܫ�]E��	�-��=�|���R�����a�����`qVțb?o�p x?)ܔC��-]����N�m���4`Le
������)Dd�Y%&t�^��vr�-x����s��+$��6v
(��M0j�c���[�l)���i�ur��I+������l6<TD {�6�x�1
B�H�-�� !;��\�AZ�ȃmR7���>w�z�0���u-�c ��Ȍ!�$�@���Y͂q��1 H=������#��f��ˡ�j����2f[6�O������}��|�E1UE��F"�3!��/�u��).��f��i�~IZ�(ed;�p�R[5U��_v>z���)S��/�c_f�O���.O�2u�1���s��}N���1�s�󘢯��
,�D5�E�O��(,g�O��YLX^�b!�s�nV�T��b�
��t�J`ek�#�z����uj�w�L��+���������5�~��o�x6x>�|���|�Z�\�jW������"@�v��]�j�]�/U�>Q��'.\���2�b�VY����j���h�ܨ��� Qa����7(g�"�������ni�\�;Y>���:�����֫�y#a!*��߂;��[8x�J��G���.���k������f dv+��R� rW�H����E&��g�_O�,�,М�t(I<,]�E�~��m����-�F{1(����멏��8Lx��۳����?�$@�p�-�!�]�j׭��p��vU�I�#�׍���;̹�� 1�����3uˍ4 #�*�B�� /wY��z ����f�a}^�{ ��aB;�i�� ��?�eFJ P"R�j�E.���3�\5�S�ŪB^�o��������s��0;*�P��1�Ev
���e�x�hX>���5JY�{ط�*�������%v�M��h޺7�d��(�>@�����d��HY�t�(�H�x6 ��`�KW���mþk��8�'v�2`�E�]���kkaI��@.	
S0�OA������U��ط�TF���*�f/Q-K6IH���,��C��
^+-V�M��㒩V���\p\���Zig�"P~Ɣ��
��a������xخ�9�g���)���0o?�8vi�i=<F��%�5[sk�j�	���׈��@F�nސӜX:�#�Ӓ��[xN� �b���e���I�����0m8M��q0��o�ܳz����	%��]��W~�����:�O�r/�*�5�LAp��F{��jI��X�Ϯ��:	9(��ٌ�n�2T�ZZQm��{�}9Y���eY�����bI�i脎�'X�O۬���{�gI��H02���G��� ��d+͚�dkc���5?��HZ�vF"�� q}�WUyDn���Ef51;�#�AA��^U�������:9��7�>T��:)�*@'�E���k�6TF��~�2��I(�'z^�__��)�N�>���j���H5f� s�m��'��.�,.oNq�T�A��3�E��Iנv�K.�[RUv�V(B"%x��a����S'3�����S��C�_3L���zf�,	���W���^e�x�����Jx:�������Р"�=�
1�p��
�ԯ���*�K���K9�2��*�TH9��O��mL�g��p�JSKP�G�z7�>0lx��5FA����s~��WT���E�^�P]��nmk[��־ym#@����mmk_�v�᪢%�<����b-�z�s���}"� |;KX��X]ݔ
|�����_�	����N�xM����HW��\�/D�\c�a���i�?�V,��"Lp@��%��r:Wʷ�-" L�Ϸ%&u���~b �x���� �"#���<��kET\�-�l�.c9�� O�����
�&����X�u�<J�pб�5�ķW$3��N��k�/�ȯ[��f�����*���dQ!%���DR,��4�� r�p��'}� $��D�xP�����v�׏�D�Z5-�XWᳮ�P�k�U��[s���o;Ns������H�#;2�����ÜA`������e�d�fU���������]3'F�y�j|�R���и��K���xK�^烸%��v6����<���"ATHqr����ba2�FZN�U���BNi\6�'kTM��<>�T��>��ue?���9�Oa��r���e���6b���'���ϔ �b�D��y�V�\^�	v�<�2?#��Fe����>[e�8�i� ��t��s/�h.�"u+�c
V(��L!�`��4Th�|�=��Y��Q|�jv,�~���dևn�x9���bt�>�9���j�\��P�׷�>��Q�a�j�1u.7�|[���+�/��|��=ķY�
 ��}트.�
�\Ɓs�EuQ$XF����t��*Y���ū›3k �MP�ײ�pͬ/I�ȵ�w��q��	��ѵ����2F��XH6<M�q%<}uM� p?�%�C@7�izP[N,�Gc�5pE�:�g���%�5��1�Jc�'��]H�8��ß���{�k�}�9��so�u���}�^T�{���HD� �g��� NRy�/�W��%/J��"��C����(�����b�㒳q9&e{U�r����#�?`#��D�զ\��������L%EkXZ��]�H#�]C��.
��q��]w��p�<f�X��}���e�o��?�Sa�d���XҭȐj�3�\/�[�q�p)e��قlAA&�?���m��kZƽ)c�J���&|܄�$��P�X/�����tt\�k� ���X<�^�#��2�f
=�B�T�ڒ�Le����ҭmmk[��7�m�ֶ���m�k׎�#�M* ����(V;#����.T�&��讦׽�~�+/m��HV�%��K���qg�}ҔV�P����� �R����tAZ<���|��Υ"�� ��{���.1�@�
3m��F]��ږ'{�����Ou	:g&G _��I'2.6H�k+����+�u�1�<�� �$�GVݡZ �Q�ǘ.���lvZ�F�Uv
��N.R����s�pֱ�G{{sK!�$�EQ�s0�EQXX�I��.�KK����VU�d*_f9�$�˫:�_�/�N��/��bUS�M����+cݶ��P�����*��t��g��X���B�U��L�1[�����x��=��գy����2&�@0爗�ni�Vmo�n�e�Ʋ�Y*� �B�Wy3��^�ũT軒��P`�7ᶰZpTρi�����EAU�ng�M�`��l91����)LQ5�*��F�����.���e�+�O\Y֑ 2<�����>�j��N0M�IҴ���uv�Cv2���O��������hjLR�d��h5oz��Q����|#���v�ee�W�w�w��G��βT��9(��E-��f�& �ڣ�%B�T���Z��;�X�z�SZT�U3�d���E�2"�Dh!=��M,�m5���*���}Օ����d��y^do�5�J�B�?N�ݲ��X֥��b�<?�I��>���=��	�d���a�!h>z��ʠ�6t�rZ<?G��4N�|��gZYH�D@^E�9"g���w�p8�OΛad��ph�W���98��\U�;�-C��ö�a���D��5���5�+*l�Ƒq�fZl��WEY�JV뷵�t&����z�H��Ӆ�b��z����v�e S!(u��T2���6����1b�Xg�C�7c�0��)+�##����C!&��絫�D��|	�(f}-�6Ḫ���``��ddI�yۚ�p��B��=L$�ԛ�j<���QȱČb�_��x�/W���g\q�h���aN~��gVS��l
��ZeD�+��)�J�I���A
[��:=��г�cQ �cIv\�����\��dU;S*d��yn"�Q�9"�J�cĈx*�� l�5��]^+�>�3��)�C�y��R������H�R����tk[��ֶ���� [��ֶ���U#3�Z��O��Jrf,$��t�j3s
c���ٽW3'�D�����۞/N�����.(D/��(K�T�^���:y��b{�4%�}��j���+έ���p��ѲKl{����un�_�By>�ܭ�7�+Q��q��Iq�m��������s.�ؓ�����]��Ý���$%꩐ �����BX`B�X��<�<F{T�xH�X��F 3s`�T��A������9>�y��_c�<�����"���&J���@ݴ2�����I�y���������Y�W�Ÿ��w�l��y.����Fޒ�ޕrt>,ג���.
8�6YU�])�V*��Y�e�5�J8PS��=�c�1.�?��C�I������Y��h����#�Vݒ����B�����U�Cm�J��Mӟy���X��*�m^���y�S2��R1K��S�U�I�;QY������h��X���x���U��[� �t�Ӏ���v]K�4 ��O�@a4�|��||�5@�\�)T�@y�"�
i�5H5�d�O�= ��~��)�_ȁ�f�& O671�p1��F��ޠb�+n�dսȠ�m\x��CN�����6�|n�%�CǦ��J牌^'%���u���Tl���=��YY;y��0�DE�'��Q��9�<�J�8�[��Χ�V$���XKh��{���Aħ�{�]T
�k˸�uF,������@~4U�C�+�-�TiP�c(��z;T���~�~K�{45X\��,���JNj�3ù}-�;AF���r�E*��gn�4KF4�:c	���m},��Y��5Ygϰb�,���~X>LF�y]9Ѱ(x�i.kòV�y�iм�������Z2r�&��y�p˧ԄB8�5pB�-���^y���/Ma.���b��c��(Zk�����_�r}8~-�g��E-bE
y�HEh�З'�d�isY0NSyv�B*&��OX@�U����U��ܢ�y_���?��zK���T�E}�ܙe�u\l�ܒ�mUi�6-Y ����uˇ����ΔIf={%@�֩�3�[#6�)t���L-2���*̞o�%�
�ή���9Qϯ}?�y��mQC�w(D�Yt �Q'ު�0���������>Yȹ��|���{�����K��ֶ���}��F�lmk[��־~-.���k�y88���f�[����mB_���%K+�Ǯ��k��w�n�����p�Z�KHl9��Ն��n�b��uPA�ßT��cFv��Sy3ƿ�e���M���R%������X���� V��܎�V@i�K�92 :O:�B�0�R�/�+��A�(q��8q]V&� c)CBҋ����}h����f���^��<�/�U�"`�e���y �^��u3p����O�izլL��&����(E�����Vpo(!�勸���R��)��U*U���S�rV�!�g$,��u��U#��t�ͦ"���5,���@k'�{��sԟ
>��1�P9��Q-�\a���|�ޔ�+�w
��K���Ti��V@眖��LY���.�{=N���~J�li���/w�.D{��*���/�`}���
I�X��Ţ&Yf��Z��������B���__.њ| �֣�ݪ�+��,����8r]�\�Bi�_B�T�qD�[������x�;[��d'�V��0_@��qTmqޓ�AVՇ���R���гD��`�F�X%����E�ŀ�X�%�~�<����r�R���}\:0-U�,`����Ul;1�VJ,ė� �6�es����usvR�~]�n/��⡊��V#T~�
Y���jmkm��<���W	�Ř�xb����Ҿ�|/-i��2���B&�9�B.'�O�b���5�L�H^� ��ug�w�>�sLza��?��a������Ơ�����o�WK:X�V>��,%W I��t�|�V?�KP�7�,�� g��Ȏg�����T�B޿���3�E���v4�,	��	e,���"(�HLE10ϋZS�'��r�&˲rNd��ұ,�s0����:��P���!�BWcr0�{��5Z���	 �0b�/I���d���%�����˟��~6+.<+�5��� p����#�Ty�֫�<��8�z�Q�x't�"�DS1=.���^2;��I$I��TMQ�~�L{�ߍ�(�</���(�4�H3^�ѥ���3�2kʹb�Ȇ
RuC��"�q����ĹT�q΁�l,KȈq��Q!��I�Y���(��H�֖����ֶ��oj�V��mmk[��ק��̀�h���K]`�9�v>��@&����V�߼B�{�I�|����������z����8�~<�^]ma�����oN�����"&�h�t%K��1,�ƞ6�!������"p�T����"SQv���='ۧ@�4Xf�(��q5*{�(?�c+�g����e/���(_�$[(԰���o	2gu"^�+JP���`���j��gk��G���*������E՛M�,�3.~�5�p���[G�c�K�9\\ۢD�
J��P/�v��� ��U�$�Y~�#�5���׹���DuL>��X��/� �ݴ�j�nK�`2+ăYz�hj��NߚK�:�p݉61 �L�i���=����H�� � LS o%�7��n���|�&��F ,�1����|�&ި�|J�+�
o���[�֗k� %�C˙|n�*�yNS���9�ۃ̢�+��e���.T%���A"�U��^�늎�^BΩ���y�O$W��ZP/�-���wE��9v�T8w$0�窐y��:$T"�`s��F������E�~�ۢd�'�:U�J�d��s��ݾ��
d �}��U] ��8-`nr�2����⷟���C%�1rW�e��9�{X��46�<�3�|יzĬ�0NS8(ؚ�܆I��D�A
%�c=�'ml�
d��(�&���l����Y8�z��vϝ!1d
��H1�˭�튕�<�9�p�5�-�<��(�\c	�^�*j�mK�*����c̲��}�<\Y�c���m˹����jlv[&��q�������Aa���Y�"��@rM����5:�6�0����������e�[�q�F�N����-�+'i9^�;j�Rܖ*��>�*HVU��C��=���՚2�FN/�6�Om�ֳY�-EV{&�2=�J�_f�d�>�9,N�`TM�4��*E# APr�'%Pɀx����ǉ���j�b���U��lQ�9�3���AUx>����<�;ˀ������_�6�܋sQk�ngeE	TlZ��dyk��IRx�9���e=���_	d�J.�lvjN�c� ��״q�ʢ:����|N���䄂��6Z�qP�Y�(���ʇU�
O���[*�j)�Hdq6R9A�H���LF,*���	���q_^�Ip�gW6��|����e���!i����N�kLOr�)*�e,���A��~7��Z�����=ל
u�g�+8���y[��7_}����mmk�̶ [��ֶ���mCE4@�Oa���O/^*���eP��_zvm���ه>�$)��ߵ�p:J���H|�ܞXy̠�$�yxC8���Y"��wSL �O}�����\���(�B	�������a�@�������~��������ԛ�Hl���q�[X%*,�ܪ��.���w�'(��cM��d�,��^p���km����)��F �ʈ�)�rl�,\U�`�aI���9Zջ��N��`��9�
J׻r"!PWR�4f�00p����,�Â�'�,�Tm�� :PB[��_��|���^�1y5�.�{�X�ш%����0\�V���T�`b�s����c��{�=xhv���
dT�6;�
���zA�+0eځs��$h)DX��g������H�.ϫ���Q��(��AT9��0Y�,ຽU���*�$hxu�Z\7�͕(���5)@f��������{�K_ͳ��[Fc�Ng��Y"a�G��*���F~`�T5� ��L�}��7�n��T?�͉�O��_�W��m^s0o�y�co�M@~E�:�i�
xT����.����9���T�F4�"	Y=M{�d�0ɪ���y �<'�c��0��{~�M	��zo�� w��r�D@���`���Pٌ����!ϛ�&�bX(��T'�h��`k��JI���J}�W���y ������n��C!����$�0&wy�?��R�=1������y�wE��}�aZ�5�I=��H�1;df���0����u#�c�B��@r���2Շ,�5:����\�:�k�B�0�y"'�m@-�k� QW`� �f�������Aw�x(��~��S22v�1�yo�D��\�E�t{<qMĚ�no$P�*,6p���F�"KV\"�H����*��\Aߙ]�[��3 ���zt�C��Ng�#7!�q{�_)�	��"�e3	�a�Jk�%̼������M�H����_C ���h�׳ʾ2�*��#�=�Ji�{�Ã�D��BDa`��ު�,��D�՝��q}{s�}w��ʫH�Bѽ��P7`����&�x����c�Ν�FR��jwP�D���|��������Q�C��Y�s�" ��9������nQXẓ�\���=�$��j�@i�$,ג�us�U:��,\$$@	�s��&!,*�$"7��m �D}�������k<�PmY�0�y�ț�G2O�<S�
d��R؎�a#�J��TTMcF"x��2����Hh(bs2{8_g0'��3�)L�]�;��q	i�z��<���B��w&!����I\��g���1t���4$e�4���=�1�Σ�a�F���k>[�!�̌R��Fx>���!������B%�1=O�\��9'��e������B<���QS��䮽��k�:&lmk[��־�m#@����mmk_�6|a5~�\�$�y�8;�f%E����jmQ�MP/��N/z r����H��a-@~��	�x�I��&"�C�U q�֬@���˵j�+��cys�/txa�GT��"UA��(`*D��;�v�<}p2�+Y^ h���Kg�W������N� ��*�5_�i9�*�UF@y�X��k(�.SI�a�{��e��RQ� �9�@��z�;�D��9u��nnde[f��Ƌ��{���x��P�"hɃa"��T�c�Շ+[�����B��o��ҹ�w�>����<n��ߺYK�I� `���pݡ�Ǻ��c��h��'`�m4? fq�����{��(XW�G��TZfM�?Q�EچU���B���b̨b^�P~�R]xI(3e��\_��jy��Ke���h�LE$�IBMK&�U$�����1�V U?��N�pu`?��>w���|��"�t���ӑch�u{��$)!�3�Qs~*�,��ࡹ̯�1�R0"x�>��� `���S�J���
\���O�$�ZSy�XzKkg��<.�dK�������k'g��-��Z�D���sM�K���LU�F��̢�KU����U,vDu5�"��Ϊ��2Zd17D�X��8�������@��'�� ��Ȧ��ñĝ��+ʬ�?E��U�U[-{;E�y�Q�0�R�|x�7��hJ�d��T]P��/�������=�u��
�I��[aކ�o��M�J�&�Q϶&(��dAݴ�����4�����V��>��AǓ^�r,�;SΡ2U#�}_�:*�"*|H��<��y^��_���������Y�ח؄�6zu�Ƃ[Q"Q���e[���ڏ�UZ�H_3g�VAӅ�J�n&�z���8k�-�l��ן)���ā>���˻8��6f-���<�6
�0e�z������\���X*V�?o��A�\�f��|i��KRT������{E��.U.z�oh��5@�,Y?u]�2��Q�H�R�zÕ3�2ZO�\�L�5����N�PR�)s��IVv��Fy(�Ɠ{Ԗ=r&=����9 
�lQ��q5����&��\]Y��䆢�c��̒�R�H0S�ZaJc�Kf=��!�e/���q�Od�R�{���<W���xVdH�NX��d7���p�*��.��������c���l��(j��<����ޟp����ֶ���m��6dk[��ֶ��k����_lhWs�� np�<�b���J�����
�YP�C��.,!��4���X8��PN��ﺭYն�/Y��]�J�ƪ���*�}�{��l �m,/nK y��6�eU\� �)\ne��y΃��.�	�]Z~*�G����X_����܇��>ӕ�Vć?n$���~0����u!*�*X��'~*����y �z��z�sK���a��r��Jd�1>"j��fҊ4���D�T�+�Օ�S/+2> ������a�*xɏ,�@_�U�GnD��O�DP	
ڮ례-+��A�G[��,�Y��P >Yt+|@��&Z��E����Y�|�aI���]�Y%��·��@��.�	�3-�P�5�Xh�g f��	�[��Ve��
���W>��^�)9�V�/i��`���>�>��i�ÿVc�jf1�αȒ�W����5UV��
�A�)H��H`S4��9�w�'��j�Zg{�H���Dp�X�= ��2������ep,dcp�66��1J���p @�0��P �jN @8��R�(���*�E@qwI�ؤy����E@@1�[2 k*�8���i�<S#���$HC�U\#\�����5E��X@Z�}��ڪ�eq�����dܚ��gT�<�-���XI�'bn.*%W�Ae3{���f����&WT"Ě�"�QT\�
ё�%�W����[I��6UQ~C��:�+����a�	��V�4�#����W7Z;��O����E�A�I"e��Pǒ���B��J�H�dk@�\�g86vR���2��3+�������)�3�-�_�>�s9q?H���7�Ofϟ�d��k�HRP���zO�Mn����5G#�"�_�������G��r�J� PS0J�3��*L�v�)k%Q���M�KUH����D�渓�1x�
Ǽm��s��F��ɇź�h>F���<��+|\����ܱ�x�K-�Hn�U�]l�U(�m�n�Y�O�~�=1ٵ�{���pC�-��bJB�l����#�1no8������~���M��c�
V�GZ�KK�s��y!�׏z�Ӝ�T�
�K�FVf1�bU�D沄JE=n��{���	�]�-�%�M'�K�}'Ph*���b�R-�/��&����5��ómm�����<���q��g��t�l����������,���F�b�R�]C���~lmk[���m[���mmk_ˆ*��¥�t�=��:�^�_�S�����ﹰ��K��E�k�-+ǉ=�R�]�g�Z�����b���,@�9��@D���?U]�R�WЗJ4(�v0�T��%*؊��4#P]m������2J.@z{�P��L�П�c���@�@_�  �1c�O[w�
�{�Ѽ��g��p��-�S!;�.v�*��s6��Iq�q�1,���~M'�QyT�ZM	�tP��p>�<Q �����g2�͋Ye�{�N��FSg��fZ3�}>�sP�U�U�~:�^{��<�]�S34w�U�V�I��Z������  �� :괞C�S2� �T���*r�%G2��t��Z2�Ǭ*|+�X ���^��
�[_�� �3OK@pe�T�y��2Bd��g��7!w��|��r��c��ס�V�	�aM�?�޽�a�4�R���y
�m7 ��4��:�h �TT<�(�r��}	�^r*�ٵ���V��~	ֿ �A��~�d��Z, �}I54��Q�*"�W����Vs{V�� ,ƪ�)�L�� U'˕�SE�C�Ȇ��㴧��� ���$_�̶e.J-]��F��X���DJ&- ��VU�;i�69R�%��F��8.����'S��Y1Z���# �δbdr�M���\�9��z*����x��'�N#���?[���~�]���*.�)s�$^2b����YFRf�bk �L��f
�C%��XМ�uE�W��B��%0<�2c�GZT�տU%>UʃI��V$�����p��"����ȁ���p�C��d.�m<���3�Ґ��,$��-�=��	�zZ��V���\���f0�G�'f3��R	h�%���	��<^�J��y,�?@��~�9KA�^�N�x��pu8�vl��c�6b�1ŝ^a!R���8��:\��ϫ���g؜��� Z^
�����x�� ���u��8�e,3�	%_�vo���v��'�N�.�	��,WgQ.�YT�9����X�b�Df���î%3J�K�Q�WP��ި�;{֚P8RY�BE���.�2Pp�j�Ѳ�:�Y�l������|ڝ�T����%� �S1G2��|��G�:-�r�\8Y�O���r�d+����+�-�T�E}2��ɮ3Ǖr�����-,�v��:�2	ZQ����?�3ރ����mmk߼� [��ֶ���e[��P^NX�j�X^04H3%�F�)���ޘ�<Z ����2�ϸG������� /fc����j޳!V���;@������Pa��^	��r�\�l=�,
�-_$2�<��=���!�K[[j���1TG�|;�s�C�Q�8�Q���=��Ƕ����J���B2�)�8j�	=�����`����Z*
��?��:��ŉf���&��\��6�Z�A�[Z�3I5Y���������r��J~�J@��+���Y� �%�B���H�ݎU��* %{��n���a��V5�&��Y)m��𚂸2�w���3�r��V���k���U6Tb *��;A�X*�i�4[���֘UZ������Vj��v��X�z�X-o@+2:f�s�����U���*_�b_�V�t�k���Xm��JV'рC(���}|:�y��ܹ}���1�Z��8��#�?�x�w���w?��,�Ud���� ~�\_[���4�g��EFe@j�6�3	^�w]	T#!:{@2����
���!�h����S�%C�0�g��,)�\��.���W)�-ϲ��lVk=��BcU�nF4��l��Fv����q{�<N6kf�$� ��W����0s���"�@�[�F:��-Q��ǥ�,��$1R7�8ןq��$�u��d������o�3T�����5a�
���([�J��
f����e��q�틐�i�����ټ��8���{���i^�=]@u,}YY�+�iL�Uj˭Y��24�)[�\��9���ٍ �%��x��T_3���>I[��H�(�#�}�4�j*j���qB��7��v��Oi���a{d�z4��݉Hn����wDc� ��	*oX�x�̶��q^{ZO�\"xl�,���n*Y���	��V��������'��몬���9s͒���d$�{�d�$�''e����Fb��Hs҂笮+���Z�Җ"�N`��o���9:99-
�Q�T�ٽI*Ց�����U
^ոZ* ��X��'�Ȝ��`�l��|m[Գ�Nrѫ�*	��"��6�H�۬��/����l�O�����md���e�ՑYD��0�Ύ�sb��yW��o{� P��Fsr8,�)x>����C�֋��8����f_>�"�9r�P41�dd^�8��M(
%������3OS�2�[*��=8��<K+4��:�[���U蕭mmk[��7�m�ֶ���m�k�d�C3�X�:�ExC�'֢�+"@��uo�ܺ���*�R����Du�hE�M�JU7��ZlR���*&�"X�캺�����9^�{�gu[�
���#���s�7 !���6+����߼�F&���ߞ���g��1�]p�Dc�,z̟��؊��v�/�����r,k{����$S��`!��"����^�7�~��5�9wk�u�	2�]�[K��؇K5.�V-F_��Y����d����2@�Y}�6���@q�o�j�]�0s���a����"���H9��͎v3�[kC���V}�g{ ໬�u>���+��y�V
�������\�LK�U�<�]�[���U�W����;�F~	\�`U��뀙��&H�'#�f�5rg���۪�i'&`O��Q�	��.�j�X��=�G�1���R��%�9:jkʑq5ƙQ��~�fYɯ٬b�+@<Y�*b�P���Ed�R9^r\��Z���i��G�| ���H�B����a������%��[�HeE�,�	����{"#X�+�5Y�.}䇳�ڈr#8�B[fxS�TU[ a��V��R1O��$`�mk�U�e��}2Շ�:{F@�Bғ���R!&*;w�l�k`{������$L��W�>�ܙe�9�{�8h���Df��(�vTx	"�1P����1�4�"�5��)�f;�`$J�U�ue�,	G���8G�u5�sHP�i�%�;���2t�]��j��Ʀ��P������?���lՔ�R��X'0�=�7����"��n����${�z��R�%���q�����r vO3��N@
��:��d ��s��D�yk��+<c��ӭ�󤴀͢����\Ӣ&S�E��!LV������	?��`;X�B�,����#�2v��Z3�|*,PX>�srR�U4ި�AqG�u��j��m\_������]�O����!�TMԴ��ƹXs�dI6��<� �U\�9�u��ZjL��B(G�So��bW��0@�߀FH���uU�ECM�mM��d�õ-Y.U�GLQ�C��x^�mh���1W�5B����ճc���S�� �[
x����|>�݁���$��9Wm(��: ���]ۭ2p�06hC��됟���?�J����w�[��ֶ��on���mmk[��צA���j��Ń{N���' %��o�l���|?���>��6 �D��aŘ����W����R(�Q�W��2��3���� ��R�����X��-d�"�;^X:�� կV��N@��%F��&*^��Y��zy�� 򅵕YG�ϕ�a��`����J�JD۸��>\�4<b��f�������Y�ޡR�,)��u�M¨�w���SwE*�ica��x�F>C�՘!����)�'���/���� 0�v���L$�@@ O���aZ�Eƾ�H�ܐ/���TR>1�;zXo��k���(������Yl��g/2O�H'o��9ĎU�sP=�!��cp+�q�)�G��x����+��<_)@�Q)]�츰�u{!�j~fܴ�e�[�:�L�m��?�eU�+Z��B/�F�E��ڨs��@�Է��˂��XX:P��t������;:.�A���;U�.��K�1>7�o� �L�`}=�*@����[V׺O�8�
�4�s�1��Q�v�H-���$�'�1�Č�!�@��u��`��i�V�9���Ѳ+
D:��V�ǁ�o��g��\ ]����*맔\��A����n�����L��?욅�>��V}����+��R�מ����[�a&�����ñ�k����/��q	/
_�W.�;�"k����I2�Z�p�t�`dݴ6�m��YV#,�J�ը�Vc�*�vh�� ��)��qbZ�Y����V�S��6b��+HaE�¹����MM$��3�Xs�3@F�$B(�r��.�y�D� �b,��q�ro�-���k�|�ML%�di!+['�wx�������n��tIfg���Yl�<߅kk���h��*�F������8��f%�c��h���ո�u�ur�Z�WT8_��^��ɋ1)8��8f��(ҿ�D � rFJ�Q�S��5�*�5Zg�s-��Be��X�WY��S޺���<�h[�g�U���'��Z�	�(`��C�\�5�2�|%����j�2�ۜd��bX$��8峄�k�����>��stF���Ty�s��jfQ�T��
k�T���N
�)$��渧s�'����Z6l8ρ9Z*j}c��di�̖�d�Hr%11-U+|�u�MQ�Jk�0�gpf������&7�+;�Ű�Y>�dd��f��fQAu�J��Cx�ҋ6��ֶ���m��6dk[��ֶ��l���!��r>`-�W>��4f�b����VnӞ$����f7�^�F���ucpg&*|���@9��w��D� ���@�{�dª�ю��l��Sj�I2&rk���M�&���W�HCI~0��7QJM�f�E+�b%����]���b�g���s���R� m�q:���C����i�.b'�g�et4�s����J�B�lV���@�mT-U�W�]x��6�ֈ#N�M͊�^U�
�d�0І��f�Q�؅�� ��9��T-��� ,{��:�P��� ��dc�	��#���>��l����d�~�h�.TM�C��N �����>Ae��	�fӅ}�V*/�6pnf��h@#ZeU���$�� Pt?y'H, Lp��/YU%�}� � �� 4��YM�SLm��*� !�˹ی%(�A,�'H��]�䡶�?���U�Nʸ`X8����6[��E�����6������a�4%�A�����(z�޹��� P������ǈ� ZxX8k���g6髰M��Y�/~���às���ͤu����?�Ѿ�!�5�s th����p�TsG$}3ǌYL�z��j�N�/�m M��~��05�
�������k��}������,���k�<������LU�/>�7����z��� ��]Ǳ'��@OcJ!'wTq?�m�f#h�b��/@�Y��k������S!�|-'H��ˀ�hWK�>0�%�C��Y*5�7T4���]�v�Ea�sr0��ۇq�a<���켴{Us�Vt��T��,���&irŌ�A�RKpUY�D*?_c��d�l�W�^�_I^?����Y�hj3=��ʎ�a1��_81H$��P��>�@m>��r)�N&�]w�q>Yi�4�r�Ǽm��2xdG�5*	����=i�7����B���E��nH�{�O*~֊�� ;���H�@F�9Q�t��d���:���l���Y����J�X����T+;��
	riwIP��i�{�mA]5�Κ�� a*#O@���:����8��$j�ˡ:�穲 s?�h�\�?GZ@D�UFTCUȏ�	�r_V$�g����os�^��)p�.		��,e��FI�h��05����^d+������d����&��c��΃����Ģ(�L���3 V�N���;=y�|hi!ڔ̰HҮ-s~���z���g߽΃�*���Bt޿� lmk[��־�m#@����mmk_�6�4?N}��(�mP���Kesu�?H����x��/�m~���H[@�M8Z�2^���Jc>�x��̿�=�{��5_��������"��k0u�[V�^^��<��T�ӑ��뻵T	^�g�VX��*��5]�_�(�r�9H~�1�����XC�ʋ�7U�8�S�WVR�D#4��^S��F`",��D�����֎~>��@)��ɑ}w�����s�!�t�;B,/%����%��h �`M�TYH9��:<:X	�6r�\U��r<=v)x���dʣ� Mx]㻷ǞU��n/�
A e]���|F��M�x�q�s���c��YN��#�#��#��	�z F n�$��l�A��*gQ�y&AETc��w�1Q��� v��㜯@Zg�d���p:����J~�yPD�ړ$��*`bnnn��=�2�]��Ck�<�l�a����}�,̊f�7�p�kU�R͕��h�d���.ύ��6��>�OǛp���<�$q5��@���A��!��L� � �U��TTf�avJ��x�(hR:�y#�1��)���יġY�%%݇5� ����a&	,����}������~"y�t;�y'��,�z��3���~�5�rM8��eEg66$���E�j����3~-/�[� T`9+k�����p�!Ȟh����&t��K�z����c]�c׸���bf0�:�������W�r�Iy��n��3 �����l$�1��%�c��N���cMFaMм�iP���Z��כ�"s�1&2�DO����YBP��s�E^>7 �M>W�w�ڬԂ��r�q�u8�	�R�RZb>�$���8����u����D�79Wz�>9��Eצ"�~8\�b`9>�n�U�e�(�d�n�����
��w�'O�rM���1�2�X?�M�n i�I��|�\�>�܃�kXU��0��hs�!�#����	��-�O��;;�;�x������[ê���Za�>�]�ᕩ" >�YbO���D@�T���d�������� Lc��#d�w�G��r�P!�A�p�O%
���k*(1^�<�I.#k:��;Q�zրr�<֥s����n2��Tr��Er5�B����UAD�9���O�?����CXl�hUUTq`��sƦGN��Ȧ4�#���y��#?,}�)�gk�(�"����-**諸�1ў*�~!���
U2x�}��Q48�'b��yQ�Q}���`f�l9g�|��
�Hu�ƫ2��A���@U�߫AdTR��ɍ׫�D��sT����z�C�y$�������y��h1����e������$���&aq�-��� �f��M%u8�?w�D��ב����Bx��Ų���_�)�����mmk߈� [��ֶ���e���2D o��W�|ⅽ�E��I"2�;�ӵ*���5�5 Pi�x5������@�%/b.�ǋ"�����z���
럭ޟ�Kw'� +��rև�~��� [�#���z�4��^U�K:��V�/V2�/����41l��C�Pl�֟أJԴR��bP(Y0�[W�c"�$cJ��:w�P��OZ1 �o��� 
�EG!?h��X)w,�t�n�FU}���F�rT8n2pG�<�A�<�1��h��G��㣏��_��(ܹ{'�o���Ǐ	��W�t�AL��q��}|�OC�9߆#��W����ݻ���F�/��;�7P��:U������u{����gv��H�r�?��R�!|���ɓ�TAk�w���|����L��z��E������ ���۲�DI�9ou�oL�EK�֬����~�}s2@A��6��O Ǩ��� ���<����mX�yP������|LA������6��>������? �LA;lcEpS^� cS$�� ���浈��sQ{�XO�GiV%���p�R	��v{��D��jnY\�B�2��<��A���M8x��.�6��zLq�%L���?�gOnK�>�|y�'�+�(�CVA^�������
�P-�Z-���2����&��)����Ć2WB���Q���j�q���9��}Tٛ��WV35%^:N�zb�|	)Ap}D0����GӪ��"=%�&l���0��!�C����i'ż����*%@],g�����`sv��A�G��𢊣35F���@9��z���Ƃ����K�^���<�e�Ss�����k@§a?={�T$h��n�F{����_�u����N^}e?�aM���Q�Ԛ
�_��1/�b��]x\?�'��ek�e�&�A��m%"�P���`�o۔�q����!0�-�� ���cLˑ	6�ڎk7���y�2����
�DR�Bc0G(kw��-2;ܚ�kp���=�SS��B.H�w{HWt #�u�L;���R,�� ������C�2[Q�ݼ��DH�du-�� �V���eAi�)%�K:*Sq�3Vl-B���e,�N`�KM4k��®&�3Uz����TAE)�}��r�%�wl͋R�(�d�!�r0���Z�X��Ҳ^:��]\�*=��n�|���������|n�e�)Ch>:b۸{�Ey{n�̏~\�Z�B##nc���Dv��J��D{0�)F>s7��#{8S>%+�]+<W4���='�j�Cf�9��z��d%TƆ���l.׶
K����D�Ui.��b�!�{��ěg*py�ዛ�ck[����i���mmk[��7UO6�t>�\?�$�0R^�L[6-(F��0s	�H�P_ �P|��~ŗS�ѳ;����� � ���ռ2m4_zVҭ��R.~N�=~�X�/ ԋ�AAf2P��>Ҳ��/or�B��1����F\�?������%�FN�EU�E��myFH��&���y!��\PY�.K�H�}T�(�1Z����n�fF�&w�f�1�eW�Ix�Wh�E)/ɏѬ�@v�_��{w��dK&�e��P]����!<��Bx��wÏ�~x��G�����w��]��?<�w�+]J��'�
�nw�����g�=y>����,�������/��^y� :�����ն�*���.tUS���/���Y5<��V# ���<���L �{�������.����_���X��1�a�R�^�1��f R��`�+���|�����C'�����ܻKR�ٳg�����ގs�%�u{{�}]_본�77G~�ue��Џ��x>���R����<�?����>����ͮ�&�&�R���r�ߗ(N���Iz��߽{/ܹs��:��1>����޻��?y�Ď%�����!�9�p�y\__B5��~���v	�t�| 
���6�V����(�X��{"����E�g�'*�t�2sK�O�[�C�x�P�KK�d �w;T �ni"�N���� $��׼�s!`�YA���KM���^�eF�2�`/$ }

-�!π�gL��~0멉�9����c@t�KߩX���A��+*�Hҡ���V�N0�5�X�w�}��:�`y��� ��V]$�e�|��O$��y�5����d��t�b[�a8Ҧom'TB�K����T- 'Q�M%~f-Fڈ�}�1���Iv~n��Ԥ*"�t�XA������H\c���{��>L���ʔ~X�Z���3�f���}o���$d4�K�J{o�����rl��E 5]��g���~^Ϯ�ޫ�d���q�V�
��HcQT7ϸ/g{Xb�>M�K���5�e؃p������_�m��b� r[7�%�D�be����S/<x�D9����'�I^�F�2����OmQ�y�S�j]�v��̅�,�*���φ��n�����+>j�1R��yL�*�ΌR��`?�u���,�kX�A��������p���vs�4��^m�p�m�IDHIe�X�vR�N*�}]��~��eU�.:'��a4n����?s�+먈���R�zJ�)ؙ�4�%��
��&M��1aM��u늞3��\�9.%�U��J�
�6UN!�o���}_��� �B�$�g(|h��9�B�;�Eu��?/�:��,�@�{*]��j��㟪G�3�)�k�e�����mW�i��L"7�\��.�L<>{�D����3�p�gW�{�
)��L�zP�R^4%2��jv�Z��<�6����k+����Z�׭�E����mmk߬� [��ֶ���U#8m/4x����-^�P%�Ԫ��,P<)��qo��]C��d)$����oW5�R�
P�6����E�JX)
�E���˗%&#��.!��P��1����
�\Ua�8���(�<Iԑ���<g�U֣E�R�P�S�� <7I[˛?��[�1{���`]@
��R�!"���c8��[ʎ�?[��om�n�
%���	��"/��ꅺa�:�\[���jȀ���WK�D�$@�d������;����/���?o��Vx��Qx���P	���O>�$��� ����W�K/?d���~�<������$@� �����p��0���s��Ww�x�ߩ�W�o��$�ƈ�j�K�\�J���a������:��qp�a��T�h�H\��ԟylo��V�˿������ �d�xJFw�t сsap0[��?ǜ�j?���C"�� C����	J+������7���?�����)<~�X
�^`!>󓟼~���`�����c��AV�����1�|Q��|����Ͽ�1�}��G�Ϟ��v��ᔷ����>��	��W�Lb��>���o§���!_�/ç�~����,��i��kQ����dPg���U� x`�sK���p�W^}-� "����&���O?�ǩ�(�p-A�} )�_�A�Ѭ�T-`s��yIh���>ꘐ[��R�`���Sϵ����D[��-}�Y_Me��SW�&YBI�� 0���N��� k����:�B �6������h�f$,�a�h�={�|��d�e�R/��wدP�1|�����Ƚ��]ޘ�2{���\���7TA��P�Q�F(��ܻ�����c�92V�ݹG��;O��pm�9vu�<��c���Q�!�qt�����]űB�V��Ę�٪\+�Œi�
q�r`?-a��l�F��$k�{y���	�$�k�k��<�_|��|��p����Ӽ�LC��5ss��O� �) ��7vO�W"Tiه�o�?ͣ�9�]����1UڣW_	?������_7O��_��F>�{�z, ��L��9�[ú�yU���<��X�-�)���#K_��VE}e��0ٵ0�N�|��r"x��)�����3��s��R����F���(t�ߟ�)�����7��x#�TB��`Y�넇�'# ���R,����3M�2��3�q����@���{f�c��&k˳�¾d�Ԧ�re)Z�J"+0�A8L�G��HD)��;�6�l�>O��}>W��1�r x@:F�� B<�@�:ܒ��\M鈱�RC�G��k킲\�%Mm+�R�R�_P!a}VϦn��V!�_�W�Y�O�,�̞aao�3&�:�A�l�� ��6��1W�N
�֬�b-���w<�c}}��Y�ZX�P�9ۭ��Q��1C;]��_>�=�<v����mmk�ܶ [��ֶ���]��74�H��������̲t;M��qg�5z7U��3_l����eU�x��Kqcv)���/��l��c�^r�Z%q�V**.VJ����#sF���ת�C�J=1A��D(~7�Ra���N˦�z�"mH�?BX�a�sN踢��b����@q���X.9ɰ�r���>�S�;m`%8��oUo�vm[H/ �����<��8vz�mRP|����=�U�Y����AQ!"(&;`�-�D� &�����a��ڮ:|��@����߅7�x�l�T�~}�n8\�!��.\]$\ݽb�4�����q{s^�� :h9�H��u�nk�Ȟd���P�I63A�<����y�%G�숶�P���^x!���+� B>��3~��rD�0�r����/��8h���|'����yx�wH��
$a=3� �;����bJ�n#	G0�|��89@iU7�0��{���]V[��ǂ��W_}���_|�E������}����W�W��^~�a�O�G����-Am���@53�B��C�����/��5	$H,��D��1������8&>|�Г/?�}�<���)|����g?�Y���|D����Y��{��9K;�D��:xۈT�xCu:�Ů�*��b�V�O^z�%�� _s���c����ۏ>}���${@�旿���W��9����'�t{d��Y�M~�7[�s�*��¨�hJ�J�d�V��TgX��\��q�t���:�B�����Ǜ����g��
Gi3�T_$e�B �Uj����+ �Ң���5n�jF�c!9��fƀy�,V%��k��a�ѹ�e��+]�R���^� a���/Z��T��X5O�>f�$��[i=�Ah�}�۝)i�_3s��!�3ż�^߽Λ�	�u]���[�����'_~�=y�׫��՗_�}�_|�e���O	L����^^�@T��'���6|��l"���s*("ff������z�@����Z!� ���r�$Y���ܪf���]��*uW�D����$p�����oq�c޽���yݽC���O��y᥇��]�ÇZ?�$|�٧$�������; � ���NƑ�L�Z�(�d���	7����	��o��o�k��F���7�$�����?�y�sym�"��(��߱�Wc��i�"����<�hV��7�\��֟�D�3���I���ߑ5���k#��<��̖L
>@-�
���y�£��?���������u�ڇ�?�4������߇_����R?!g��11��b*�B �q�h-瑓��'m�5I�q�E/z��jr�ddҼ�z�b�����2���R�J���C,vv ��I׶.�c���38��5%�$-�I�]C�����
��:����^�{�Z���,b#Z^���7�T����|.�c���Yw�l��e� ��R\TCTZ��6�J+S��$զX����3�L5c4���Lg�~��ccd���f��k���m"J#��*hjY0"BY$8	�^d���}�׼���� ��ֶ��ov���mmk[��צSO��;���޽��E7�4  ��IDATk�a,�j��+��vRU䗤C���_`=�`V $ Xb�E�%�X� �`o��㱗b��y�߇�w���jQ9WM��<�]�7��Z��4�}p��,����L��~H	�"1��t�z8/R2<��'�W,C_3ϭ��Fm	�_�(ȥ��w2�xS~ |J#?3k���dy�-���%V�>�,n�qq��Dv��a�i�_ĨmnD ��T%�PoZU����BիlU |3�U�x�G��X^�5^�_(!�( `���[o��_z��vP ��E: <�bc
7���Z��M�Y��(E(1 r��@k�s�@u�C֋lB�JS���I��h���\
(��ڌ�����7��ſ�˿��ϞY�k�0X������*���o����^����o�����	�)�y��܊m�?Ng�c%?>s���弒U�ʯ�v�j{�C�q�fV �����~��̿�ۿrۨ(}p�>�������s��ǖӱ�$&y�޽w��~=��bU5�x�`����)@+��i�lV�C�:Ud߽�0ܹ�"���?|PE�?��?�>��d�͕[O�^�ގ���p6��|Yk�
Ȏ������x�M�+ٱAY�c�y��Y*�Y��2��{�~�
�>�}�#@��i���>��s�8C���O�0�K�'Һ���]k�t�=bU����0��Ax��G᥇�pL"�s ��/����J���3V�����<@H�] �ooNy�4�@�.�W����	�t�e�a�u��3���mh3�����70�2/ ä��'��B���!M�*�9)e�l��Tܭ�����JW�̞�I�cp��%�	��H�n���+�<����H|a�����ﾝׁ>��<n�!�U��u��c�����?�$��>�����ׇ�1��7��Q��}��O>���D��dև��v$
G�@���D���'�q0'D�Ѿ� �D͕�d��/�܄�<�A�ݻ��0,�>�z���}/��WËym��lw�*XFA
���$݆<�0Ab~���O����_�<��Od�y���Krd����2P���q�w] ���#s�Pbmx�78�q��2��c�$H>��AVE�Z�"����+l��`�s����=����g����iUlؘiű&U�{5/�Qs0W�qN�Ĭ�no���p���7�	?��O�_��_�w���a�G^}�����,�����o���U�
}��b� ��4��I�f����2�p�̜b�4e���(K�ʲ���s��u#�1Yi-
��	��`���F�
�Bx�4B?�usҵ
AR��_��=�r����X�R��Ϙ"b��r�<��6p�&��5��Ͼ��N�|��/F��x��M������=�
��'��R�-̸6���3'
`�x�t��u��|�x���&���-��)1¬A��u�X5�ȟ%�X���Y���TP�����Q��ݜ�p�����g�Ⴧak[��ֶ��l���mmk[��5X ��k�����:�0������A^�#+��� /��!Bi��\V��p�Wꏉ� F����22��I�P�����E�;QH� �h꽅����Pu|<�h�B]9�o
~����h�Q�Wb?�II�E��\���{����mK>2������9�C�a
�����UƇ�]9��u��Pa��w��Z�X��83�th�e��o��=ZLQ�`룈�z�$�E�,��)�pJ�@ �2 9 ����j�f�\��ںTN4�����0���� �hk2�t�g&A�D@Ǟ���V�~l�^�i	�d&¸ؿi?��f�j����hg]/�����q �G�� �0�k�@���^�ۿ�����0�����v����nnA�y�-�/n��c���w8��ئx�K)�35Ne�a�,�� +|g� �����_|)\_��}�e@���£G�
������Ϗ]��ʏZl@��`�,�%+��)��v-�[dk�T5�Z05 &���!��J{����ݰ�_�_x)����{��oK[�d !�����,����܆�&���������?�G�t��>`��3>�;����(��c�����+�=bu������G�{���O���������iBj��̓��Gx�@�B���������-���������{��y���[�z�6] 롒�wu�w�^�����/»�}�`�؋ A�>T4���o��'O�0�9N	���yT�ت���2R5I>1�9YU�l6T����k�K�ɱ��w�$4��[��f)ßY��~ߊ��t���|��a;i�h�L��@FйhrX�@�q�s����^~�$�~���ʣG�Ӧi,�g���)<<���|����T/��Jx��7���Lb9�[����w�
�g7��8�<��w�_����_�<|����xK�Wgb�q!!p޴6�Jn�P;�9��m�p���_�-�)pl��^X�`w��]�9�}~8��1?'�hA쵀n(��{d9����F����M;÷�z#|����|�G�_~��	���,8�5����:	�y�P�@{Ǘ�~�����]���O�%���ZǸ>P�]ݹ����Ir�ހy �^,�H�ӞN��u=��ϒ5��y����XH����u�k��J`:�"�����L*�����s����'�ڣ�uȵEcµ����O��S�ʄv�Q��Qc9T���|��
��hX����� �xk��
�X,���m�����$,a�x�/�xW�`����W����_%���A��,�b�I���px,�)U���2iM�'��6W���E��:J}a}H�����bI����Ҕ��4~Gݧ[�pH�*��8�M$r6��.��V�+P�Q�.�p��ق�u��3�(�)�j>�D7D�u����1�qn�ev{~_�]��I�R�k{�j�?�p�Ϣ��n��W^y=��wl�ֶ���}��F�lmk[��־V�}^ݘTո�vaR�9����Ӊ�B�6�b;x�[��m��5�SUNz�E�c�_;�$U�7U"?F�;�Z���PTj ��?�Cm�L,U����J8{��Gl#��}�H� UѰ"�ϡ*�m���C ��L-�.��R4��-�H_�`��6����Z^�k˳��;`J�/�+ �XX�?�K�ަ�j��UO�)�i�� ���y�k��_z#��r�qeمl�D�I)��<n�C	��GGg�F�3��14�!�u>Ң�$��e�6���W� ��귩k1e�Hu�c�K���P-�d�E\,<f� ��}��[���]C�ڙD](�LeU� �  jv��1�H��g�)ܹ��m�K@8��!Q�p�8*���w������_���|� ��t{q�
� j�js���u0��8�U�xaD]Y��FWE����0�ͺ�\�uX�3�!�o �������a�qpss�ㄍֆ��y�{)pUT�(˧j<���&&��	6H�s1sC}@b�bZ�-�d���)�H��#7���˯�"����b:@�H�V��9_+�U�d����Z��ڇ/�L�����]x뭷��@e��E`�5�3�3�~�RQ��Om;�l�����w�½�Ls}�1AU�X�����h6�]8NA���nM-'7U߻� ������~��_�7��6ɚ���0����w�O����/��w����eC2䭷������$B`%���Ixq�k��J��x��y.�0'�)p�+�q��U���U��������1B$��&��BC ���1���x��鍨),��<)�<����D��v�'B���+���-��P �����;�|;��Ǖ�c\�ZVe]{�����y�X�z�r���s&�T��s7\ݻk�ן'���x�ƛ��K��1������Ex���nʙ`��Z��N�6�����@����;��u���{���}���pqe���|}nO}xzs,�1�sɯiE��`s�!�������5�ʗ���ߨ����Yy?徺��d��$@����vy�PD����B�����eQ3�w�{?��p��<�����?�g*�X9�9��jSAⰣ@���H�}=VS�����r �R�T�̒��?�'Q�R�ǂ$�x���{�.9�,I�����Ҩ�� 	�@P�����y���9��L�n��	EZ
(�2�s�{="����	�� �����av�K"2|ܾ�]�����{~ �N�Bb�%�2b|�:ڗ���|^����/C�K�q���PRK�56g��ڛAU��o�~���"p�~[�yk(�j'b^t�=�c�ͩ�T�:��d�n0&A`����8d&?Vʐ��i���ʧ��Z2}�>�k8���T�+�t|����ڨ�1�=)Iq���G<ڗ������^��S�s=�<+�N�D�����^h?�i�E�G�$T+�� �Y�����O`E��1�!{���s	J9ڦ���^����WҀ|B�Qe���ʽ_�u9(K*C|SE;���Ў��,]��yR�ޑxV ш��y�oݥU���翼Ӧ5�iMk����!@�ִ�5�i���@[�?�"��b�JLXR���t�U� �ےXy�`X��y��ш�Z5F�$TS�����i�:^��RK���EjA@�܀}��|X4A���M�HRL�!.�b�r@h��@���=�X݉<��hL�	�ܮ|��A���P_f,�^L����:1��K�ꢲ��,�,�H�����UyN7�a"���(���ՍJB�aȥuH-H�)֧�KU~����!�J8������a�82�I�2 �c�{hl:��'$W&Z&�2�y+Q���e��6i�%4�!z�[E��������ۙu��+�@P$g2��P���r5���Ҿ��9�^U=�H�����Yu�j�^����:�B R��IMAC{�(�����bOh����;`wt��]V�����lgKs���'������K�?�,Xe��y�?�Z}B{8B��}��$0�����@o�Uծ��=1�,غ��� T��U�fwk������4�c^lnʃǏ	�&��{��ܦ�R�7'ۻ[�W e}X�W����y1��H9-��ջ��|����0B36��d+�K���ݿ�z�]��Q�.��<�­{;X����/�vWÁ����Ǽ֯�;+�;���eiiٝ��;��A���՚�|�j܂�;���/�j�|�z�f���c1V��y�����#33s�a�
���Pm�����?�{إ��rcJ�#G����K@��(s�y������=��	Hzi_�\�w*p �����q!��܂9yJn\�.ׯ_cV*�;m%�0�*T���p���r^�u70[oa>�Q���; נ��ߓ��������D� g+iW6< I��~"TjAq�x��U�R��]���G����% ?r�>�$ �}�y��7� ����曝�Q�0���,��� �y�G���Dv�!@^�#�gB�NJ¬�kS5��3��*��K��d��w��֍�r��m�{���?@J7^�^��noo�v����BZTl���;C�i��6N ۠u�s��Yy�W���S����Y��;>(>����4���x�\N+Җ�p���;���euu�[wt���/��O��_�*������@�eUAUJ����a*]7gi���[Xt�����tb����NܑG�;��u����7����%K�˒��j�
��dLad��lgH�Iܦ@�xuG>I��x�K˚P=Uߑ(���$��2��$�/"����'�}�Sy������5�e<״�5p�4�ܘ���3�\��ʃ�*�$}�{)�p������I�"�K$!��=:+
��3 ,H���*�ٹ3���ü�������a�Bl�_����M-���A�{['��cFI��%O��:$�mH�8��$��VIUq^�T�Ю̊1_X�X��0 �����C������-/�m� n�*�R�v<J��e	�=�f�y
���c��j������I:,>�u`�X�{cbDq��KB�C�K��R:q���j����6A�2���Q�5���j7�5�9��1�K��-�:�#��,*�� ��|�[�{�y����w����Ҵ�5�iM�� iZӚִ���Z�^N
����I�/~b@����
�r.	>
�V��a�����)��Ee��`��`*[��U���_I�Օ��R�/���wݷ��J=QT*�i��L����%~��B�!C��"�ê��bj�S̓�ަJ��RD7�+r룉�]�AEo�k�@� ��(����&,4�#����\�^�O��Q�7�g�>h�}Y�:+���G�����
7nƹ�lþ��Y(�Y%�$�Fn'���+��״�EY%���U�8W�<�R��; n�98~�{ۻ;�;rC�e ���]G��?t`��~����,���rdɳg��ƙ�����}����ޕ��M�1ș�	��`�xGv�7�+��իWe��s��+�}ey߲��ƛ��ۗ���$,H୏ j�Q��0�`�R�ld*;cU�1��Y�Z�P呙��P��\Zm�
� �RF���u���ܝ���S�3+.�������y��q%)t{�+Z��Ҋ��?�UYQgG�q��k���� V�`���q"w�U�Ǭ�?v��|�����768V�����uW��� A�֧7^]����C�9��Q���[7C��n��H�!�cX盔f)c�k�6��K7f�nB�33+�μ���ﲺ�L`*'ZY�k�+!���L !�����8ݷ�*�O��O?�Dμv���`Or%����%������}�Ee��YQ;���%y��b>v서8yR���?��{�	�)�| u��c��.T0���׊hl�Y8z?R�3�*�,L��~�DJ�7��
�.HBh�@D�h8���ۿ�L���Y��c����vDf��sd��\�xQ>��9u������@_c��uk�ZD�\�E��T���.�T��LK�[(1� -+��P�(�K�! �Y9z�#��yy�s$A���[��/�[�p (0�}�ƿ�Å�}�7?@
���H�D�2d�{o�'o\xC��<��>[�ܶ��TI�0P%H�`rZ�o�(��l��`R�[��h�{i����̺k%��&�����w��7�����.¡��ĸpkZ�$\�BS�A!�t���4H�ܝ3r�p� 
���w]�ﱛ��nM�}��P�@�`V
X"���0�2<H��~0�_��,#��=ƹ�.,��[���L��[�Q����?������7��=B� q@�2��e��|Z�Z��Af]mі0&�FEw�ÿU�5r��	�W���I|���B��Y�w���� �:5�Q�Y��gs%M��,b�?`|�:N�����݂DN��#��)0�?c���d�U�u!���B�U���>�|�¬�@�x�?�z|�qОV��K��qYh9�\o�;̇)��M��y�����ȲJ@*�����T1���t}*B֌�Y��TYgPn��ڼa��sf�
ހ
>��X��Ȟł깂!��2��
0h���9[n>---Hg�G�ִ�5�i��� MkZӚִ_W��Q \(]�S
��C+���80uѪL�1���Ӽ�/`�'+���&�"�	�Ef���I UG���{A,&�&ڵL�r��tW���
���U�K�Ww�ԧ�j��i���m#��kT�O҉Z d���5B�����Re�ض=�@�G�k�Q��0�NL��}C����S��h�\�_ qj��[��3F�h\�|�[�ǰӯlv� ��B��F\űY�5�25�#Ki�{[���"!�4}AWO�\�l�"rh��:a���&P%�������`v��q���%���b
��?�eyyY�:LP��N:m9|�0? ���G���K��
�1z��9?ulq��� l���wo��������*!P%���A�CT�we߾~�m�vm��	+n�G
T'oml���]�Ndqq����ɜq*ss$h@���
ǎ�3��	 ���U�}5I�2�]ޅ�%�u���|�*���M�w���C�q!��͋ !@E���*A5=�+�r,8��5h�թP�7V+T.O��54�U��j�B�],��J0���*�ϼ(h�3;7+gϝc�;�-vv�����[�`������1����~ '��q?s� 3��
��h�����G
r1V0Q�VJ�V1�n��25AZ\�'|���[\f���l���c��V5e��HB�����%��vV>��'�0� i(S�lDP���T}���L����"Ukўɬ�@�<��"!�uwk[���͋��-���a+�8�P-��M�����V�/6P�\e���f��+44����B�HU�*��չE��2��&!�A�~5ȭʯT���5�ȡ#r��[����˹s���q�1�(�`��2(��k�L3A�:s��&mq%F��>��P��PD�<��p���EL�7���[c����B��q���n?�1B����r�1���hq���
 T�9vT�}�=��Ïh{ŰnQ��+ݨ������ϒ�'�EQ˃1�>�X�1%�P���0^0oݡ;v��{��I�}�'���������
��\a�%'�5-}��b�[����rX7@��vϭ��Rﶻ��mϰ���7ݺZP������*+��H��=��4+}PkD�����~�������[����''O���?��]��e��f5��iE���a�fe���g�����ʋ���v7�YXqMX�X.y�x]c���C��ӳ�gO�Y_�����Z&�"UY��T��|Y�FD�Tc�b=ɡX-}�������"+�Ȟ�r��s��@t*E���avXR��(�s�>��f	��8�s���PC�Ӊ��/��ȃ�u���q���J���P�!��*S}ކB�b#Т����q��^�7�W%�ܳpWA��oaE5��)�R=Smw��@�g��l.����
Z���`���4��kZ
�O� }ƾ�@�+��q��ydI��!ȏ�`�>�~�4�iMkZ�~{�!@�ִ�5�i��1� edk%m�'pb��,5���G���hE��M-��Z���jI�ʬU���$��FC�W� ���k�ޜ��\AO�X�wZM�2ib C��_U���e�V��ZxEH�KJ�����W��vQ��r�B��!^\=�a������RAnE\��? :�Z9b_="j�UL��ԾLzL��K��+���m�<�Q�9�4 :�	��6Xf������Q�B_��Jo��^j�v����s�9!�t����kE�-kp� x�#׮^������0#������c�Zv�~���P=�����9�)BHy@`v*s�s|�G%�`0�v�-�n�bU? ���-V���9	8��p̟1#�7k� G���302 ��NP��(8��|���e o���|���PTf���;��<|t_~��\������[Y���9*S@� �Z\X������FT8��DQ�CI[&#�n �0��G��V��~��>�n�����`,w��b 5��>�!�\��*�j�lo�0�A�s�W����v��G;3�(Rڞ�<��f^�H�s[^X��?��`���₩r�����~�<oD�%��s
�6LG��'�w�u��� ���3�V��^,$�����(�{kk��
�mav^I���"5�W��lɃ��ޫ��K�Z(>���~���mr�]ZƩ�
�`r�3p��
 MX ?uB.�}I.����+w4��P�ֲ`<8��1�w�`��>�-M� ܂�)�w���� ��9�i/֟�RD���B#�< ˕�R�i%�gD}>�nS{��Q����K�k U�rLл7RQ0�a��ܘo�P>V��-�@&�;{V.]��ker����뼙 �U��mk��
qpH�V�o�9��X��f{�$ �V
�Q�L1$vy`�A$�\�ݕ�Օ�U� ��l��/s���R�yJ��$(�b
�[B���y	�dż��$z ��/���`�9W~��\��ƹ�%|v �9��J��y�� �S,߅�����)�n� \�ܹs��h%�wk� ��HW�<�Y��+�#��@��gO�T��!� �� ����������c>㴱�p��&������A�����
LU��я��l%�r%��C%�{3=^�ݍ��g^��?�H�8^��9�ʠB�,�@����*:�ǖ��hee�k|�i_�jk�8�܇d�����@a
,���1S��{Y}���d�և�c^���#/�yNF�c�u�k���i$/`�cS+,U�����A�'��U6�s�%���RJPa�c��I�!� ؋�z\� ��bn�"���L����G1E���V.�j[ӭ����j�ZF�@���jh�[f���H��ᜊ���37-l���P�i%$!��(*�P`Ъ�S]g�R�EYl�cR)Vr�@~压�VQg�$�.I^]���xܚB�9^\k��rr`���_����4�iMkZ�~{�!@�ִ�5�i��F�j�ʇWs�*	:F�ZH(H�C�cV�j����e����v�KU�m� ��m�1(�0��?|ї+�.����瀨�CM�s��/��_:���^đEj��&������-���|�:���y��½���>hU{�A�ͩo��a�mTY�@�m�X�^./��٢&K~��J��[�YM��4��l�; "�aۢ�o}��EE��a��yl鰳���`�.Ͻ_��<8a��,�k��jC�@�f�f��f�����gkr��e��_�(���S�@1��O4иT��9���? �jݑI�} ee�ྷ�P!RN�l���G��j�:�4��g�<^ັ�mwh�A!��x��;���+�A~�`�j�|�������r��������Uy����ڿ��4�P��(�����6��hoY��sj���j���2��z�=u�2�$I�
���d0��
�"EZ��y�����;H�k�/_�Fv�� �����vhҊ5�*����Y�`�fݸ���jʵD������%q���O�>B;�ޜJ���ʩ.��m��r[�<��7870�ñ�@��6�\ �}�;9~�Z���*�����e� x���]�����c��>����?(gN�fH���� �bc���< �Ȱ���y��X�;c% ��ae�T���W_}E�~�]9�j$����k0��ǁ�]Qo{*��D�w|!��V������k��"�u��^�u������ύ��_����4V)��:͖�m�J�z�h���S�-jJ����0�
�b>�*D �� ���5��}��q ���ʧ�c_ھ?3"sr��1��O�⥷���W,���։\��� @$A��ɘs�?P��;w��ݻw����ʢ���|��0�9_����L�@`}�_Z�w�}W"���ꫯem�	��E�c���LeW�x 6O�V��ۿ"�}�|���ѣGy<�fx.hqʨ����^�rݙY*G@���������E ��Ь�p|���<��Z+|ص�/(��},.��w��6 �޿{[v�:1��e��-wVE@�OxM��n�aɵ�gq<Z��/������WV�[��_ʋ�5��#�_������3%#x�/�92Ϧ��G�cg��U�/( H���$vc�|�o���,��Q�U�L�����x�5YK<�oyu�z��?�%���0՗j��9��%Uy�@8�K���y���;)MmA˦L�9PV�F�x;0�^z?��1o��"�m.����>��~{���t#U��S�1����z~aL����dl�WظI��B"%R�����fՊ�*��d$����Ș�N~��3�`Ov0W�l�
�2�Ͱ���"�(��1�>S�@�o�` �|�0#ur��5H>o�囒LvmhY�ن�s������[��#7F�c��X3��lm8RkN�l�;ܑ�5�iMk�o�5HӚִ�5�W�$-�i��u/<�?��)�*�`���l������p�F�@�C��l������*h!QU�U���Ds2e�W5�j���ma�1�寂�_n/���3VUgʔ�>�~Ȧ��{��jۿD]��NMN��Ϗ$�*Xuw�����Ϻ�R������-�*��qͳ�%<�s��I��q˾��`���SU����p��v��t+���x�&�`c���V�&�*�|E�o�!������>�J U���s�S�3��l�, /��*E"T��,'}ֳ\Ǟ{T��u�]�b'��< d@05�2��w\�ĮUЮh��~��j��/��������W_��_}+��!�;�$�(�����Ĺ���>0�\�B�k �+P�2Y��K}Ĳ>h���e���rנ=�!�G2be�X���(c} �4�0C[1("h�<[;�_[ۛr��5��_��>
)�9Ns�@kY8lHr��V�N�Y�)P���0�`��F�rd%	�sg��G}$o^8O�	�����c�a���]ߣ���Xz�e���!M+���W�ʑ#�,�D�\�9���6h�e���������A�;�ׇW�?L� �k��ɩӧean����9%��F��������S����$�`��ͮN�?�S?�UοuQ�~�=9��(Y�Z�w\�&��w����T� �c`i~I�% c7�,�|,4xiq���?�1	�� ��wg��哉����oMU��>���ZQ�f9SP�!��WU��z�kت�Na��[I�\M�vZ���=��nla���63@4;#e8ȣ�/����ü�̢p�ݴU	;\iI�����$سg�tm�*2v�_��Od}��L(�`��� ����Ȳ�s��ٷ�$]�w-�%����y������������dKIK��L ��5(�I3���k��V��� z�-9~�8Ƿ*�d���	���+6(�Z��,��?\���O�\k�|o�
����Th9xHN�>���՛$Q�6$���N��y�7ȉ�?���z��o�q�s}Փ�`W�fv_�J��H0]Gu�JV$���j�V0X�-�+s����y��Õ�����J�ce�����z�G���ȁ�sV
�x,��p�+7�P�2����r�.\z[=V�C�,�˰{��:��0��ߑ�ڵ�L�h3慷Tc�%Vɭ�����|A�f~	sFJ+����3 u{>���e#v/��a� 	�+,��͂	�i�ؔE$k��z^+��U-�n�sλ4uF�*��d>$gf��/�����b��NZ'�إ4r�U�R�D9���D�k�T�l�r�L۽��{}�,���|���%�R7^(]���}:ۈ�����N�$�R<���p���teu��߃`�G�׮����n��:��`�������vWn\��$��m�N6�}�'aT��c�ݖ���5�iMk�o�5HӚִ�5�W���	{�`P��Q��i��fՓ�'|���a[���JI��O��v1x-_�k$�c_a�Tү =~k�)}��;�'5��9�c��R�IV}�Ea�j��4�"�W�� K�"���2;�ضYd	+רF�+i�}Y�W$�D܇aŁfSV<d�ŏ��Ue�z>c��4���	Ox�$����GƄ����������
\�8��Y�.��O�1תҢ�����b*�$�1�P혚uu+b�����H���`�фY)��tB�4����F+&iaA�^G�2j�aƝ��L��@+�}u$�@��p�-��I��A��R�,�4,�@h�^���q\���;�e��S���,��W1�x�K�s����öf]���, �T޻1����T�Õ;ݶ	ȒL}�s��nn�>��%�E�"d�۷�~�$��( �� ����r ���G���'��� B�o�	P�X�ϸT�T������;�m�vT�f�'�XA�Ny���*��� d����l��q9r�à���oOh�����#(�"� .�An�F�m<ߐ�������7n�h0Rsp�����ɣ����>�{���U�X^={���_�h��/�u��U�p�-y��\�>[gN����:
�����A8�����)N,��vaPLmmmq��= �n�7G�R8q�^O w
��
���	����"m�N�>-;;�n�x���(�I�i23�B�%ܲ�"9�^��#0���� �m���Y�}ob���wc�|n����B���퀸�*}y��w�:�y�H��	���o4q><]{LB�8��ܕ'��h�9��I̸����#�G�|����@�@r8N?��nd$n���|$Odna^.�u������/�����?��Ӷ��z
���ŋ$���g�� ���u�{fM�Ec�]c���@֞�����;r��=�����6��ʑÇ�N��	�s�=�ő�i@�V�J����y��)�^�ڵk���C�]��FTc ���eB�ʍV]l�?A0k�D�s�<��-w=O�9#�^�����ߵup�u/����>��
"�h�*��Z��YQ�m��*�Xi�q�����像>�[��և	ϼ��]��P��ۈV���/�F�[;z?q�6,H�l�q2�-U,pn���Zn�{j�M��q6��C?�
�FƼ�k����X�F�/ƶUfխ�(����K���H�6SW�wp%����gW�P7j�E�MD�V>��yǤʏ��7#�/S���9\_�Z���&�!Yð�B���ݣV�S���BI��(J��ܕ�P��
\�b����s��B��-�13Aẗ́:�ڏ����x?���
[P��@g٘�Pq�Vo���*h*�ڢ*����:��3��*P�y푻�u.1�{P��6�XӚִ��f[��7�iMkZ�~u��Z�J��{�T��"��N�d�Y�V;�řd�J�@0��X	F�!V�+o%�Q`)�}�- y0��@;��^2;�>�`�Y2���J�X�
�D,�W�G��-%$r#*�G�����K*���Y!�2��gQ�2���5����k���ie���R`ЛGY�g�")�q���2;�3�~~NxL��g��jOj^�M
�~A���^Iƪ�P��VH���C�ε��Ei{,�J�B�2�Vf��*D�>Z�=��B�zi��� �2xl Y�mj���o��u���8��IA�3�J�&�5�5
0�1�Z2�EHɠP��m%��E��2�/��ڷ�b
s��ߨGP7��`S�I�@󎁨 ��{�<�1�9<{�T���k�r�;*Ef{3.����H�1�	%$�j�Q$ \�:[�\� ��~�2&,�>��
� �����Hh�J|��laq���A˹�@7����t��:��]AU5�/�f��j[�| C �ܹ `5���Q�ٵ`>���*Z��!X�๏��wW�� D�7|��\7���ϳ�G�?S�3B-���c��1@%u�$��uh���\�|����}G��~�T�ggf��IǹG}����&����B�"��9��X�~������]�A_a����	2�I˒�o�R5��O<VT���q1f%�?� �|��ܸq��K��Q���UZn͝�͓z���ĩ�$W��-���b��9�~��Z>zDN�:%7�!��M�2��	u~3(9WK�(V�r
��ª�y��\ҳ�
fV	�^����3�O՚c㎕�$��n�6�j�C5��>C�
�^X} FV���~Z�8y
�����y��f�J���]�ﮯ��O�n�/oݸNb	d��^��ܯC�K�U��Y,;�۲?�
�=;;#���H ��믓�b�'>��Ĝ�$l�����o�f��ۛ[$R��M^�p�*�]�+�Oȥwޖ�/r,�{���
�|�� I���޾}KܻCE,�>x(�>!yE�j�#Z���L�|�6�O�>�;��CGr<a��X�N�?�g��y#$��K����*G���7;�"s�]����XK�ꌵ�?r/�B��4ː��:n�i3� ��ʐ�c����f�簶loo��Ʌ�	`q7n���g�~Y��#�JS�	Tz��; �1.Ǹϕ��s��1��w��'���d�yU���Z������);F�*6ݵy��1�Հ$;�m-�uwǑEj'��22zڼ���	*~�m��C$�������R)0�)b��;��J��瀮���	��M�P����m���+7���P�:���#ګ��q����G��۹Yx=2::�><B�)Y����s���Ǫx��
˷b�y�y��Ȟu̺K|ѐI٦�����g�I����S�~p����lꙮ����:AU!�Oy~.���!���]b�ϔωxn��4X���M��(���D����a�KP�3�G�6�pU�z��s��ӧ�=�'MkZӚִ�^k��5�iMkگ�`��M73x)�eɿ��2Β���<�K_�-p����<��ږl{"VD����TV&�T��7�y�T`H�YA�Q3_ʐ/�?��v�-�;��"`8���I��Lafɑ �;<�{��<��̆��[Gp5C��E��0GP�zn�y���"���f~d�_��e�Ab@'T!{��z���ߓ���D�Qgu��V���g&��ȫ���a��(��i�/���c�U5o�5��a[DYb�}f����&��7A^yˌ���y�3%:B��Ԡ䄠\D�*��.ͻ����*��[��*]j�ړ�fA�Y�ޭ֊��G��g�xL�D;y��eyU}���A�[I$�����̺sps�}�
��6���" �= F ȍ�}����%���U1���t8��7:m���(��3�&�\���������0��%g4��Q]�r����&������h�UY6��! ZhH03=����uh�2�ƴ!��H"��3�6-j�0����v5�`9��|A�o�������p�� X�ϾH}�#�I�:;���"�L
|g��%�Uݘy[*����
K�|��g� 5p1`5���͵��%�gd0* ��&!I�����ڥ�,--p7;;c�	�������aڽ�9�o�f�d'�c2!H��Ǐ�_�Ӎ�Yy띷	��n]�u���<s �/,,�Ç��z�2;�����o�Ȏ=&gΜ�����w?�P�q��;�+�w�m�������ٳg��AFeW�֛�R֋g\3_ll�m���}�\z�*�0>%֠��Lh������W���7+��������Smm����Ü��EY(@��A��`p �nL紳R�Ġ�ƨ�d�Wu]ȍ��$�W�a<b�zU��`Zq��� �b����|�����r;^1�c���u߇R��?��?�/�����z&�P���KXَa�
'����\(�n��nn���'r���Ih���k��oʁCi{��O�f%���ww9V��r��+�؍*_�q�}�uz2�4=33'}������ɓ���W^s�yY�U�\=���*)��?޺!�_���Or맛��]�mw�̄I,�Н��B��n>A�*�-�w�'Z�>u���]��Q�ǵ$+�V\c �}��_�?����??��lm�p���-E@T�U1�Pn������`���2�����*8UT���?��+��;;[r����ĭ�:f'��'�;�q]u_�5�r�+��BO���#U��!�j�S�n�ͻ9����{y��wI@�&	[���3�Wg:j�Ux�A�,�I�k(^�F�=�͕�ݾ�%�Pra�e&UjA�/x�A-8 �KK3�6��x_s����r����ד��P2^��ٛemWxF`
�{wm�TDi2�0q�u�ڝ���vܸX������3�s���U�g#�Ё�מ��r����*"*�r�B��[��6��D�S��eD�9U�P�P3���Up?u���ݟB�J�bDj��G�9odS�#����yZ�x��vn�f>ә��NI�pM����T�2�*�U����4֋~_	�!:��5�0�>�}�S�M*j[	�V��mZ|��8��cx��δ9.�_�i�d�#�&��,^�ִ�5�i��� MkZӚִ_W˵jO]JjP�eK�ѐKVe5L���y
 ���Pf��V�I"�Za&Eeo$|�����q(,4*](�j�*��bX��z�QUj��vV��3&��Aod����[L�`?��>�R�ߓ�!��}Y�Oz8��0�.�JYS[h����M���^���ڪ��nL���mJ�:�e���x�Llx;�bQ�+�&
d ����WׯB��[:Oĕ-����{W� K[��(�@,�Ğ���XU�U���HΕ<�v4�Z�H�,�Y��Mh��X���ص��`Q�Qd�#b[ƍ�ױ���%m*F|�,�E�Vo na5BH��-#�HT��hۨ-� ���`#�f0 ��1=J��Pc��v��	�J]ZjB@6��02B����D��Y�`��;=H�d��tD"�0gU���Nj>�V��b 	+�'���?T����$�wPXdYV�j� ��!�$ ���Ƅ̾!ˢ?����:	T���J=��d���	r�bU�1�z Ŗ���5�'i��?�r�ܼy�� ���qͻ�Z� ���shw�X�~��m��/����e�`>s�	� ������(c[��I��*�ٓ��$��Α��e%����ښ|�����?�����	z�Ơ6J�i����}��׎�|G��2�0Ϗ���t�0���*�ӯ0��$S�X�S�cj��9"�-��W���i�+���@����_�W4h�����&n=I�9%e5�K��A�ucaqe��y���r��i~�*I�:���q�g߾%����5�����y�?�oVD9���pm��)�J�7��Q�1k-�����ئ�
Z�Vw�E���Çh�D�I�V D|_D!�af���`]����O�yUxv�Y]Y�'N�|�Y������nw� ��G��O��|��g�������&]Z�[!�t.v�21��	3X
��Hz��mݐ���+����8&�iF9 X1nN�>#}�1�$?\��l����=W@q0�*b�{U��b���/f��4�jJ7&�v�9x�|�o��������kin�%�%Rh�6�O+��h+%,�hE�?��	�s�s����w�țo\���E�]����5c�c�5**�Ǽ/�ʍc;*�'c����a���J�t�����KIAL@�#�oo����UB]�������_lʏ<���n�9sl����F�[�ψPi�2�d�j��\ d��ͪB�Y1��[Q��G �W�uTw�տSSh�w�]-��,K��vG�J�� ��g��!��J��|�|�!yD"��C�S�hQ��N}�@�w_{@��Tk�K�"�Iι�E&���y�ܥV�����*�Q%Ml*��c�p�(�G7{��,���CiAb%�m?q�8v�����Ϡ{U7���]xn/��}q��a7��^iZӚִ��6[C�4�iMkZ�~]/�E���W��~�E��B<BU���^4M0:�eI�*��g=�h�����,�kaV��^�*ߔ �E1�(�N�P+a�@���jWk��W�FU��^"A*�����w/��ѠJOt�q�ͣ����T���1��v���8��[��ޕ�x�_���t�TŴ'2�H%8v�9]D��GRU�UV[/���f��V^�AG�)/j����X��ٞ����>� I$*��O
��:*�2��x��W]�g���rC�^��|�b� (� ��_�u �q�:v�b�K��W�n>���IG	%0��#����+�Mg��V���JQF�A%j�3aB�&�C�O�d
<xxWv�7�X+4��.��Pً�T����ʰ[tET���h�[�݅�C��Pj�o�  V)㬰�fV) d� � `��x��R9"dT?�TD�;l�y�
�/ƪ�Ѱ{� ��P[h8{�qΠB�A� (b.��s�V�5�r�j�2���a�����>��*���,�J����1�$Աӛ��W��&�a �kO�������%��[��vJS�2��%�������w�r��7r��S�����;����n�;T�,//1s�/8^d���(WC߿����h��n�7�o�5����y]��HS��Q2W
	��n�P<_&�_�̟/��Q�*�-z0G�_��P ���у{zmHvO{�K56�w�������d�ϊe贪�	�i�+��fQ��*��U�ޞ(P�؝��X��e�����`?p�fK�p02���/��_�&kk�I�C�CP dlĽԹ$��_�=N^7�<|�����ܶ��Z�<�{��[r��!*���6^�&��6� l��'���M(G�2�t�}�o�>��f�ލJ;o����+@�oܖ����Mܿ��K14���~]��H���祻n�n��1��R��賵'����h!6i�0�H���L=��>����Uy��!����<�_�X��{�'o�|�5l�`s�|%���K�M�Z��4��a��ej]7C�	-]?~�ͷ���c���6oX7:��y��qEZ�kY���P���c^=|\.^�$�|�,��J˭1P�Aa�%����u`�J�!;n��p� Rq���5�O���c�k�۹��ZN�ߔLӱ�0O��Y(Y��u�@Ir�4�+��Ic���	�쁟UVV,R�yq�@Y2�=���{�����p$R��̸�37;#������s��G��T�ܶ�u�ӕ:���J+y�JPu\�a�*���1	|��*-�&��b1 Om�B1���ɪ�YO�P����ψ��qqsO^ih�?���%�2���q��b����h��W���z��'�ytL�� P����V���Miڭx���j��k��l���\+]�C#̦�3���%�uh�{x��W��D*ΧiMkZӚ�kҴ�5�iM���Ds8|5�� �i�M�e��K�T%�`��. �VZȴ�RU�WU�����q	���
$6p:��G�3�0 �_d��B�b��aV��/�*�����,g�J�A�>\�J�D1`�M�8މ;|�U��0�+���eQ�q��V>D ��|m�h��އ~oO��T ��^��Ŵ���#)����J���#�<�t�0ʫm2���`���hB!���DfS�T�/�jO����]|�Jooa��� 	��pqZ(e�Zl�B%a�4p	�j��� @��z�`n$L��/�����ɫs���o�1'4�W��G6�b�3d\h�.lT|@r) ZA�eB�%lFE�䪂���;|0�}@8��*��+-�PkX����w������ ����a�
 ~"�z���P3< �3B"TWy������
�}�K��k��HF��6�5�Ȁk�G�@k,�|�cFc qX}Q��Д4�?���m�F i$�,��qX����a��pW�>}����G6+�#f�h������*�(
�1�/�X�S`ׅ��Y2�c��~���I%O[�.�7���>W{Xm`o9�n?�����Zu=xx���<]�TW`���hKBS�%�;���r��U�t���ˁ���u��R%����;~R���G��s{Tɴ�tZ�T��.���q�,���x�Y�:���F%�s�RD�M	�J-�I@�r��Qg�l\�@3C�#���r�x�*�˗�����Ѧ���ph�֙/gϤ�P����v�s�j�D��V��]��)�n=�"��O'�N�P"6�:wwVVV��������ds��,�"�$$,@$;v�dաI�e㉩QԮJ �׾�&���!���sU�1��	@��~�"j�Dtd
f'�r<���ﵚ�ђ�/����K�7'�]�9��� 3v&fŅ�r"K�K���oȷ�~#w�ޮ�_���猒�e�Z���O��@�����XPA1��wk5��<���OX��q}����D�R��2�@���*��G��pΰ�ߥKo���.�9����s=n_���L]_߸q�sJ���e9�ꫬ�G���+|�0��rgr_�0���{�:Tu���^�2����P��t����R@�y� P�D*���\W��%�<�_������`����L%d�P5h@<�#�O��$�넀�15��)7������=���0� ��`m������D���c�5��2�G��� �9k��9�B[�T׌)�kޡ�e��:���D*U��b�u�L0އ�P��J~���d}��`Y��H���0r�@�wa�	�I�R���3�a9Uڪ�d��?��lnm�Z�oyJ(��̤9$�����D���`�]߅�%��"�?A����ߦ5�iMk�o�5HӚִ�5�W� ���`(h�/�Y��Ɗv9_a>� b�0"����Y���Ƕ�p�~�պ��zh�H�jq{CTрmC��A���ˊ�J[Q�`}�M�A�����E�K�OU %Ua�Y���'�׻8ҐVz�
�$fZ�E{�?lbj��+��F�LUO��P�ĈPR��O�����(*�C�YXEdQ�W�I�����P~v��:�XW�NkՍ���� ���b(��Va�V�.�x���Ȥ��9èSZd�V�O�j�P�ᰑYH��/�<
 �U�h�v�H�$60�{�I����Hf�,�5,���1�9�Ҩ�Q�B�	�`�)�H�Ւ�4�l��&湏y��a�z���YJ�nu�~��PGep��#V7�� �� �a�y�9;9(�}���P�F=��
K�Ɉ)�OI"�nmՑ�3ii�9 n���Z�1�G?2Q��
�	���T�X��H�$`�:m��j�U*0%�1%�y)p1�6B�Y�iauo����-ԖY\|���ItX�H+ր\�����kr��	Y�_PE����w�ܑ���o��l�B���L���>S%	T�Tp�`8 (���r}��bK�a�u�U�j_28ݝ[�ד}��$c�q���^3vH�VM �p���֫A���㏷�Ν���bC�&Q�!�a�)�ZqT��!΄�.�����ƵkTI�"
n�@��A	�F��/�=}��m��� �j���6�Ҧ�(�d��aV���m�R������ =䗜>#/^$(��k�J�ʡ��n��W-��;�]n����"�Ir��h�ִ����گE���ޢ�@<��v����2.C� �4�	%�W� @9ߛ�9�>}Zn���,� �2�.PA�q��9���������Y0�؆;}��g�p�}���s�"s��#�;�$�0�0���QU��}P�d��qR���Ύ�x� ����j��㏲��L� �.�l�u��?��vn���U���
*�k����4�Ǉ���@�omm�W_����7e�҂�_]���9�#�,����C^�<U(��o��Fn���$BՕ���z*w�Ў;2�i�s��)@kF���������$�O�p��6� �Q��� �hs��`�_�9�`�8����Q�xO�5����K;.�%��Ŝv�H�I��d��-X��"V�c��[8�� �#���-��C>+�`vWh�N}m�f�
ʙ97fa��-�P2*(�@ c�>3oL���wr��3��f\X���9�a�X*���E�r�p�ȑaA�	f�G<'�_��>�r�3-3��ѰP��R�>XkEv_�\����������R��Y�E����ǭ3�P�N�������O�*Ѩ��*�	E�%��$lf�i�,,�ɪ�SX3H���ע%��Y�2�`�R���m�[M����@-2�Ϊ�Ƃ�h��,k5�/J�v��dq���x�3�,MkZӚִ�fk��5�iMkگ�% �| �����j���&����(� �Eȗ��Q�[�n��h����+i<��P�X(/����L0�w���ճ|��
�����Fd���q��I����-�T�Q�!�-X�e�]ZdAA@|[��UvPu���C�'9�K����)[��e�!�π ��M}N�ע�kʙ���_]�95�QYW�gyQY0��"?S˥dJ)R�Z�$Y��m���`����v	.(.�	�!8��/�Vlơ�* v��_%��� <T\� ���rh�*�"�d���8ġ��J�A�Z1��LdZm�|��,�R���"i6�uZf)У� B| �XGj�1/eZ+G~�R)��"ԟ��6L�6+��ތt���G��x2�jU0WA/�B�uO���?�*e��X��i
���g�lU�f��f�Sj�Q��$0ۮ��V���� �8���۾�N�-�Q��9�V]L�#�),��<�%-YY�1Qr�f��y��מ���Z�@3@e�����KZz��^�@i㊙�dZ���벰�Hu@�}ˋ��]�A���?�W_}M�+ IaS � S!�f��[3Te&!h�:��u ��k�{T�L�Ն��糳$�zhe3@r��ّǏ�?Z�����G[��7��������C�CZr�sa]s^��K�扤p���*潼X���HV��0&����B�������!c�x2`�ϙ�S�j��m�#�K��;�����*����J5�@S��������y3�����8 �^Cξ~N��/�A�T��" ��5�����#ɏ�/H��bY� �V��j�@�(�Si�D)4(9RK8�>��Y��I�址�Ն�����>�Xz�˫y�)%;%=�	�T�h2�� N�:Cr5��j��s����o޼I�۟�͹cIE3NB�JC �U�
��O�t�a1����6���+0�����I"����o�ʻ��<��@����%+A�[�'�ן1��|�s������2�c=���[7���;$��m���ࡃ�ΰT"Yf�<s`&c�k�����Z�L�֞I��e�É�,/,o}?vk��;�4'ǎ�/�[�-']�wf�$?J�[�=-R�%d�vv囫W�t��+��_YY�*kl�Ɠ���*�8j) ��B�@��u�Z�*P�����0���Q+�u浰�{GFeg7E�{�F~�U�����_�	d�$���	l�I�8�ԋ��Վ�Y[��z$��y�#���3f�g�
	�������L$��|(!ZIl�5����<�sQ,i�Wjt>o�F[><��|7���C x�,jQ��+yk��Q՟X�Z�y%Y:�`y��Ls���9u|T�i�Y*�',��RMu�� 'SHF̩skS�]匌�CS4&n�T�iQ�=٘��&о�"�pC�3�e�=�����'q�7H9;�iMkZӚ��hҴ�5�iM�մdJ��J����E�VQ����VDz�UK���\+��B���pJ��!�?�?+�K��(�����!�h�E9�b���}��m�Pۭ¿�g k�6oeNT�h�lg�0��-,2�()b�k�Wj��2Y�6��MĜ���7��b��c��	�cW`=R��������ف��NoaU�ܫ3Z�T��R �.{�1����d���b�)I��%?�_1����|ڏ�� # A�|NE�\T��(����D�����1���AK���x̃�?�i&Gh�JZ0�"P�������0��L+K+�8V���R?�0nQ��W�DF,�R� Dx���.�l}�*�����Q�ࠬ�?gE�h@:���_��Ð��Qy*��g�|k�C �R�C��i��%诮돒6^�L��
������*��_SOՆ�A�(J�Jy�*�^���O�]y�C��jk��5jcdE?!<e��ȇU�D-�p�e�4�P��L{���>+��iQ)d�ª�}�5@;�. {F[����?wǽ+/ޗ�'ORi���S��s���狪^�Q�'�"�s6_1�3�uԍ��6����6ǃ|��uǐtZ���M�}����4�]C�`yX�69i�$��b���dG������e�{���
K���RF� ����& �`	��� [�I�r#�h�y����b��z�նUz����P@V|VF�a�?h��jm�y;Š���r۶����:Q�ϮD�	��֞iS1q��Y�ۘ,Y:�CK��?=�%�����/���-C�&ȫ��y�v_!*�C�x�ڡ��V�`m�瞒��59���
2��#���r��U����y��3�홮��Gr��=�}���5�����rP��gg�����1���Z[�'�ţ域}.wn�r�p�>���<�霦4-y��-�*%Q����E���� ��xv��v��w��<�ŅeYڷBk���17 ���A���']IX�KMx�}�)�� ���[�޿#��_�6G��[����r�UBy�����h�1ЛSuͻ�O˺�W����c���r��X���]��k���{嵳r`�!��/D	Ѣf�p\e�o�u�۟�������n}��:�v/� ��d�=�f G"γ�ۼ+H�W׊E���y5?UI��Ry���FX�0�G �x+V�u7+K�F���B-p��(�/�eF���iv���K�Qɂ�+���Iz�zK�c6��<Gޫ&J��+��|Lʪ���ϸ�4��Z���l��.��ʂ֊��=ʾ)%�t|G��g���b�����E������ =p�PR���~:���`�y�T�R����&�������ȍ��XUޓ'���C��,CM�b����l��fQa��Y�]\��������2���(��K����5㬤�&��Z�6$Z1�'�w����K�5�iMk�o�5HӚִ�5�W��G۽������^�ye�V���	Z�o����N`dR{t��A�jU4�o�f%
�{ר�,�b�ً�םV7x묬P�De�d�}X�O�x-��'aeߤm��e%��:�l�i�)V�
ЙU1�8�������/2G#˫�s=TO5ԹTL����H��_��_r����H��D�Z(L,Բ�
'')�?��DU�T��a����,K%}�ϫ�����A� k�� �u���JN���+��J:�j1n���V����N�,	�ָs��3��>���)Pd��7Jz�c��n���(x.������Z�A�B���D�}H�@��|�5F�a_%�X%ڒ��K��$l� F��,	�x ��S�N�+�_������֖���P�
��,��K0��9�y ��H�k�"$px}1	hZ�O�B���X ���j�u���Ѱl�H1�Pz�j����0��ߛ�ikE����$�M]R(@j *��Q�g<�h<�Yw����6���*LԦ�̽��!���X�+p�޾YV��[]a,�L�!-���u� ���g���q�@%<�a��=�c�����F��&F������AZ� �a<Qe
T"�D�?���Օ�zμU���`�3�k��ɚa)��p��$�\�������GY_A�1+��ٰ,D�**Ь	��>�����V�_����Iݺ֊�!�0�pm����4��n��K8�|�XQ�rn����(A����eӀ)��P-���R%5����ۃ񶢺{�D�N.���ڧ���CUk��+mY�P>��sW��] �^��{��ʍ�d��+�h����������'2�E�_q��y�����/�)��&�3X?塝�������dU�d���.��{��7��:B[��S{�����S~NlMa�5Qo~��Ǩ��^�Һw�|������ �aFǥ\t2�te�W��k���Ӣ�&Xc�P)*;#(�vܺp��C�u��<X�(�*1��C����-Io�KR)��^n7~�:Y	֋��zo������O?�$(����9x��,�2w<#��8�9��}��%~���� ��\u?��뙹�=vL�~�Z��/.�R�๛Ǹ�F-��:�#���ln�����O��|��dZ����h��[%�s��+ｂ�g)�Z+%b{˂L���
���A��>3tm qř��b�G[V��sM�i��yUT�g5�;��!�-mUa$	����a?�����:��1��d��	�GJ�X�2%����M�*D�^?U&�����f4岵�����3�-�ngZ��
�<,L���GA^r�`fHBRx0�zʕ ����c�FW�5q}���`��G�U���`T�>�~����y�s-� 2��z��:e0Ax�.ץnd��.Zr��z0s
g`���΃)u]����fd��<6��9}�up�HTc���yu|�D�����쵒mZӚִ��6ZC�4�iMkZ�~�-3{���b�|q`�ޮ�W���4��m^r�(� � d�4���-,�n{c�Ͼҍ�#�Hs�Oe�@��$x�+O~��.�Jܾ�C�M����-AT�k�5R	�E�b#��c���-���m�<���^�a
	Ѱv 2�K2�JB�X���s����_KF0�W]dz�����r�x۫�@�"��[�=Pێ���@���������2Q�wT��	?����w30�m�$e��f�Ğ��<��y���	�쿸c����۝�� �#��d�=�t��HB���B.R��¤��wQ������IZ����{�ۑ� �����~a���R}3ȇ��!+�qʨ��R�8g����PDmw^j�D�U�j��c��C8�6}�OF�Vq¶)���\$CNa�����V$��]��L
�������>���Dx���9o��"Y�<I-�A� yt�і# `\ҟ�;ۑ�p�6Z���EBW���H<w��$&���]�8��D@�L���Ƭ�5C���t�3o:��#Y]Y��6S���P�$	 \#(�����r�>]�N:.]M
�p1�#T��X�����'_9#�KjO���Q$P���m�]{5�6�[�2�h��lwFv�w����q���2R��e�ȡ���O��!29�E���;1+�c�:��-���o�~L[�t����'+��8�z�!W��"?��Isp���:���������֋粱�\�Pi����8�
P�XCB��3�^}KH��Ls��`����Z�#�u�:��w�5x��P]ѝM,M�;�7Ɓ(�>b�o���uU���i�(qs/dR���v#�x�$�9�sqA!�!��=�,��qܓN-�r)���c��z7��@�v�ݷ�Rl��N5�kn�Y�\~�v��/ �SdE�1:?7���]���0�+�և8�ʮ-bAj�%϶@H'�YI����X��
2T �+(27?_�O��|��?\3�R*34�����j,D��{�D��e��h����S����Cv�mw}f�9R��ck -�"w�<�v��H9�T�s(�
*��ڔ$=J��3����5��zNN)	�,C7%�=7?��gH���n�ߕ�\��l�`3֬�d\�#����J���qkӮ{N�~�{����|r>�I7��^�sG�M���d0��^W޼p�A�3n����(kk��Hǚ���C���r�����ۗ��#�Ǯo`�d)��n.a�<������k�w]o\����j�B��Fen]��qڛ��Z�dƺ;OU���+b�;��s��	�ӑ��J��x�{������|��TSQVV�<��JR~��E�:q� �cp��=%����A6F��	�k<�
�JU�d��+kq>{e	>��27;'sn-�nm���辕E�DG�!��^�߁Ua�:r�ϡP�����`��{Ȗ-���揪Lw�A_�N�w7v�I�/ֵ��E��A����ix�z���7w�y�XڷO��I��^M�R����OX��322�j/1�b���9����Y�f�M�-�"���8v�g�7ᙛ	O�|��n���-^�v���� k2�}<rm��h�D����� �P�\�<�*����t��=~{�R��\ۊm����N�瑔�v�xF�^�kZӚִ���ZC�4�iMkZ�~U-�k�u7[pe8�h�`�
:��k�2��I�/�I� zXDV��b�&@-V��U����pM!��F��*�e�$�L���1��tO~L[8���G������)�
+��B�r :���� �j2F����+��J���܇���ʗڦ����#{ɏ��SL���?k���BhU����Tej��z��Lj�F��+Կ�SV���������㺒O���$�H��eG�֨���׳��IKJ�-�m�ܫ���8�f������ͫF�z&�̌8Ao�����V�H3�ڿt9��DE�����@��i��3K�Ϥ݃�� �  � ��!�R�;�������6�ѕ��Y�0����P��t� AK���?!xɪq ��V?��R�Y�/> X��$���Y��@��t0d�*�.XY[����ܻwO?~L /�)|`2��s ������?��[k=�{�.���.�<���~J릊��>m4\�9 <�If�f;��*�`��*֚��>úr��R$Hc�� a%�I�`T�Ta��"�4����� 3�wv̐[V�$� �j`u��B"q�U?14�*�# Mui�	5+��ɗ@���peE���;r��%7��L�a@ �v�E�z��� �%|1�4?E��B����TW Hb�/4�E�~Bp��{kV��De���My���䷿��;���E��f��ѹ����k�!yp������]����mP@~ 8���D���}��P]U�5��[����B1Av�ݸ�!߷���X\M����|���j	���'��t��P EHb����>(@��7M�L�uڋ���w����$a� ]F�w�9�
#�-���a�O��FD���/���>7Ԁ{�1ļ��^�ɓĜ�j#��'no+H�y҃��eќ�Z�h�Ii*ieC���R�wmJ.\� �6�j��!��[�E��c��+��5�������t�;��*����+nLC���VHԉ���_� m
�@m0�&�k!WP}9p�J�̞�����>þA������	dԀd �q�\M=�V+��9��A�ڎq~���vKP��X}��k�/ ���Wrv笆��z����޺��e�����g���{wMa��e�;�����!����6����1� I,��*�'O����;�����a���4|<'ɱ��cn��S*�^���`�kHLEeYN�R>�A�Q��+�W����!T%.�O�wye�ON5�����)�֜���	�·(V�GT6
���,?wh�UAA���~,M����JD���kEɽ8u�1[x�)�����@��ޒ*�En�M��l�+]��K9��5(+�q��eVy�_U�4�J�������ݳ�$�VVVi5ףJp���ùe^����.��ND�e��e�@^)��^GkYdfeU��}�Y���syU���=�''sw�c�_�$j�&�I�伿gl0s��w���*3(���Nf$����>)����+�.�w$	/�V"I&]�Z׺ֵ�b���u�k]�ڏ��A�z;�%�@ob��=+(PңJU �Z9zV�Z�KBU>�PV���߲������/�ȏ% _�/&���.Bb�� �N�t =Q�D�
�W2˗HKt4o���(���@l�al��_@����#�����l�c�|}�m��UP�Yx-�ik'�����}ߕ�Ջ����4*;�6�1��p6 E�;��a����C���5�G2&���ǔ�z�&-uD���a�JK�da@����[[�TET�ڏ (x��ۑ�bg�@��d|D����Z��)j	, 6P?nXrA����OL!�R�H���>|�Q]N��e��Jh@�'�����3?�K�w�b ta�sds������#y��9?���,� B��_xI���=�s?��S�~�;�X�T�,��WA��gt(i����:��@���ܒ�2�;�K�~�
�6	��?5��Ï��������U�_����;9�?`��kR�k �Gz��HQ��l^N[)5�掁�8��/�$W��&���\�x���am!�4��g�� ��9ɠ�yI�E��E+�T���q5r
�!� ^����*�P�[�x?឵�՗7�xC~����믿�*��l�"�0�R�� ���ݗg����Ҹ	�'�n�E�װ�ΰ3�����7�qゆƾ����2���@�����<���={�D�V���A���&�D@�x|��X��Xu*[	����E�������q�v�$1Q#�ҡ`�Xi~O���
����
xq|����2����@�]�E����`���Gp@�j@�?��\��|����"T�@�Z��TC��H �h����������B�c������>ȯ����)���*����p��aK�����*h�����y%��f[�<5#�� �؂�+��&�R.H�k?�*-O���0��v�e��; ?�޻Mk�3gFj)X�D��3ܾ�c�޳f)�����i�ȟ'-�� q����7_-��ɯ�y���x��ʫ.�2�\�R�FnO�Bv�̶|��G���=V�CY�_�Z~��F��pl�Y2Ŭ�O�Tu?�b�Ƶ��O?�/�������ApoI��'$�<BͽA���;�:¨SP���������\0�u:i�*�γj,��bs[ɑ��Kas��m��B�y�{���P�k##̠��uc�����������Y��2�M���>�����4�TҸ���|Q��ڊ�����~I��>�������-��P�|� ����BY�cb/��o ��vЯ774w�jZ��lNB$	�W���灾2�h2ˍ��TL�Y�xq^�-!�.Hr)A��M��@�m���~GkĂ���#�o�{�;���{DE�}�������V|SK��ȕx��	E-�-N�;8�k]�Z���Һ�k]�Z׺��j�E�UXRt��9�v�=�EEبA�X�IK�M� �Z�/�*� � W�-�44 �) |ƒS�r�������@�ҐU)���q85$?���p&���0��l����&�YTKDV���s��Ğ�q6o�����I����6\��ƍ	jH�d�����=���{/qS���L�N�
V���TK��|�W���<Gkxo����ZV�,�g1�/��2n��q{T5����joF��͍5%!�8�:��N4��
�N�F�&��n�V�7����	��
��}��gϝ�dR�U� LE�0�7cVnNe��a�3P�Fg��٢�>v���	T�L&�0�����<:���x|L{!�a��� ����R-0Й}Ǌg7� ��m���{| ��Pvw��y��5Y �P�Y[N�l6�^ң��'�i�絆���\�Az�+���	UҀa+�%j}��L�lA @(,t@�z���a͂q~����kW凛�er|,�Dye�әZő����YP�e���i���Y%rϽ�I����������W_e�o��X ���9��Uף ���3��=+�0�P��x�����`h�����2ӊXf���csk[�\�"����_����ѯL&����ذ^&�xz]�ȼ̩ѐ����=����qcAB�����`�ET	��G�-<\US��*�yh�t�|�*�1  �������gY	\�j=F�������|��Wr��~��i��׍�!
ڽ"�QM7�*pO(�/>M�0�	N�=0��ɓ�U`��U�� ��U�m�A.WV���ǩ�2�fk�ϙ������[�'
��*1_�{_����NI��z���@c` ���&����nI!�k>%����%�yV$4k�3�w����ц�bU7S��!<� �=ܓ���q�9�@�SK��k*�2r����u�`R`T�/��v;-��,#�����������:yU��w�~��"^a��<-�*��(n���c��T�{U@�@@�n��T.ݺy�}ނa�[[�����l���y
t/����<._�,������gO�2��!���n�5�Z�YŚ�p��L���[����ڵ�38��d*�Dm鸜�������F|	m��h�h�*��	�@I��ć�G�7T��T����e��q��Z;���gn��8,�zT�ex$�p���ɫT��I�D��gϞrX__Q�G���$��w���� z�\�G̸��T��3΋��B�
1T��IJ���#�a�i2�;����+u��H�BkRj�=5Tx�qF�㺉�E1�4BQȆ�^Y����6�miji[�XG��d���SAB���@�	P��5y�[��[�I����IHT�z�����S��M��!�B�YT��}B�S#��{Xt��R��]�Z׺ֵ�~���u�k]�ڏ�1�ѽ>����0@��0iTs$U����x�[�����}kK����ѡ�<%~���C�m�2%(hy��� ����;����	�p^f����2@Ћ�0�+S~�?��`� 5F�`\� RQ�1��(�����\������!ELA"�mVa1����N�u��L)���?)e��b�Bx��^�'|/�/7���ȏ8m3U�Я5�{8֪�2*�(PPP빇�� �jx�s @ڐ�����_�J���Ϟ=��{OU��ll��h�ʪK�O�j��[����m��
����g��핵U���0��5�1 `� O��7�[���ϟ�=� �PVFk��oܸ._~�@(�=&���͛��?ȕ+W56�lZ�(r��ζ�7|_Ο?/�=���� 9�Y_Y���M�8����p�gE2 ��|F{"��Li�Eח����	^�*��X�m�6(��Xs��ڔ�b6�~��V+��9X��\�"���?ʅ�/�Ç�x0
$A8������)[[[�*"������D����<9���B��~�իr��U ?��adYQ;���y��W_� �����=��TC+ʈ$1��R+�\�M�rm����=_Ċ}��VR�w��e*?���dww�,b��������޹s���wZL	8���U,4�&X�D�_�ڬ�����TC?�i���D�&P}��¤R2l1+h���ȹ�����`�c)��A�\J#7��/>s��& 1l�X]���53&��|�1��(�Y1��	��֪����J����l�e0���b*��焪���L���.�5)7�Aܥ9�����x��-�w�̳��KY+@��h�Gsf�T�X��]�hN�*������PD��]��f{�g[u�Vj�\�k���y�5�~��%8jJ,T�V�^�3@�����zΠ�:l��\#H�F$�=pY�<Q��'�1�!���w�ON�um��"����D�$)�>!��;?ܦ-�믿�������$�'C*����g�[t�-��rv{Jh���1��Hsܾ�{W@���>�1���;�ʕ˲���vCȮ)�S�B��b1c���νt�yN8���3�T
��ak�G�,r��u�˟��|��'<w�� ���>
I�&,P	��f7ƑZ{2��2�2�^y�ZCƪ��3�U�6*�l\��>]�U���8��$ �����:(i��(��r�RU[D�(��
`��)�D�٧�$)-�[�\\���֋��t�-�X,T	���0��m�"��Ӣ�S��h����V�F���bڹjv�eH�qMdμ�܎��<j�	ݰ"%c�()�om6w�e[�����4m�#+�����c��C����y�Rv*�N֒T��h+
[7w\W1��(Tu`ka>�4��(R�ϯi�V\X6HyJ����p�+U����I#�K1H�#���Ʒk]�Z׺�Shҵ�u�k]��4����ٞ��M����Yjx��%r��j�h���Y!;����y��⠵[A[�y�PB���p�!Ȑ�y͸(�rIq<�5UB��'��Ӳm�vy����& d��j(��� ?*�=9A,%K��Ԅ{�Ixʭ�~Y�{��s��֋5p����Jߐ���"�S���c�_=@.��?�UKʄ�,�gzJ�R��Ar���C�ި>��T5����	�� H����T� �K
iI%��4U�u��q�]����7�`�~�J�۷o8�=*�Ϝݡ]	§1��77�W^���3�a ke0?��(�5Z]�`��] ���&C��d,iOV������9��E���/������g�ԉ�;�e>��w�}';;;� ����
��ÄYjUU��@��֦�9w֝�U��9�D���"X��A݀s)�L��9~��������,y��`���do�sF ��V+ R�z,hI��k ���;�����͋y,����<�_.]�N2y;;[��}��!�a����� ���q���w�s��d}s�}�&�� ����LV��t�ǭ[��������w?G�u��,����,|J�Q!���&'%j,�r����=9{�����������J,��b��W@5���=���/䫯��'�5����hcs��T<W%�^ch�@��`��ٳ0S	Y����y�+���s�[��á\pk����`��ŗ/�ao�8TT���Ν۲�����_L��v=�
S�~.0���g�K����������r��R�女�x/Ɇ���~��ؐ�)0u�>�ϋ�[w����\��;��$�����y3�
�2 �Q���Q��}�37�^E��eq�&�l*�[\���[���Dמ'pZ%�*�p�D���se
N�mUH�K�����^i�j�����u��^{��f��~�h��j��'hu{�TR�d�Hke����wF2��d ���!T�5J�Ƒ)���Cۓj+�(��U��8��1u=�-���P�(i"�ڷߒ�)��b \��1C�H�o *�Z/�9s�9G��q�F�����󅑅 "���I�|���r��od���2IUHB;���ڈ^�kTg:��+���_����T�Z(Ь9�憎��x�P�-�1a��h�6���i�c���Ϸ枅7t:�$���?�	��ǊE�� r��'<�G�+��U�ڣ!�&!I�YbE>m�SU٨��a|O�:��Tki��T��E��bCM�����,�t��a�i��T�� 	$��fQ����}g�J����y6�X�ɀ��2Լ�(Pw�w׽I��*�N�g�8��B�3�U6�B�:(���n��������&^���x"�5��]i�r�Oa����F�h��*HR��r�ޡ�'�ѨO"Z�u۵�u�k]�_�uH׺ֵ�u�Gժ�{�|�Q��B"<��Zm�+��ON��L�BOk��2��V�Z�zě7=l���yx�)E�fa�����q���X��أAM��?���\ �h�P�%13$j����K$D��RaE8���l쀼ʡ!^��|O!T��CBS���x;�V%���` H%�C���E�W�k��Wvx�ǋ�����d�PA�� P̗^,�����=0���<�&s$d�D/�އ��@C Z�� )U�K��~���>¼�@ö�)�_��@R!�u}s�
>��
������cXe�YIN���dBpjX����M�r�7� ��V�C��.���d@%�$ �㈠�'hP�j`T�B�p|tB�e=���-ķn� �ɱ��9>~�H>��C��]��*A7 iL�����R�m �W6���!� F�!_B�ͷ��`�����/�2@&��ʂ�̣����[��w��X�G��Z��U'T��T5$W	$*v�#�Z�>�&}8��p����0P��T���������1���8�#�8���'W0�ަ���~b$���c��Ϧs9:8�o���$�AX_a?@e�;����E�6P��s1j�В�BM��
����F߭��7ސw�{G^�p�` !T-ӷ?R[.|�l:���_��W�R���SC��5��Q�P"���:6��q���o� W��lP��͕0%� ���\y�U����r�t��e +g�Z�4-y���#� �W�X�� -x��P1P�W�
�VFdv]�-�	�߫���_�����_���G�$�K� ��X�A+M�O�p���q󄠦�w�j&w�ޕ/>�č�=�%@����� �����iV�W��@BĈ_Sy\�wfɈ�ӉT��T� c�vE"+)RD��HāP0@�笠�$g�ߨk+l�J#�R-��"���"�����'�ˬ����W^ ��e�p�Ȱ&��B�Vd%�l�?pѺy�su� ��_�]c��UN�&�4�/d_`�)�c��s�ˎΟ�&�F�X��k�� ����qU������?o.�^z�{���V�$W��4��2���@���w�z�	��6�'�������)�ަ5"H�,��B�I�{.�PR	����Q퐴/��.��)���@|��'"��M�D٨���R�ֹ*?�>*�k#V=�+6���3��W��R;)\���1�"S$���s^IL^�@$�V�wF�Փ[.Gi��M�EU�{ )�*��}E=��k%�r��$0A>�y!��s0�����m"�Q]��.�b���`�ϕ/H���8���S���Y@����2{I@?�8���,-�E	��9�B"Xg�c��>�Oi1�^�U��q�걂�\�aRZ䩒�{��Q �p_���X}	�mҨAxϜ�"DlT�ýn(�Z\;S#��י����mH׺ֵ�u��:�k]�Z׺�#j�d-�ά����>�}�K�(h�����<�c�*β��f�+b#��*��j*�,Z5�3�`�J���i�"�v  ���$6����� 0�B6l� ��r}����>�F\Q���ʆ��N�C�2'�q�U�才6\\�*o��T�Yކ'~X�\y�6�<.B�1/R�����XnD��J�")`�.H���>.<������ٟ3Χ	Do�#�:���6��/�O`�Y�K�4��0W�s:��"�� ��lENM���<谹{FF��{ �` ����	k0�u ] ���v ��� �#N�6	� *&�5[����=�z��F#$P�j�`��G Nr�n]�xA.]�$�kk��ae�Ì��|:�k�}�U	�kλ׃���	 �ñ6	�j��o��!�ws�P�gvHR�=n\�D�ޠ��a�H���l�l˕+W�����k�����V��Ђ�#���������K�)p(�?�$2�\���XI���,�Wõ����s�K�Á��}вi8��]�_���?��o�OU����3>���ܺqS�ݻ/�t*�nΤ�;���ɚWL����Ho;W+��� V���}���
�`��Bu��]]Y��t��ǒ5�%]�j�����W�,V�߅���l.�$?���Ӫ~��S	0����YH���P�@��׽���?�7�x�m��/)�nM%���k���^��xF+6*I"fa�3T�����=��:E@��.ܚ�����ԲK�Z���K�/��~���-�>�0r��B�'U4���,���üP~�S`�C	���4��P�!����d�f�~J�i`y���~^���)$t���g�I���ZP�}�ͭ�j��I ��
p'f]��E����82Z��?�&��j6Q���c9 ��fk'^����� ���x_`4:�E�Z�' �bS��-}��_�c�A�O1vi��]f�F+���U�]JT{�'�y7�'�8r�^���3������P�6�dv�vs׿��yճ>9�e�؏5k*X�^df#q�=U*�P��ϙ��z�`O�������S�Ɛmw<���
*%�UhUf���yn�kܐ�eS����H�,�	A~\��ý�w}¿UaU[ы��yN�ۢ�'؛r��^�4P}6ko �2+2�H���E-O�]���BK9ؼ�g��a��	�!���L*w� �f*��)b�H�s�*tM�6�bS�`LuO�,X���cP`������|b�!�!��nNU3Z@��}`Yql0�率�J&ɒ5��'5yQv;[(߳(���*j\ǰ����������RB���b������TR`k��<&��>A_S�{B�V�}��w��R��G�1n�%��XǮ�b��ƺ�k�dxmw�׽��P��:� ��u�k]�)�nw�Z׺ֵ��x�e#�}��++�j���:��|QE�2�ag<>f=�� �XLX5��7��lA ����}�p6��)�X'��= �Y�l��ӽ$PS�������� �=9ƍ�D���ߺ��arU�����L��8@�~�2
�x�)=�������Ȥ��Y%��H
�)	c16�f���_�9�TU5�{�TH4��α2$l
{�]�
H-�Ǚ�j�BЭ�@O~^ت@xj�Bȫb�����@�E�/?C�k�]>��@m�D�q�o��a?�"8�N�XAKp�RrTW��%��}�|&�b�ߣ0��JB{3�U#�2���  q܇���Ѱ�*T�0\�$H�Xh� �`������h �̸p��i���l��+�KB���Ю4t�p�;�E�� �̧/P��ʥ�r��M�M'$)���L&SV����nή�R���$a�n��z���:%+��Qc_��bVm/��j:;Qۮ���y ��� ���N0�f�5���榼�����K��p���ڵk��g�ʣ��	p'��	d������VT�KzÞL�3���*Y�#����C���+r��Ǳ^Q��=c�Z�L�UZ��ᜬ	�eՀ�a6yh�#�V횰>�t������O>�?��/|]��u:�q�b�	���X��A�eV��w81��[����Q�8�5_�v^��Q0W����1�u��9&O>��C��-��@�oo5s{K\%f�5���|z�m�81W r�^�Wd]��7F�oP|��ȏ��5�l� Ȋ�B���g�i*����C�>����sMc%i� �Z�:?�PyZK8O��f���|��q�W�wh`}�ș�@�?T�,�sS��p �%����F�5��.��A~�eՌ@l�1��'�Bzn� �0f^LJ�۬�u���� -2W��;O�c����ϑ�X�kȵ"[sCj�Uk�;)	��*������8�n��696�J�U��z���ߛ��T����Sv�����j�%1�*\G���"?�E��'����(VR��w��el�ΚN�{!�ײ��I�; Ȏ�U�f1K�mJy{E�{��� ��3���I_fV�j!)?u}�����s�W�r�܂$���'��* �뢪��@kw~��̸��2�yު�����'������k��J��3�%�/��!�,J6����{(��o3U�����ʲ$ɛ���$����u-84�%>�F���/�{1&�Yz��ױob䯘�(TG˶�|N�Fm��9�/�$��/c
�环��vQ՘$9���v�'(�@�d�Y�NUS@uR2�ߋ��c�b��p��nY
�
Z�	�XR�p�\������͟��]��� !=�8��~b&��~���@n������T��E5TdT�t�7���1��p�>?IUQ	߇��=��d<�u&4�+�'�z�Xe���
KU�2}�5�kѫ���e5������ebM�ek��X�Ė�f�E2*�����D�㱬�����k{k��D�Z׺ֵ�h���u�k]�ڏ�s�FV�Gԅ����� ��ʈ�&�=�\����r'��Ӫn�%@B �
#�:>����q�� ��0Ơ�J����$ �Ϻ��崄���E�::5� �S�����Q�*��Vk9 T-�"ɪV1��s�߳�o��q�ZR}4U�m5�O��y��yܴʴ<u��O�խ��ׇPV�*��4�Q�S��0�J��'����Z9M�
��;}�C�D��v�s+_'".�C4��؇�V3nU�|�6�A,P3�5����Ze�T�� ��
VךL`�HP+є��|i�x�Y�_���Z���n���<��S��:27���J�kl� � ��7~���M�sr���M���5���,���� �ш'G��E�|��Y͟Ii�  5���ġ�JT��\��om��YP[���K<����rx�/��&x���I���o�����d��ZPYV@]7^��2Ά�b��(T/��T��q��A3�S0��P���O�4k�+@�������裏�O?�^��z��\�n�	�{҄l��Z�p.��<'�$YU3/�~�!��U�)��`n�>�l�r�js!���ܻ}�J��ÁZ�dF�b~ �"4���u���>�`V�&�:XB�R��� }���s���{����=�jpO��Z�[�!���w�w_#�?`�vBŉ*V@~֤ټZ$帢+Az"Ä
�(4������{�^��;��G	����D�~I0� {��w}�skd
�ϽVb��4T���ύM�c�P_�t������z��TnVc��J��B���� ��{oI�Ϙ@jhj^3�6$��y	 r�d��'���@��\Z,�M���s��(�P �VԮ=�7���s�s��yy��>�ʹ�Z�d>S[���'�a������}(�"��E��[~��,���^�cwg����D�'J����y�o[�ۜ��8"�BA���38�R \4
���NW�<�@A�`vL�q��=�!�'T���o�rIG=�Tbh��
����Y�78g�fG�,�#���ASl.�nݐ|��������=�`4�Z|���
W��ɓe�,xM�vG8���f��:��`����Է�� �=��7_�c!a���-b�U>󣹿H�fM�gXk�V[v��106I�7#+x�I,�M�;�\j^V�� "5�q���d��`
˶��J���+�П�G��s�h *�֋ٺ�J��d�/M�|�%F��A����a��ۃ�n_���8_��y߭�L-OYT���̭��֣�4$!����ƚ�jU\�@)�j?�*�t�t�C�:
O0ql�.�X� �_ !��8_{ ����Uk�K;̢�W#	��`h�
�!��x/��8Q��çݳĪt�k]�Z�~��#@�ֵ�u�k?��m����-�S+�=��H�?�� <��� �'t�ZLDؒ
��= ��2?�O��qh��PI�S.�3`z�sz���ɵ"K��������=��X���
zxJ��XVux+.�mx,�[Tf}�_ߨ&Z?mZw1?�%$�:�=^U]D|hG�D�~���z=숀�0Z1.�#�� OR�B����a:�5gD-��s�uBcٵܿ8�%"d�������J�pROt���	���[8�H2�-�Qj8ze�j�Ȫɛ�X�\�ml��!}��K�`"`Q����
��n����P��6먤$��ا��	���Z��h��I>�

"��蓧O��/>#(}p<�˗�ʅJ�z���}>� :αVeGP�MFpE�����^)@�j�H+rae�#(ܗQ���뵍ON����V�\���c�� p����TP����di xݐxI�C�iOTkRD�o����f/E�U��g%�V��}�4�k��hi����M������#�\[��֊9c���ꠐЀ�&�a�>�c�x���F�X�c̟>}��<����2�%�.��
�~X[_����g���=��&O=�0kT�/4��-EKp����	��5��T����f���:/P��\%�f��un[������������6��l D8�=M!�<��]2����K֗n�1u[	���ROV�+kF���T%�|�����w=�ہ2�}ȼ)�}�`�O�>ɐ��NAͥ ��5�:/y�naB����9ws:��>Ԭ)5=��-��;��96�E���P��B��:����j���2^"*��^x��</-��1{�P�à��-����S��2l�$D*�H���� kA���%��<�����������{���"��(��Cڜ�ڴ��#;;�T��c�C7���|=$���a���јk?G���C_?z�D<�OU�[�-|��\�|�*8�{a��a��/�J�U���Ucg��œ��h>��˱~ <�^%�L	���OT�3�_�����t�=��3�}�}9w���y��sc�,,h�-�����	�}��#�����3����8@�"������T;Ī����k������}F$�F��h�+��gI�^��|�LY.���0�Ӗn�H	���j��H���������A���*SXw��&�O��W�a߆Ң�"����ZP�@yB�93T�C5� �,����$��]b�)A�dS��Ǵ�Z�Eձ�_���=
�2:z�Z[Y&��*��� u#Z��fŧPa�:���^7���U+��[0:��U���f�5���f,�z��[��=#5��2'�C���#�u��kk�H�ܚ���0A���#��ao��d���FfӅ������������lf�#[�,��]W)�'c�PЍe<�ț��*]�Z׺ֵ�^���u�k]�ڏ��M`�X����bG�(@�$i���F�_Q�J°��`�u�%�t��� ��n߭(���^
�H$���O,�2V�o��~[������3EH�\��*𾵿�?YxZ���_5<���b����8����>aj9!y��:��BRR��§H�K�]�'?�%�hu��� #��Gx�/�w�A[�K�j���ư���:kI���%���Wppv��$����a;���L�_v@�CRk�k#��@�p�J���3x�T\�����{��s	B�6,�}@��Y�0H��o
֥�1��l|�f
�A�P�d�g��oH���}��ܹ{W2�9+�5��|2��`�̒�#���O���=���%h��ꫴE��Z7��� ����7	o:+�
LI�gM�I.>��0��Q�yP��\_ې7����������{��W<�X$��ڐ ���J� <T���/X3ŚB��!q��݋)�^ꎣ�L����Q8��s������{'ӱ���s��,���0����XVG+����\�����c<f���C�#j��-�|�3I������%�@5�˘˰�B�������6�YtO��v�`@�_���n����Uy|hT��8��E�Ms@��ș�
��A�X� �Er��*�ɶ67���q��s9�{Vs,J=6� ��^�P�0�������In\��������*��PvfwWVW���kn�9#[$<�1st2&����a��X�����~*�Ν%����3�{�.��4TI���rpp ��ܗg�{���ά^��O�\=<>��Ԕh�*��O�WV��/�/Q�c��Xc��{+���o�J9�����<e>P*J�I����J�F�D�J��@�:��v����r=�	P.��L9��}zW�q�1�A;&�A��]U!��	��o���\�|��F�B�ѧ�����c�� s?�N��6dJ<���'k��.�/|�����;�9.�Ɂ�Ԛ���f
=ϝdF�T�WFBR��B�n�]m�&7��2[-���ޗ�3f;{Hy� Q����P�3�k��q��w��c|t"��ÿ���Wx�~�L��ܡTm�@ݺqC>����|*<�ʝ�!v��e�]TkQ#�8�*S����UE���g�����:3�P�יЮ�h�ShV:�_���G��7Ue��9�ܲ2bE�#���58~����J`�b�X/�&�s$汨�3�P�P55�1�=��G���V
d�އjQ�VD�$V�v��Z��͘䨪�p?�=��(��@�~W�XLŉ��9c���IId��_x"��D�ֈ�����Y][Qu��I�D�-�~@�g�HS�5d�*wW�=��S�/���0E��s6�'��r�������&��r��gw��12�˷�a����i"s+���87�|&���E�I׺ֵ�u�'�:�k]�Z׺��j��C}hW89lH@
�-�P��r��apB�Ͳ�2J-X�y&b�53���R�ӝ!��z?�$ԧ��}&��������f)4j�z1ܤ�eu���r�4�Ч����Z{7���i_���/��T�9*^��$2�:Uv�E�J-U��X6���6�(���<�؝/l����� �ŃH�y��Ј�R�U�wTa����JH�Ѻk�"`�`U�(��g�q'P2	�0#�h��t���DI�[���>_��
i.�Ĭ�5 \=����|*'��>�����P-�6wemc������rttL� ް�Z�¡���U��6e!Ӌ�+ � �A�'����*�FC](�ΙE��b�!V������y��|��r��]�����O��G<��`���7��ȭnɝn��wޑ7�����lm���14Zm�zj�$�HZ�?w �0 0J t�Yu����Ə��?9�O�YTA����*ww��y��>�o��s����Q�u�@�"F�F��q�����ʾ]��l�iL x#j��Pg���e0�;ߺԐw�-����H�={��± h�����Ͽ����h��w�l��v�s�fe,��<a�٬�WR�ߋ��f�[���9��f9����1 ���or�r&l� н*v�y0����9����?x�,1s#�	�i,�-�8�O��X4�s@m�f���~��K��/~)��������h=�*,�3���J����~(7n\������|r�bN�w~.��o���N ���)����� ���noQ1�k���4g����hU����Ǐ�� !��������p�<�ߗ3;g��ի<N��o��F=~ O=v�{,{Ϟ2�%E�E�3r��G�g9�pcc]��y8Fv��5S#�aH%���'i�Z�V��V�O�@@p�������u��*�n2���c��0\d�L�Mt�(jm	Th���m��}_A"9��7P��˞�a_mװ?`������x��c�����0�TZ�c?q��6o�c��������ʙs��.�z/��=�%�M%���j��~��1�5�V�S��Q�Lh狆���C�q�t�}2=��]�Hv_n�߸~�K��9����ѼҼ�}�a��5�����_�,_~��<�ۓ
�]�WS��p��-��P���2{��Rۧє�.��ƚ��	6΍��:G��ϫ\0�5����yqZuid���4��
Ip�ͯhf%M�h�q_���'@�A���&����WT�����5� #@���DER��b�7�}ҦO�
)j���������X$�k%�.�|���W�{"��A�U�k1����a8�� ��d2�zP�9���	�U�x�I΁ ���\����k�nެQ��1�J��uQl���*�H���OxM�
� l-�x�������ޗ@�����ڐ��mYsk��Sf��B����̩��9�6�}�G����Ǫ�B�),u�k���(b}�-���J87��"�h�|��t�k]�Z�~z�#@�ֵ�u�k?��܃�P) ����?��GjE�b� M��f(xe���`�~�JV��Wb�V%�������VWm�z	'M垰ڻjh�YeA��L�S������&���B���U����[�[����ϊӆr�o!�)g���%��K�1-Y��ae�Xi���U./���u�ߥ=��Tc�8�B��A��JF��Zv�
�l�ΩX���?�!8T5���+Bi���w�Y�E��V��̇��r&�h�@�R������Ս�2P�&ݢ����?�.���C��ӣ�Z,���U $&��d�����ߕ��HN�'���#V����B; ؽ�O	 �F�9�u%�Gc�!��U��ݕ@�ɉ���j�5�h4����?�'ϞI���_��+VK���̷Q��A�&���X��Lg3���yP^ l�܅sr��e� �Pu���#}�� �
Yp-����3`��pm���ٯs?�}�0HYU1��U��AJ;��^}C���� 2�jA�����|�m7����^� ��e�y�4��-*j�2�,�����!�J�%�Ưb���T���[��V���/�X�@֭ѹ�[ R�LX3�.� cP�G�/����K{������-fܫ-��^ �1�d�	�b|q<�B�
���h��/��H}�2qcw��-�}�>��c T�w��R�g������ߣ1�h����^]_�w�}O���?���@��~�EX��ڵk���nߖ�{?,P��\7f	�ԝ�����+����	�S*8����ڔ3yf
�����ٗ�JA]���������}x��p�b^���U7���A�]|�e��<�&��ܖ/��\>��Xfn_��Ԏ)g��,����8@�<~Hஶ*�$�e�Q�m`����:��
L3Y0o  *љ7�WqT���d"~VG��Ef�S5�|��FĨu�����J���T����#\����F�d�t>@sի�p>O��8N��-�'��0;I����*�T��+���I��r �	 ����D�in�3d0����}FCk�*��*���X(NЌ' �8fX�AU6XJR=�kq`���[z�PF�X����
+���o���3�}<�R�t��u������;���8�Ywq�9��j��HI��8Doװ���Tѵ�=&Trd��cS�aO��B��Ȧ�(dIM�����9IK�|��f��~�q���Q`�/"!��X�E>o%�$p����,�{�L�D��o�oFB��^?���X !�����Uns8�=)��{��v��\83X<ι�(Q�资�.7F��K�} ��<��p(�x��k��U7���h(ђ�5�d��=�׾�8�l�Ø߸���^��B���V����ʺ�WB�|�|���>"����{0���sONƖ�4o��Na��Jv��]����Ց�gؕ�.��}�AВ�jG�{�Д.gϞ��]��y|t̢�!��Հ�*Kl}R�k
]f���r߃kF�f�UJ���^�����Z׺ֵ����:�k]�Z׺��k*�7�g ��(h�ϳlF�����'2� V��އ�Ҫs�&���x�����d�V%�'jU����sk�Dx^�j�����P̀�~෦��$��t*!
Uk�R^�ᒼ�N�d��;��@K�V�����XEn�hY� lL��T�r��ޏ�	D��� �>��3Y:TK�����RU�=� �b)p]?���c�~�/:�W�K2��͟�~�e��P�ai������4���Zq6A�,��BZB�Z�}�Ve��7�'?ܾɪ���#� D{x���UV�fS𚐠¿AUA-2>>&X���!�^Bp�����>��b2���Ώ��lnm��'��9cvª��  tt2!`�d�p0�2��FR�z��F��B�HaG1$���ܿO>z k?��͛�e6��W�qllo��������6��5�c��Z�� �W#���ސ$ə3�����d{{SU-�]X�jQ-d��H~��������!%���ܚ/y�Ț�4� 4����?{�G"���!�K�!@X�iEj��R��2Q���F��?G��b>���r����_���׹o�pAEoQҶ�Am��XI��)ȵ���� hiE͟%�W���QY�����sjYZ���.諯�v��$�g�7�"B����7 �w{�ȍ/��y��d�<�q{t�~�b�;`U��"(�"K]2k���E�޻s��9+o��M���~+W���,���0�%P��9n<�ܾM��'��*%��Tz�>���Y�R��ޕ��*���5c�ݚ���=6��4H�y�R� =���9��7�
%��y]�����]�C�3�����^���\�� �����Q�Y&��_��6xY�ٓX�/�$���h6txx,�ľ	���K�x2Z,�Z�쀙��R2h[@�NC��:�*�GEm�5`#�|U�P���G���t]H�1G;΋��j�A�Q�D�����j���4IɃ���)�.VK"�/Zj�?�E�` '+�⁖��D��q,x%筁�P�֦8`� t�wĭuSZ�Y��x������D���S��E��%��s�z�4�2��U�s� ���F�����ZJ"�d:W����~��k��~�n���/?u{�}��f�۳�A�_e�3+Le��&����e����c�'Ya�58�f���z��̛���k���Gj1j�
��y�I�89�*����|�������~���K�Bu��C=�eҼ��eH���U��[sXHu�`�s���<�s��ݵo�嚙�^�b^�Z�����o���4S���_�?h�Wr�h>�
�[Y��3w-�q�M�,T�w��h�łw�u�5O$]d�=�Q�2�k�$���"��{P*(C���֚ƻ��dH"�'6��P�jie��)��'7p�^1�d�Ϣr���r����|μ���� �q_U2#��i5����\=tt�g��7�v(5C˳� u9UԵ�u�k]���� �Z׺ֵ���p��V ���� H0 !� <��!���S���|x*��]����I��������j3DԱł�K%A<Ӡ���O1Cc�8�D-�ѐ%�W����6@�{�/}��)B� ��q��� �,D��(��k>����1���Yd�Fm��Q��7�)4�,b���������ꨘ���U5)�RȪ���4�* 5�&	��*w��\L�@bܒ�_�C�Az4�M5����)y�G�i��[�[3QT��$y1�*_��� +����۝�Gu���ۣL'c���j��/<�I�~|����!I�l^�b�&�踔�g!����g'�CDB�=n yQ�	�rp2�G��<a��6�$�ܥww-����������cA�n:H	��)*-h`��P{�d��U���l�=x(w��#9�u�,y�HP[(xPk��q��v���'}�#�����!����+W�ʙsgY-��F2�-�J�<+�P.�?ۣ����[��5,�a�G�c�������}�v�|��G���Xs8��j����⮟�Wh �z�͊�|.++�ܓ�D�U��E� � �d����}��$����|L� *�J��Cu3��U�cR"��*��[{2N�����P�Hr���}���!+�A��>�+�\�� �.-ه��]�Cu�ٳ���ȇ/�hu�l��&,[����o"��]���c���U�^�^�XQ��7�ͱf�������S�w����$�=%We@$)���ٙ�s�������P��ĺ��|�7<�s����B�A���Cf���� �+�+���j�YX6�.E9���-�?��+�D�X��I�.}HU!�ƐJ+������	�W���|ϡv�>Uf�R�iT���(�vN
��~��+�u^�A�� �X�M���P��w�9�f/�!2pP�>_�ʈ	lj9E�#Cj�6�*��t�˦�'@HVY�}e�VK���y���"ݳpuj����>e�`���X#�KŨQ���Y$-97�F�B+#**B~����ڈ7����=�r,4;!(J �fP�U��9�k�3EC�����X~�uq�߻G���ۏ/�|�
B���7�ˍ�7������n��e��%�I�@�9�"�a����b���oH��V�2��9���:J���	��Q(��*�|�*Ҍ�$���0�B#8���M�����IF�ڔ�
�'4��ӫ�|&���U�6TU�ip�P���}����s�k�V�����9�n3�� ��(. ���3^sC�8&�VFH��V��޵��64��@��ir�0�n}��)M;���'�B����!ƹ��i_�8�~��^F�0+�q��+x�'�5��gj�B�oc�-�8�T��
1��s}��}�ҝW�c��ؽ��h:Ș�
'݃��e��P�f�Da�k�hR[0UA��-����+;��Y[���J�>��"��2JIj�\_���Z׺ֵ��4ZG�t�k]�Z�~T���HSVyՖ`�=�� ���ڳD���� �t\)�����ȏ�l4�J(|)++ �2�Ky6S�F���K�p����V��?��2���e�RN�o��JS��o���(�J�$h��"�!�a��!���G�,	��*�R�����^�����l=���~3Q��}�}���x�ǃ0&E����Kd8�����"I�	��@Up��%XU`��T	��1+Ŏ�`�f�Ħ��B�VV6�b$$����3X�?q^iu.�K3]\�[7�*�ZOU�����v0�U{��������u�_%���W��x,O?���g�Ǽ�8�,dRju&�6�kũ�z����̠�U�DP���/�[�ZR�
$P� �5	��ʺ�  Ѩf�������A�l#˪�
� �A��!D <�]���aqs���/*31�Q��9=��X�"���LU�t�r�اЀ#	���Zx�g�M���������y�|��_�/�[	w���BaQq
{muC^�u��ۯ��{�r� ��nʼ�4�b����G ,ss��'�������XA��MF�ja�X���8�
U���J�#�Q}����2d�Ǭ���X�X�MM���<�*X�� �Jȳ��U*Q���(�{��`V�M%%`�^��+d�����,� ?=�WP�������c��Oi���?�����T'��#������5�~��ڔ��U9|�����fB7�:rc��s�Ô
V��\2���HH-���X�,A��;'��ￗ_��7��@V�' ���:�Mu���?ܔ���o$�N��Dm���:����� 8Oh��tfP�lkǦb�8F�DB�{<�5�U��Z=Ł㊤Xld� ח)@A�>�>�6Xq��|�5Ow�CZ�\�o��'���C����DO�h|��հ�ӭ?��W�q�T�=��H��V��8@c� �x>$ �j����͹�a�����H�Ub�\.V�'1}̹A2�!�*\pxe�hES� k�$�Q��>)*/{��U� 2b�-P����;����YaaȰ�k[��	(HA�x;��T�q������OC�+ǡ;�a� ��5���i�ƪ�4 H�l��nJd���j4�K8e>9i��1�Ύ��|$�J��&�c��ͩ���M!M�>fVX�g��'�W]�7���>���nP���9��̐��f�xI�8�n?��12CNA�X�n�f��3�{����Z(���nIB;��lB��M�L���|�׺0hs����~��$A��!x�%jE�9�j~SH�t 񇹩

NQ�X	|swLm������-��(�c��������\D����Sq��|e�Bp�˳���IOI�c�6/���$������<u�]�c\�=0��h�kd��u\O�z��P1Z��3PT���ޫs\#���<pm�|3w��$8wX޹?v���wȀt��3�/|-�?(bp{@��������1Z,
#m�U����XՑ _kw\+��N'\P��n��}���:[��L8W��@,�<r�2��;��=��x/����5!b�*RX胵�{3�7Gx�v�3�A��8%��Z׺ֵ��$[G�t�k]�Z�~D�����CC\i��,�y�/�!02�"3��ѵV�zU��L��� 	�8V5��m8�j�	?��8�D�$���� ����l�"M0̪{���*)�H�7+�2_x��t�D����H�'�� �EEs|$BRSK�w�/ٻ�!��!H��tu�Z��ʣ%Q�
�H�G����>�����
c�يC��=��B}P��͢Kɔ�!5�;Z�oJ�4�EpS_����B��!��m��c�cE{��'T�9��{������PA+#��m������Wj�B'h��X�R��1�vC U���en'���
sN> �
��<��T!.j�&ɃLj��5	�I�9��� �r��st�h@5��L5 @���:�4���
.+C� F(��p��m���Ň��}��̦��U���%!C%���q�S�
� F��Od:9a�)*�w����˗8���-���>�I�|��Uc�o��(��H؀���43����2eW)�lB�I�|��v����G��bք�p@7���Z-P��W3���+�*�"�xN�/վ�\�F"��y-�W�����x��1�e]�^$�t.�ل�) �B�� c4�5�j���6p��1J�={N x0Z���-y��7	,bo*|�?���"�b��ybs��mX�J5����}���d��l7�8�н~�̀^Oַ6������;�svW���*����.�"�خ�����w�|M?�2�Wa�<�Y�@޺�������#���eYY� c_A�
������������ޫ�+ ��"$��D�YnJJ�Ǆ�Nݼ9>:d&,�2(�"a��(:0c���V�P"�<��ƶ�u��`O���$_L�ȂU��x��H` b�ʕ@wK�NM�玱1��&C���l:j-�:a?T/5���k���|R�x9i1\{�AQ�܌��B���5?�w�k���|9����g*D�
G^
�K�����Wx�B �ڒ��anL��O� �"�Y^��]�h
��
,4=���C�j��j� h�-����bo���� ��:�2B*���Z�D�NE!��J��@���k��F! ��MEUG�JUph�:�C�P��0ln]�n}��*��(-�B�u(C��۵��G!i�%�>mn#����X��6'�f-y����\�N�s�aO���t�f$z�"n�#�Hxϡ
@}��p�M$���z��ukfA�Yl�r�`+mM��GSf�h1ζ�31�I<�J<���mT��hnI��~�<�q��H���{�����g>=!Ʌ%��7.�NB�?T�မ+y�dR�2�ǣ�)��0���Gf���5ײښ5��{NL�Ԫ�H����k����T"S��$r�vv6� ��	2��Cw�s��MQ�������JȒ�r'}2��8���^��ֵ���%�s-��j�@��	H��YNP�y�F;;in��ֵ�u�k?�� ]�Z׺ֵ]� S#D�X��A�YRy�g%?j�K��޳X7z��3s����֚B�B}"�p�1r"X�i�$���?����:`��ʃ�ڣ]H�
ֹ*8�&jՄ�@����L�=��b����j���\��,���*B�����+_�\��`Ɔ�WF�������(~_�xi뱶J��a�P�?�*���8��U�#�I~n�?���c����ȩ�J֠zZ-kR��
F��:�yh�7����s���gxgؒ<,U0]��i�Q�l�a˙�@�p��B'�
�\ fפ�'S�8����e�+���� ��HS��ͩ-�2I e*�'V�HQ���<�����G�I`�2
v�<��9<��f��Sm`���Q�����,I4hC�o���� q�Jй�O9���2@�ǏI�]_^���VGr��3�R�R��`�;�!#_a{{���>T��\��ELaV9�Pg5������	��Q��K �Z�Y�1+T1W���`�0�0����cΩ2HA�(T�a� 5	�co�%T�1DX��)�GQ�r	�&n���9�iccM�=y*��ޢ
��
60�;�ꋄ�3�4�8 x�V&nm>~�Tnܸ!���\}�U	���ؘ�ΝK�7������ex�t<e�aI�K�yj.�*�8T\C�����kW�kr�����[o1趟夘��۫��2�bڬ<~�@���G������sY_Y�%L���_G��DXE��Jn޺.7o�&W�\���eV�|�~�s���B,$@�5��N��B��	��:��gO���J$Jװ��1w�ɓGr��wr�|_�_��a�a�U���+��2��M�뇝�m�\_��?����d2>��@�~��
�E�H����� $@�5He}5�Q�)I2(z��� �B!�(�c,0����\�1���2�ٟ�"s�{('�Ƕ�4CC�4�	�r2�a��!z}���0�D����9��sAl��)LB�� 6x̅z���#�\�wD[�ȓ2�9=Q��۞b�s�l�}XC���G%������bY3�*=�N��{ؘm��������j*�5����Md�U����t%��p���M����D|мZ�q�u^�Y*$��w�=7��*�B��Jh�5֏���F��A_cd�-Q��!yٕ5��W�Q�T�Rq�M�>a�JlTl&��Ǆ;���,�*{=��G�H3��ʈ�8��|H ��~�5��5�@24J��ު��Q�c:��̩�����Ȅ����ƭs��d��kDAk����~������(�IU�RQ��*C����eｿm������I���r@"A�"�%kL����gy�d�#Z�-S�( ����:ή�o�9�ɳ���������=�{�����s���r�s���l6f�VT��3����B�� 
Fh�&5UT�P�״=YI��1'�R*<�LVz��GGGv|���g
FO�öZn�Z,yI�+;���m��g��RKo�Ȧ�Ԍyֹ�WF��~���1E�L��Ӽ'���)�#ڶkhC�І�]j2��mhC�V6��4E��6*2Uy�A0%��{����Հ9U[����f	�҃>Ŗy�����5e�c���U�]�Jn����6�R�Q�༦T����g&���L�Π��e���r�ln?\� �B��g�� Է^�}��D��-J<&Vp� Y���~ZI�,����}��تDp,�Duద�~PmTL�o�AK�&^��=��lnq#��A= �
�ܾa�Y٨�ЊU�|K%P�ܴ̣@�o��^��|�M���-
s'�O:��&p+e%s���1�m���dO��b�V�x�&�?�⥢�@hZO!� ��"�:Q�n	϶RU��2dl^�l	�����w��&:��P�4^X�c���Ly!�א��ȳ{#U%�Na��J�M�Т��v.��2U�ү=�{>W>��^�yi�}m���C��ܖ��2ڲ0ǥUe=�A�<y�L�ٵ -�R9 !ƪ��W{������6^�r�g���3�2�/�����J1? ��#U�z��챺�Lܾ-�R�o�K}��9����"� �>|����?���Hj�Ϟ�?����������*X�#c��@���<Ǩk���$`5g<�5��KfM�N�8k�;_�!�z`� x]PK3';e��c�sV��ν땷���9������G?������<1�A9�[�T���K�^������򒟵X\�H[W+�ˤr�mD�`���8�/������ߓ�8:��qg��g��m�s��1�H�Y(�1y���j_|�9��~��-��׾|�Ҟ<zl/^>���s[\^t�d���2��]��٭[w���VS)mg�I���gl�X�e8���^��Y ň��	"B'@�Wg�ϫ.���|��\٢�d��C8�,�$LQ�]d�D� 0��7n1�j��0�h x���OC���./��B3�	y&�	�L[�γ$̾�j��I1��x*9�w#����1�p���=�@��ʙn��X���>e>�B�9>�#(�p=D%=,���,d���W&� o�N=l���W-,�>�F���:�/H'�@�Vnef�de F�@��w�Q������~����"�]���	FX�Sn���q�dN��3c��N��+x�ؒ�B׮>3�4&�3�I�5��x
�g�'��Z1����t2c'�#Q88��EX�"�r'DGTa����IR���rB�n�~��J��	?�r}�{.߯��-/�HAhx�b�KX#�0a���t��}���Nt���J�V�s6RJ����M��9�j��YY���hR�	����|�S��m�5L"��I��������������6W�c[��"+U�^�{(��O��-q���
�,����KG��v�捰����)|m����������S)7�NJ�ZV�ڙ�E�����'�=���T�$NR֮�I�!��t��i��$"�Cc�X`5��mhC�.�� �І6��}kZ�P=	OA%����N��x�C(���h!`��wR� o���� (�D���m[���VX�W���?�*ɦf%$}�+W.�|�
��j<H_5-_F���>��!o ?&NT�1d�?�K��,�Fe(�����nmŗE5�5�dk3Փ7��m�۽�m�EUI�	�x<�����C�բ�=�/��u�
?ձ_��\��������P�k�ъ;���?@ S�w�!�V����6��Q��C ��goL`M����)�Qx*�-�j�X9n�rȫeR�t�.�����=Tx�b�4e���hwk|�<�DX�:yA�K�vq����0o�`9	s�.��C}���#��g������Zy��{t?��HLƐy�oĴ����+T�����F�S�
nW�@HD�HS��鉽~����2��%���
�y�*м��k�v��V�bu�{�K���_m�@��9>��9�kC_=�ڬ\����J�?J��T�уJa�BR�0� �[�xP+��ն�� �'�d��j?|@�ãC��'��_��?���¿����?��������fϟ��
��/�4��Z	�,�4H��dfgg���=���d9���Я�Ǧ
c<�l43_$Ε�A�RLU��-U�
�x&{S��:'H��t�����_|�? �1�ޣ��mr�p, 0@|��������p"y��paA�E`�~�nqC�)|��g�����ۋ����ȯ��+���*��/�?�H�
��@nY��s^�xn_�=z�-�W���T�L�{|�y�ߗ/^���R�,y���Z�;����� (�]PW�r^J"T2�Pyp�->��k�����g�_�(�e"��qC�S�h�Z��W��=0q+B����&��� t�J���MY�ޒ���5�ػ�o���'��O>�;w�0+�;�1쁾��s�x�SU��B?�.���IA��..N���+{���c��@?� A���Sߧݪ���?#��iON���h�TmJ~�:ºaz8&(������{�~8��߮չ��g��p��ID�W#uR|���N�zM{�	z��\�q���9�{�	�=�[Wy1Ȯ�@6���\�9eY$�2e�ȃu�PI�[2����p� Nt_T@��ґ����I�vN�s�Mr��FI���������J�W^[]�k�>���o�'n5�&�m)7�9�)�ت}EnJ����A0�Ҹ�h�f=Y%���O�U�P��<�S�1���dX�IEU�u�ޯ�=ؼ��0��i�,,�5b��m�)�Zof���I9	�x�z��m��p^ P�2�Ov�A��s�Ҭ�m�;�|�e��¿m���R��7I-��TELPT��"�E؏�DMm�z�|�c;W���DFT�?�R�Vn����x-"�EFm�gi��U��	Tl��X�eg�%<���І6����dhC�І�-j#F|G:�T�ʉ$��#d�
����_�Y%�'X�4��1[�G�l � ��O��-�@���|��# �ne�+�8YW����-��&*�)Z>؍n* �� F���Hݪ���N�+x��k��bǞe�nʳ<��-	2��r� �sIy ��8w�h���e�V��3�ޔ����$H�G���u���s:���g�����7E����QI*�H��n�$m����*K��
L+�
>����t��Z�E"��Ҥ�H1�f3����-��8û��lw?g�|������0O >)� �bވ�R���� �+�D�jb�v�A���b�
�L�#�{k"c:٧�m�1� �z��.��:�C��k��� Z�����겦� �b���FT'LI�,��A� g)5BL3U~��������Q]Ϗg׫`oζ^�ny�sص(��:�\���t;�]�VjL�U�wS�"���nְ�WFG'?�)�V`��7�yUj�*��xX%��I�N2
�qg�%���O�'?��ȕ0�7n޶����)acra�od��ь����	�n͕ ��b����k@ek7�u������nT�\��Cx_o��y�J"P��?�mڒ���sxx�>��c���d��K���� �VQ�>�����w�������HA8������B(u  ~I�"����<�{���.�.� ��j_ȭl�����9I�a�C�uJ�J^ !�0OWW$8vE�+�d`�tq���$��N�0؋G�D�,���WV�V�.]m��|L����vx|l�<|�6�u������~�����}Ü�Ґ/�%kS�S�3V�AT��"��'��|2f��9%ყanܸ{�>��ٿ���n|��^I3�}��a����+���Iz94��U� ��� 3	�xm��*r�g����/��O?�����d��|:�㧭��Rs�G��ߥ
@r �űE���E	��BߣA��}CA�8�w?x?�Әs)����g]�b4�a����ެ�7)70I����0������J��s�k4�bv%��
um�O�{���27�����TV$\'�koeͅ9�Z��O�b�����
�o��~��OI*��`�G�ləƳQ"�an'I�O���A$֖�0����� H��F���W1�e]�jͮ��t�m!H�\DI�.�*�W�d������DM-p��toF2s�j{?�LR��y�(&�����D�#_�h��쮂�4�QQ�9X$"�r��"� E^��:�M���zf���ч�avI��h��$��c?�2Yx%P��bW�ຏ���l�H n�{�M�"����&�H����2��ԯ�R�eM�{��m��7��rb(�~�ڊ6c]�xӽ�x��o:(>]�t�mhC�о{m @�6��mhߪe�=�/��#,���媎n� �s�FW�IidC[�M�e�J���@t���R��QA��ZxY�E��>��uLWl�{���\9��K�R҄,�� 3*�s���7+sV��e���g"��Qy����
�F���`�7�YR��B��E>��c�+?��P�T���G���Й�-	ţ��y���{xX��.}� !�I��L��\D�d�~P�])��Ѣc۷<wu��gG�zt< �i��&���y�c�����fջʈ��d�J�U�`?@@�| �2�5�����ݪem�>�΢��R�,���T���[����8�mc�*M��o�gd�eB3u��vU����n�b�iz5H���|��L`�^6"�,Pix2�hF�'�D��?�|�Q@���=I�;+�A� �߰�1�,b*�afQ�uj˫K;?=�w��NY�sT~���)]����i��hQ��4�NJ S�y�= �N#�E����(F5���X���m<07��WR
6$�د�W;�M����ƕT"�`ͅc�t����l�����-V`����?8������/��?��@�f�4��݋��(m��@�j��
�G�,�I �]F�݄>kD�t��I
����Cb�,%�4
@9W�i'�,����w�G?���$�yp�]� �R�hdF`5��//��/��_���������Kz��$W�:'$v`�؄�V:)�C�Z+��c[��vyU����Υ���l�0J�1�� �hҫ9ˊ��z���[�Jj�����B].���G���[���@�U��m����׳�O���mQ�\�*ԱN�֦�};�q��?X���%��A��{@�ұ���-�%$k�7�Qn.�XTsG�p�oc�]�|�~��_ڟ����w��X���1��;)���8�1�~�UF�7H����PnM>~8T�'O������@8?�	�_��$&[�[�X����8��B�](�Y���I�����p�TT#t"<q����v��m�̦R>p�Km�d;���~���rWL4Y�*��-��^a�Cm�f�qE�����u�I���vM�I�W�3 :�w�R�ݪ����ߤ@ ��1���D�V��Mt��%���d&[\/Xc ��1��380�7��&*�Ҩ*�6�H:Y�v[�GO�58��3&*�s�MB���A�� u� ���S�	�M%�J�z�9�;�q��V��D�9T\�t���L��J$/�/���	=��q"��dRA�npgȠ�B˸߁��}�_<��R���hn]�yT�8uCMc��,�
?�\eCi5��:$=����X��6`U��,Ψ��9�n���{O���P0'����Xg��Ʀy���N��~�FŔ� �h)���,X��i�ԭ�Z#�HQu�s��W��R��e���q-;y�9������(�=`�{C�XsV%��C��fehC�І�h2��mhC�ִ���Q��9<ˏ�@���D>� 6ƕw>�;�����Cs��y���Y�
sY~$1��I���J^U���6��������jB�ɆH�Xi�V��R#����L�W C����K����_kQu�5�B%6��bi2�1��!XI�"���6^�.`;���`l���H	�o鱬r=,�[�H�a�ȧ�>ē����2�;M6_[�%*`l�2�D,��C��d�ho	����h�^�]DUsN ��O����e�4��V�e8��`!�����C&�iψ�m�fL��9�5�y~B����&/k�/�hRV*�2�i8 W �����
d]�*iS�F����͘?����x,�d�B����H��l
�ME&�g,����k��O&n#%ࣃ}G��Fk�b��g���e���R�T��i<a\"������$�%a�=�47�}	Z�W��j�]�	(�Z��j��bwj۷@����s��A�^�J�Ď�j?j7��٦۵����������|����w��d2b��4 ��Q���[������C�̈�x�׸�sY��Lm`�'P��HID�#�Gq�����JU 5��:p�WI��8)�lU�ttl}�1m�������[LTq��x6�]�f����S������������	4���Qݻ^.��r�_�D��p�2L�T���ͱ����*�I�Q���k��>��޾�^o��C ��|����Pnܖ{O6�:��� _$�����'o^��Ǐ���t��c1��O
^�qk��v�~8V�B�����'k^���07��µ0�VVX�U׀[N%�gq�ބcG�m�`�� ZƩ
k\3������}�1|���1�c�| �C>��� �.К��`�$$��Ts��d�Y\!�IU�Rg�re����\�jI��h�����Bk���f��F�Sae�R�#����j�T�׍�w ���YO^HmZ��@{@y �������ګ>��b�.��`�kj����@�`�TM�g$Q��IM����?���|-�2��O���ޤPk`>`mTU׫0�=3t�>�$�^I�j� ��+�6M������T����x��Xpp�� ��o-�R�sow��c�{+ �JH�hY�s.H@��\ɻ�%��������>��G�4��"Q���bx;�"�0�zI�����J�Ϥ<�8�Q�VB��k�*��O=_�ZW[��m��V�2ja
��]��J�H6I"҉Y\ �@(��-�"q��(iT�����MvT����zC�2x
���~�c�������#���Nƺ��+��؈x`AS��1ȣ�7�Γ|qe�ߛr�����V����μ;��Ś�Qa��0����l:�ٺ[�n��0@dC�І�]l��>��mhC��4<��la���1��6u�W������9� ��� ��v;!����e�{�<���p�
����a�C낲��x���y���h��2T}�zL������/ �$-�&��D'H�\�"�����4��������q^�i�)�*;�
�T�d,�?��� �A(�K"@�cIb~�����%���њÉ�,�1F^!)��ڤɘ��4	c6Aut��]���^���G��=X>�>D����mR��0�kC�}��6�j"3��+�Q��a��rÇ�	<�6ږ�)a�J;�2.z �����`Ֆ�b`�I�r/�%r*Wt��d�B��FG���+��T� d�A�uG+1Z�0󹂂�V_��e�q�5ENUԊ7]X�t�@渥Z�x  ��IDAT��>�媤��XS��q����}㻊?O<o}��I���KYn�9g�|�1s���-�V�~<�W~8�*���;ٰ��X˅���h@v�q8�2��b��#dy���'��e�Ω�М�l�X��}FR 
��+�_���վ>�7o����{T��\w�e	A��+9�i�*�<n҆�����XM#�,�'�o�5����( CU�ɹ�@����l2��v�}��}��*@�.@TL��?CV���죏��N޼��ϟ����r��^���N�H�Q P��^��h�s��U]���\8�cO�	����z���T+����\�E�=���n޼a�����W����܎�o����I��T�8��������o~þ�|�:U�z'0׉V�B�p�$w��'7XU�*�?��mք�:�N׆�{$ѡ^ 	�(㣮 ��Yٌ�^\^pl
V��X^�>��{].u�k��əo5ɚ��L�OP�`R^-.�ի�a��q�'�<���a9G5X��,�eVF�s/�]Z�Z1��8?U�v&u��"�P�;3c����<�/�̠���4"m'#�?Pl��:9>�i�s엟������º8��0�0�X��Y[6��sr~F˞���Ǭ!A�{�|���8aCa�[�1l�6���W
��m`�y�[8!�|�kXC��i�� k����r׀�PJP�h?�?�U���!�I�a�� #�-߸~�������{(Id�F�A�چ�ץ_�[Z��+%�WW������t�H�G��\]" }B�ss���#�o��̏�u��v\�{IptR�����EU�Pu�Ju������ݺu��E���0�_���9��_1�����ka)ظ�U1�kRbC�H-����?-�ʢ}U�ʤ��de��HQ8I���5B� ��3Fxk}���{1��AJ1 ��1�O֒����=��s`NoVU�Fnx�Q%�\d-�'\')��l$�z�:�G�]��WX�I��(1���}��jt�[Z��NLE�FR���Vc�ϋt��h^�7����-�t�wp0w�3�u�5�OLy��u3t��(=�0�x�M�{K(��`Y�sUR�\��;�Pe��sm��f`�N�{!���j�V0�W|�ј��J�s`ڮ��s;:�c�	��g��Qz�ާ�_�omhC�����dhC�І��iIUuI�ѩ�S�@�Gx0�P���	xG�r�j������"��K�n�3�.�*0�/_�CT�W��	8�b�l��C�V�mn� R��1��o�
]���:���\���U��@G� �����c��>�g���(A��-��:�?�߳P����j�cz�)x�-2�w��G$[ V]�����6�\������SV *'z�7$ui���(����A����0n���H&�m��H%��=�������<��n�I��2MrYe+�vIR�եE�s,fD�+eũw�*/+��i+E*Q!Q6)�7f�kB0��ue8 "��%���#�}c�]J�B��ڭ<�"��0t�X��d5�`����ã0�`�m��YI�kJT�b�T��GT��#yCAl���2��cil2��|����7����|���.�(� �e"GЛ �Рf�8텯;�q�@9����1�jrx�7�-�����v�L��/(/eD��B�Qş� :�/7�����us]��v���U�܇e����h�Q�k�v7�NPoܛdi�k�3�E�5� [֌��6(��{e��x[V:��y��=x�.�«����4w���
v%��i�R1�f�0��Vx����.��S��ɮ��̲�9�N�̢(�7�r(�U��D$#�����w��>�s�����nݼKBz�)I,��3Α�>���������~�w�������о��J�:� �b)�7f� w��ma��l��z T�G��an�u?���$a��xƘ�l���w���i_�M����H�qOf���r�� ���{>}B��G�O�����,T��y�g{s| �a��_ϟ<����R����`�{���a�I'L��嶅�ID<%NAL$a����s�n��}�����{���H�eP2B�f�E����c���$�zݏ�D4@b��,�Ξ=D �ȯ\�P��k�]ai<#*:��@۳h�j��es*�P��D`�SVy�	 Tw!s�a?;:8dQ��<O"�߸��?��!�N9E��%;�x͠z$����7X]%G�5�6폧W�`�F�ְ�9��U&a/�eUD�d��4����R1��V}F�O���R����d��	?�>��C��ݼyS�
�դt�a�H��iO����8�d�p�Q}�f�0$�3������~�,�`0@ݳO"`As
� �'
��[P��s��B�Cm�a�G��=�l����4������Rl��VTY�����'Ң�\��X/������g�x�=l��!ګ��{�8�4[ڧB��/�q�s������v���`�a����񳑵�Xx�
�\ɵ
�9Iт�cF�f��Lg'�D�aO['��j�������b�v��kj����O�{���$;��t�U|�O;��ʕT�qx�m��fhC�І��j2��mhC��4<���v?</��:m�ީ�V%�����l�w��}�t�}��b��Y1FGx��rV�Ã����g p�^��ĭjAnch���V��42��-�b�*���P����0D��`v�:T(��n��=�E� �OY�/5Ƶ��V$Σ��ႍJQQ��lN��,@�h�C�aI�E��xh���-��-�^�J�"c������4�r�!8����K�*�;}�fr$k����H5 O1�E���̉i{I�ޫZ_��P���Bȯ�"GSU�-��h���}��w-� �6��XMLU�M�G3�G쇖Rn��;z��5��oǍ��l�c���h9E �V`�N@h���mL�E�*_|& ����:P[W��rg"� ����� �l���8ه�P���,�L'n%��Z�9���N�EA�,q���+b0|������������À�{PE
2��~G�.*�q~ e� OX�M*'I
��(P_�* 5�l/�ى����hM;ˢݛ���.�	b�mY�=IJU�@����2����-��y�� ��R��[�Wj��ɳ�;����1���fs�1�?Pe���V��je��KynX��Ԋ�ݽw�������}��8|�t���ɣO��?,W\�����zI2���̭�Z~����}�'��?�S��;wC?da]i�������������뿱����ڬ��-��6\�f���%%IH�	E��h��P�x�B�=�������.�DV^�l^�j�<9j�����h�l۸?^�=�}����G$���M��ʅ�п��K{��9I,��,�Q��e�@��2*B�&Dҍ�{��+ZGa���z,�6_��e��@kw^�I�������M�^v���v��}{��];:�ɹ�0'F�Rh���B����NN�>���]�P���IUUm�TZ��¡��cD��)�K���4n��p��^�G�>�a&՘���^��I����T�0��Z�ʾ٘�^o��y�8�ef_H����fK���ΐp�%+����{3K���dm���X/�-@K���EtI���]U�Q_8B`�Ϭj��%e�F���Ƚ����<|�>����~�\0I �i����ř�������ۨ��<C,Iܒi��ю��?�K{+�8���$� ^�� ���#aZ!�d�5��M6kZ�y��UY3�\���[�N�k�!���j���x�����S�#�@�q��F���TJ��fN+��L��3*�T<"�P��8��/(��'5~��q�؟ʺ���՗ʏk�L�=�P�;�ݦ�_U�"\��j��9+���=ޏ~\��J�0�&���(vB�F����e���)�(^/m�c�j�ڨ�dݨ{{�i��BЩ�
}��Z�כ����VkhC�І��j2��mhC�ִboZ'���q�	��x\4�4�:a�a�皚U�IxX�+�i�P��(K��U5d��*0=��<�z�F�t���s�1��C��;��3>���5[��TU\�m�	M�
��I�Зf��eY�H`���� ���ݸ�q�C�xv	^[{�i�]f`�mzPV�� V��2h�yh6�пi���B
��@EΊ稦��	l�=A}��T��VU �XU��;��T3"����M����$&M���v~]w=+���ތ�
��f��j#	j��i�8i��`���f9BP� �	�A�����s��5�s��z����\�!͎�G>�s9�$ې#{��VɈ�m�[�U�*@�v�� �"��Bڰ�X�7}5,���5>)��EV����� ��1��]�Қ
T��7�1��w��$���47���l��� =�R��w ,�P@��ɟ���ſ��ݻ�����D)7 ��z���]]]�����T*��X�}%�����S�y|��B���w��L����6p5�6�6� ��Y�ʅ�3wg'Lԧ�V� �0��c��������V�V6��6[�k�M1����-{���Я/�?�r��T�[=���N�.��ͣ#��{�n�s��]��*��
@Dx�w ˖a>,�����0�c~]㠠�I@��پݺ}��N�g����ܖ+���������������s��_��~�������Of\$�s�5���$Y� � ,��wbo�Sْ�]���;���w����4�$6��׍h7�!I,s�ݘ��H#�w	�U����w�#H\drp��y� �T�j3e^�xiώ�Pفk�����2��� {S�jwC��ئ��n�@�0�eӳ��4�!lf֋���V~K����=�  �������g�"6�����6	c7��o���9Z���6��*��7�_ګO���r���)�-mzhQ����lF{_Ǭ)�2�x��h}�ώ��h�� g_Z�̮�^G Ԉ&Ċv�5�4*Ұ�f��a��sP�W�����.��룫9���n���j�y'�P���j�%���X���;�7���k���DJѭt���Z�29�:�Ŝ�\�N�����s�ޤ��������X`�ymYs.q_L;�|Ϛ���]��t;`t��g�j�x�ʯ���zP���b忹V�$��N�Td[�g;W�q�Τj�"	$��J�������!�R)�E���+Ϥ2�V��OH�l�����s�WU������ՀvV^�k98T�R���/ԪP�ẋ9�7�I���O_~?��z��Jhm9���6�ggo8����������E�^��*�َ7�NA��>����-�P	�>���7ծꀸWG/�I�}�[Y�����
Rޫk�'�'nhװ`��NAII���mhC�w��І6���[��*�n�v�U��*<��YZ��R��h��N��G�*�beZ�FÃ�9����#pl�U��@|�ǭ�|Q�9F�z�V1@�*qN�}F籴ۊS4X3�w)Nj�"���˨b`e�Ŋ�p.N�D{'��[���V$@"8 �'�Rّ:!�c�ĐgGa�h�6�
�^�A|�de��7��7�b��=4�vQ�Cꁜ�˜�C0�ƠU6Hl9+&�y],��G�Ɗ?���=k{�l"����O��G�e��.\s��^��}G>VH�|��F�_�*��n�^��E���oڽ���+ ϩ�b�=Pu%țٟ���YoV��e��]Z�4" �� �z�q�h 4���+mId�.vE�5�z��F�2��	H��[���p� ��[)�hZ�Ţ���c���@ ��Qd�0��m��B�2����/f�9�������?�O���ه?�K���d��
���뗴K�Z���L�74�����Ϥn�����O&{}Pl�y"�4�$� �a�uRy #$��'B%����)�<`�6R^UJ���zے>x~�KR�u��|I'P	 ;@�������F<'�s�f$�����n޺k8���vzrª��,�R�&���Ν�v��=�q�-�F���>ׯ�Γ�mm�X��ى]^��eY�<�l$�ySU���{��`�<�w�� |�έ��21l�����}���=��+[,/�6`��V�M=�$�a�J{4�0	��`��ł�JE�v�ѭg�mA9f�@���P7"w2�¸��ۄq)��Py��h#�ŵÌU�o�Z�#sY����à:�������"�e�Ϩ�::����4<�Dv<M����
m�w`�a/z��M؇$� r�v*�Un+����rq:ݳ��#�q�ݼy���"|�8�g�i̤:q�?B֫�8@~�|�ܞ=���?���^��2�d/&�v�E2�M�_��9] ���}���߉F��H�2�`(�s9��,�h����i�[1�4N1S�Ĝ�U�L�Ԋ<A�po�R�bo��\a��VA���/\'1��m�@
c�q�4Y	�0XQ&��˷���@̀uKD�����(�)qp�-#��������4��A�]�-�!yB�4.d�О���**v[�6qM�<�{�&ZH��|.�=���#�����S�C���{���;�}T1 ��:��.�Y��N�/r���IMź�@ �k��ĵ��T�B�-�)���p�E>�����*�Q�Y�Q�E���|>U�-�Z�/g�[���#��&�)�_/�X�B�ͳ=��slV�R�~��R^J���6]cWMo�>�w$�R����l>��	#�-�̨��Uj禒�p29����p�y�QA�Fn
3�֫pl�,�h�D+��u��V�z �3)g��sk-�ڌ&9�Ip�K�WK�'��%�b����Q�2���x"6����xhC�І�]i2��mhC�ִ[{��y�^^.�W����j뺩�M[W�j���.�F词bU�_�v�\��K@�#�C7��p L�N&@#khW�5����=���=� $A'[`�O=��Uߣ�Bf����N�&�Z���>����5V�o$H�om�ZO(��h�Ee�i��Ђ$��Ў`���[Ŭ3�v?u'X ��a\hw���Aډx���k����R��GT�D�#�<o�mWٰjS:����?w�0u���{��e�$}�p|���y��x�
P�~Я����`��Q'��]t����QM��;��Z��aNh!^���eM�U�S��1G@���k0�n����7�$Ƿ ���U,��|�4m֕�����-��G�sZ.�>W�E_5�9���c@�*�젯7�vRW�TN����F�Їm8>U�L�g�]'V��ton�G6������(��x�>F5:~xxl?���?�����-EE��ȭ+2�2N���̾��K�����0�¨��K�����gN>�劊'Tӎ���U�r	�]f�/��'�L��;H��q��9��A���I+Y�l}��ϣ��H��;�P�9�����+;;;�
��=�-G6���ۛٽ��J��}��Y蟥B��#`)���own�&�}��];�y�o�q[�*s�`�9H����@���S[,�n���MM��G`���Y��y���{�����S�&$VPџ��]U���x����z�ߛ�r�o���Q5���g?W[�s���sg�V6��ΚuI�t��	�8W�E�)�֡�������pl,�˚�6�-��I>O�"�@�)���a1�]`��曉�� h������w�	Ȉ�� �NY�^o���D8,w���k�xdr$��������7�mR䶸���z�ϻ��hK��$������?�g�5���jX���r�u�[���/;�8����x��-.�	Tbo�5��Ȫw��ɣל�il�	 �9_�8ĪX�׭�@q5Y�`sB�Pw�JJ�;�mXaB�B;Ǆ�C��Litco�Nǽ�6o(*5�>��q��|g�a�[��E$������ܢ"S�G#�FF��H��߉zi��?mX�f��j�Y��1�$����I4(�TЀ�Wɖ��*��\��;���{~��2Nn�$��+������&U	���.��8�����^�����ڽ`�kX����(�}�����F�x-9~O�9���U~�TF�EjA쭴�k[Y�uFk��=�DU)���vs&ڰ/�ς�yJ��T���m�p��Z��d��,���y:�Z��e�ݶ��R6IJ5G��yT��H�5U$I��r6�S�3N���{:�rA�܊�#ᓑ���8���`��	�N��py��͍Um[�|�
����a_�Z��/���haD+������a��ϗeT�6n�d���oT$SZ��Ǉ"	*�<��?�/*A��Vp�ҷVC�І6��D��mhCڷ�u���EU��ͪ�|5H���ݔ�{��RK�E5 #1��ß9�Oω~ � 31���롴��74>䵭���&:����y��Si�I�m�b����I�^� ��)r���@e��S�������Y<p�K""l���M
���צ^q��ƃ���A�^	�)j[U��@�ڪ�I��fo[*� L���!#�>8:�[9��׺IP�w��KJ?��p��M<�n��7+S�؟j�+xHgcVZv�c���{'�K"0Y�$sK�$q �����p,PXLaAt�`�ѫ���YN ��T ��z ��B����s$�Xuچ�x%m�Wd��"�wzzn�_[��m6�(�����LU�W��)״��54  Q[E�?�����3����w�s�s��7�vr���	���; >P��o�<��w���۷i�3���oV�u��G6�` ~?�؇�����I8�d\D� ����#����G�����=}��va�����B�z&{�i��u�'�`neCp���;�ʽ��n���q�9;��Õ:i�6�B�
.T�וsQ�*����i��u;�N�u�\�����|��^�x���0�a��?P��W�I�V!	���|ng���E��;A
�m�ycr�wd��#;<8����M�f\��a3�k����zig''����0�^QY�BeA��c �}��=|�]{'��}����x�G��Pc�J<�oN^3K�sa�8�[������^�{S��u�J�a�
���q��r]�FU6~��k>��J���,��b"��׵���	���.*��7�w���s��J�y+��]��u����%�'���u	�s*I��˕=y��!�
rL"D$w)H�q��t�����F
�x�2v�h�� xغ�Q�	�.O���س�:�]�"�1��Ϋ3���J�\2���gḿ�������	{r5P�� s�p��A<�Lc�>ڪ� �J����W�I�� �2�9ި���#�~Jd���\�̦М$���r�C>���c'��D�uo�u؇Ѫ
�˭6[ψ���o���N��K{��_��6BRSe�w���_���<����j��%L�qB:!��pM'��, ΰb�|*5HI�"�3ΟU�-������0*�B�C�RW��;�. T�z`����7�4��{�	T^�\����_4Oe��R��B�iPy͢*�����[� S�F�UP* ���"f��>�+IN4�x_�$��[Q��me�/�掻~��X.�m��0�$��cq��/�	�Ӹ"�7t֟K�6ۛ��9q\L�z�Q�IU��*-����B���$��2cN�Ҭ��ڸ*�u0߷�����) �]�,� �����9�3��H�FJQ���T.�y}��}ۄ�����.�/8@�߸q�>����)��k�����>jx�����e:���.�5�,����<�Xj�ue���~>��mh��6 C�І6�oMK�U�O�<m�"<�]'dqT���x-<��၇b�*NY��`��<��X���tOV���@�
M������A� I V��@Rg��+��|�m��
?����S�<�<��H��ٵ\S�t�� � ��\(CZ��[�/�"���#oi� �p�o��牬�<YU�컆�����,b��K F��hly_���[��E�E$Q�( -Ow*<[=$�{�H������I���"�E im��e`���ϳ�W4nك����dP�L�����
O���-�-8��� ��0쮑h�W ����y^����8�90NХn� x|�t2!� ���û�O7�h:ao� �eI9O<�~� �� �1'�
9X�Z2_�_��_���?g�7=��9I|������G?�����vpp@����7��|��!�GO��7�|�� �s��=/*����<x`~��ݾ)��t6NP��&w��Jc5�x2c\�,�0.� M���4K{���}��Wvyz�
ObAI�|t�Ihٓt�T�Xm�
�6�����_���*`7��T��^o�s��_Ӟ,-
U�b���y5|m�2�~eS��=�����J��Mlj;;��xb�^����Θˀ1� D��]�;��E��&�=;>��y���pAU�|�>k���S)��R���d	�m�U��-�.l}����%��}��� �э#�<x�]���Z�!W H,����iG5�2�{�v��h�|��@�(+l��P�V��=�+o�H��T�����^�¿Oޜ����*[�����1�D�[��R]���e��'�P�Z���EfΈvQ�_aagn�չeO�i~���a��S}@;�����a���\��ZEj��^�ze��eOU�e�� �W���֭^��R��YO���:�q�|Tʷ^-�
�D@;�^�T�X��+lr�5Lmdk'�(e	�ź�8{ų'���#{��-�/�V̖(��-����7$�i�� �jWG�t�HYQuNDt�w	�̭�E���5"� '��l���g��L�:�0F˿���Hj��N�Rإx�8��GO}/��M�p9n6R��Z�:�b���=n܍4wr�8a׀-e�tl;��l)�õ*�RW�`�IzR�痈| PNr=��P� 0l3��Y!�_�<��3�P��r5ѵ�'aJN�+�c �-��jNZ�� !P^G��]z�V�&K2��Ի�������D��Tc�����	�x-�O�}���}�j2�l�G�"7IE��ϊt�
/�|N=�j?XB��X�!e�����s���NV^�`�u��:�?�15�a�R��G*��l��
N�&N֢��i��b°Q]�x��^yqy��#���p̘KǇǾ�l���^sJ_�|�rF
�O딑�{�gϞ�>�N�V�h����0���_�=}q���D��;�y����u�X�ט���[m�s� [�ύ��ދ�%����%n}�㚬�dK\~�.XC�І��l2��mhC��4<K��Yx����0�$O��IS���$">�`�J��rI�K�l:z3S��)�J�*�:�r�Z^�E�?4�.�APl��E��=�� �G�x����@J���"8�h;��m��KV�6^��L�F  Wx��qm�a� |���A��tq�
M4��}����ai5�0? ��x�_�K�&��	�<�'�z�8B��L厰���
�IF9V�#�H�+Ws?+��I���<���or�N��~��5WǨ��	<�A���LZY	VP���Z��l��gP8*�B9V���T�p,MY\Uz���x`'�T6���l�����B�=�����ԭk�Ð����H`�zY�^�R���p�
�@�@Q�&�����۝{�o-@�پy�����H� ����� tsuq���XQ���j�՚�6�y?;<�O>����_��}��G`e�YP��2������H��EՕ�������"o�n	xGe��W��8������3-6 �����ɛp��ɋW<~|~AE͈s� &@3 K�����|J5�s�`�oW�2������T[�R�j}<\%@�f��X6YJ�I�č�^���]�nWq?A<���V$n�eFXk�3�~�f�/��������&g��?n�=bc�E��_Vk���l�s ��e�4���\H��z���%Ʉ?�Z�LBf�� X�\�jq�|��?��޼|e��V-?g��v|��ݼ���'��ܣ�ԕ� �"���@����k��c�����&{|?��bq������g�K�"��
X�B�߫�θGn���*7�@EXa*nPo�'�O 6֮R���YM�d���	��鱭�z aq�m��"rWܿq�R*�T�k��2� w�	ȸ٬W�R�Q��ᇉ�>m���ˎ�5�X8���=��{��/Ƴ�+_�rI6�=��J��9�^��}N�A�Z!�Nb��&���%���ۓG_��}fO�|cW�ʫ���p�����
J�vW����
qU}��Q&a����ݣs�I�Ӟ(��M�_���{�f�@�QF;!��TXմ�R&�2jI!�Z�l�Y�:�c2	��5� `���ށg=!�9|�׸ެ¼Z��
��&ܛ�8>�4a;�igEK��כ�`q��L�#s��/1�Ĝ��DN��"���F�s��"��J��T!�@�� �o��Z�`�A f�S��R���N ��Z��ޙW�D&	�r���Ϛ���V����6��0�F��/�0v��f*d�rKl���gJi�u]�~]�M9�$���'`���.7�^5�u���y�Q�Z���-�R�3�|��(�W�G�6���Y̫�i�a��`��_�;\�p��׌��[�k�]�S+Z���%J�}(��Ÿ�8tњ���a�!�й)���ḩ0���ܠ�d'��q�*Z�q��sG0}���cys�����zʾ�u։��)�H��k�Fb����T�A+D�/otu���M8g����f]�lɽ��v*�������:~xp`7o�:��m�p]��v�]��VaN
+<�W��q��"�*�&k`EE"�b��~q5.�^%�m8��RmhC�о�m @�6��mhߚ�<<�����ak:��x�.V��Մ��P�>�>7VV�j>�.y>A�rT����(R��{|_�r�Lɞ*s�dYV4}�f�E���[����EUZ{-��u�k�"��k7�W0���Ѿ��;dG��w|�ϩP��5��	�U��Ȃ��d�G�<�(sod�q�L))6��pM; �yK�� T41�<͢��L�ȿ���-�Z���[���1��	�-��7�.���=Z���
$C"2�*�_'O�Z���3N d�4qA�@�:�- �pĀ[��D��Q���Ӿ"1�
Yt�d��G �B5����F$���;ߝd[���Dq m���V,�a
���+*�����ܹ�������_M2`�C�߻o?����|l7o�b�tv`�7IAI�0b�h6߹�c�"0�m�
 ����8��U��2�Z�JYTR�/�" �1��V�g^��������?}j�^� @�
Zz����o����xcG J:�u�)���$Zr���8� fU��Xd8VK�yoj�v����Quql��H�7������<ݛ��>s�?U�\����W/����>C�Ax4c�3в(�-Z��xO�	�?"��@�Y!�@Y����V�g�N綾��W�^������˗vqq�,�Xa�}a?���;v��]�y�ܸi�7��q?��I*%M��M�Ԗ���j4ٳì��@/�8�?�J�2� ��f+<�q� @0���^�=}��9�/`M�9Ye�-+�֭��"�n�N2����ٸ�b����c~T��90���!F���z���
�q$�Y�ݰB��_%˩�q-��R�p��\Ê1mu�����~��t� ׯ�)����q�i���87�w�a�,D�����Ͽ\���I�/쏟��=}��?��N�NI8�����C�غ�"��T�w�0g�R��9��:!x�=���I�e����k�l`�q.�-��f�*�Z�I�@ł����p��b�b
E��o�{��5+�A�N�3�sa�&c�"�`<V��0/�Ǥ,㞘���%� lk��c/F�Fn�GR4\71��'(IÞ&�X�&�O�_�nmo�%ۣ�Zz�P>�r���`�t���Q��VM���Z��(�Vj�JL!�ɚ$9�׀ ���I&����\T��VVRiHe��H�����Ǣr����s�SD�0ץP��JB{4�����5nBeeHa�a�>��o��Ry��7�f���׀D���d�1�6�}[�"�iZ�ܪHP`"?����u"P���3��U�~ބ��}e�?���I�N�6�fl$1P��-앥�E�0���|/@�˘�X�3�V�����5�����#�ߍ��4V�ʢ�:�EX�X#P�����@?�.�C)��&-��|���P�� ��j���r�1��cGB)�oR�~�|,oU����mhC�w��І6���[��<i;����W�h�?�&�"9���Jxۛ�^�S��Gn;��{�4H�� `	 
�x���;�V�~	���߉T  1�`�Z�|8���/�1�s�a)�-D�:Ϸ�u��o���@r�d�p=��m�����������	:�FT�6��A����DR{���JY���x F�fg}�8���k��4 0VV�Zo#�C�F�`۵�B��sE&G�m#^N�	�YeI_��9�����`�Q.�nT�7Lg�������a��ϼ��O#����Ӡ�*��@�r@.AM��*�@�W�3�V���WG�o�DE�pxy�g���m[��q^��vR���]�%�4+Y̿N�&�9:�TU�]��6!�#�����?���w�����k���z�@ܹ�����U�W�.C�j��ѿU�C��`�S�$� �Ba£�j���!0�x�Al��h��r[���쓈l,�=+fw���'�����������>�� ��|�vVP u���X��"?�|ʬ�VQq
[U���Ү!NDP��@y�_�[ ��6�6�7��fn��u[n�)�����TE[6�29;*�w|���X�����˫�={a6����&T�c�otL�]J���Ќ'��	0������C�[V�w���7(�N^�7_�Ѿ��	�WT�0`
�|l�0wn޹mw�?�#؞!j�&���iS'���ĭ�����Û��M�&�ULy�p����Wų~N����G�t��.�����-./m�*�Jy �T���qi=��3��� ?��T

U�7^�%��Hs�����ym��;�I��$�=�As��7co�޻X-���oX�]���Vtw�ާ�H��a�!��$��im����4/#���E�%�ro{,�]C�͂��FnVvy~fO�<�̏'v��%��M�*���,&}��V*[:�ɼ@�҄���.B�����.��Ú���+�%�g{Hs�q�������ʩ��T�}6���1w=�ܲ�x��5$�q"G��'v��΃�&ә������^Ps.�I��}�l�2�O5n�(���v����K�T駠������EZ4<愱B	?`4��<�ʪЗ��|^�P$H��A��A ��5�;1�'��8�II�7�~N���
k�~���htU$�����ò�I���n��yU���S��A?7������ҭ��^̍XB]4f�s��/b�"�*܂ByE���R�*"Z��5-D�~�bmjY:�W*P�m�~�E�ԧ��$j�禼繲K~��ŕ������j��]Lº�5	��K��i�Il���G�O�+RA���9���e]۬U,�F{�2��3� ��"����R����js�R	@D�N��ÿ�Fp]�6�k�=/
i��b�M�y���s�#���ﳣ�%�߻4��D�������.�,�]IT�y_�����B+i�W��=Z�����І6��}W�@�mhC�о5-�;��'y�*�LF�"O~�n]��Ӳ��M�մh�CX�)��sv>���� ]�hܪ��~�0�����ƈ���L �I�T����PJ�\�if=���p�4Mj� HY��8��K��M~�O{K�v痪.m�FH�EX��X�ܶ��mt	��`L����
�&�Ү��ǋ�wC�pɊU�v�Ui�c�$+�S'AҴ��A��y���T6��.I,��B^��֫:�Aê���غ�,������]���g�nrV*��(�kX��: '�83}=ᓑW������$ �p�#�,0�s:zlǪ�]5�y���!���{��޳U�D`�����U�3,{2���#;>�?K*�@[�7�G t핗M��	��x��hs�zb�^������=�׎������ʫia�5���Q�/�<���Oc�We_�񏬌>8��wH3lj�s_I�C]
��H 5�]�_g���Q ��\�J{� .+����Y%�h g���{���:/�d�Y��y*@�b���́���AOU�*;�y?ص���A�b4%	��)��0�PB xq�~`�Q��vF����Yo����fE��7�^����_}�%	���s����f���?�۷�ؽ�� �?�W��j��'�Pݞt�� 8BΫVc�*�q����<��	�xܽ�Ӹu�6�:�mʸ�woۭ�w���G��a.R��;@���$؝�q�� ��d)=�	�= D6׳aHbu��A��ȷćVP��h���k�P�y�
[����7��4܏��$B��}@��y����~N��\A���,U�x���2F©?ZݔR,\���:̍E��ׯ_ۣo��Ǐ�9+�]�z��&��1���و]�u K���Z���D�lu������EX{P�aG�6��.8l����6n��qH}~4�,�"h�
��Z��i-�$�B�̑��^�ze�=��߱�y�'��	T ��j�}�8�,��B5b�l&�3X�!wFl<���NGx���u��+�o�����gp7$�#y�E�@j����!m��x���ls5vԇ��g��O���0�,l�&�L���X�
�l�P�@E.���hyf�2�r%� jP��ŀr\�j����v�����Q���~>s�n�:YH�Ty��T��9(����� a7�^����z�A�3��\E�mA�]���g�����]���[WC���	��Ev���8W̓����4|��_����B�6���>s�j�~�[�m��|�*�_�z��ZyF�{@�}��uZwe�� oT#i��x?�Ia�e\?	T�Mm}x{*e/�0d����fs��t�[�Vy^m�����I�\!ݯ�>-���n��z&��P 5�=�s[S(h( C�І��l2��mhC�ִ���e����,�h}�iwt4�$*��5~'�Vm���3Zq��]�^�5�N>ң����H���A#� U�k� �Ca��
������ &��|�U����V�r�j�����4[�Ho����{}F�ƺF2���i_ͭ*C< �z�Uॽ*%���¯2�(D�}�;	�����Ք��H�@->'� z�n�a���{���o�*�	e��CY�함Z7g�Hi����H.Э�	�ƚ% �;�E�=c� O���Y|���?	��/��WxІ������<����l���*�G��$!�%~f�[��
'��P��+QT��y��l?���RP�B�5�1�6�<�����P����Pur�{Q͌0{( h�k/�EZTP<_Xr 0����F�=����U�"�T�_�9��4���z���e��_��:5����e�5�#(�y@(|��٩�~����7������>��O���ߛ���l����Ø�*u4�8V�[�Y�s��d��R5�C� ���B���C2�:�DE�T$U�FM�$T���`�|����>�n�RӲ�]�F=���LaTǊV��*ܯ�\<�Ǐ����fm�7o�f���H�T�����jYA�N�~nu��苾Y-���}���o��x�ꙝ��x^��h��"��W#���		�HP����9\�u�9�sS9xM:��� ��;Z{�'nYH�וifNP�$	,�M��ӽ���ϼ���9�T�0�v@"���T�G�s68�!�+�"�!�Ѩ�I��o5�ҷ̴'��V������/�'ol����k{������܎n�x����'S��Y�,P��Wq�}$���ڙk���te)��r�����.�O�v.�����	���_�"j��Q��m��+Rp+#�ؘ�E�s��0�'am�_���E�-��/+�ݜ��cc̰ZW0��d7���ӗrN����b�I��f9-�0?2O��6Fx-�+�D�\�9V�>�������?ح{P���iξ����)sy �ˆ2���z���	Ƚ�ƹ,� ������u���k���a٤�N�?�Y�-I���q��{k�njHH�~��(A�'AАCC�?P Ab� �� � P�HH���=C�t�RK�r�̓������yD��y�[u)��vޛy��"��33#Al_�e�خ�NԢ����jf�E�<����]�'Z^��H��$���1Mq�5 �l�@�Ѿ��@��[@��f$f�!{aw�(]Kv��`��Z6�FvI�3;��i���IE
vàB�����nQ7���eAdqr~���uk�P���pƜ%���>���) ��^{>�>����r������3L$1Fd�u���$�RD����1�ݿ`�EgLɣ���OᰓZ�(֊��&�aa�U�[��ξ�1m�6>p�pߌvK�"H+�QcP9g����d8Y{�Y#��L[4��h�vvM�mh�{�����ό��(#
-8���Z�4���Y�+k�b�]�QiR�C	�@�a'x�_���C�o��,4�����(�ѭmmk[��w�m�ֶ���m�[��;h��s}����>�\s}Ҫ�������#�m����lr�
���;�L���}b�WΩx�R�Rj`� i�{\�rFa��x"`YJ���,� z_=${�[y�3�Ua�h^��3ZȰ��7[䱮�D��ceH1p<�dR�u��i���|_���M&����C4u���f%�zZ���ύ�!�=�v���X���SR&{�u������~�*c�h\fU}��*������$�<��abˬ#ppyNfs֩�{T��2Q�|8����K� �ǃ�	�&;y��~���d�3*7f,��J ��#��9��M]�:h-z���$A� ���}RD�e31�x@l_;��Q>��5��H��ǳ/�Ϟ}�2U�-��{V\�ŧ�ߣ����I��*������R�\h3�~wXU_Z��������M�G���5�<�QىJR��X���3���pzs>����o���3���(���?�[B3N�XXz�P��������Ϙ?�����w{8�*�G����8G�:n�b%��f��(�]�����,�(Pռ�X�oy�3s���!?v�ݨjA8�$�����#�t���	�Կ��lk��_|�%� � _����
�}�ax�=X"�e<�Z��Z��"��k�E��Q�'T��F��ׯ��>�����>�_���5�qB�2NX�����t!����<�E ���r5H�	������:���U��5�5Tğђ��}��l����a���4>�	���
��PÚ����$��ժ˱/A{_�}	$�@�����6O-{)6�y/;�o6�@���z������ b��se�Y�]d�݅s=�7�߄�u_z��{K��|?������?�zJT��j*'ٹ��t=��1�ʉc�
r����|�ߠ:�Mx�l�d%���5	2 ��+o��XQM�y�����=��sW�ǉD��9�3����u���9���d�V�����˥,@{X�.�uq^l�H	�<��3f�$p� �:U��:���l����u��㏩lB�ʻ�'�J퇏��'�G�'���ϨbAU��^k�'��/l��{��́k�/?V��O?�����4"�#4T��5S$���q����2���<OE�P�����B0�ǖe�}Z���_=�}�E���}�\���wn���p���Aϟ-�2)�jg��xm�dnE�uU�t��=����;��
F~�bQ�SI���R+RI�@ڋl�����F�`�a�:��g��D�2�-o�5���6����w��$�q�<��kÈ�ly���Mvm �OW� �_w�a&ز��,�R'R[
é��0CE���,�=3� {��"���$+����cK"@4r���{�L�-�#���=5��5��,�U(>X/c��9�;uy6�<�[��
{K�7�br)�N���4�o䓘��7���'鲂��ֶ���}��F�lmk[��־5m��s��u}�}V�����˵��2��A�./��� ����%�6dC<��%"�p�1��YDn+��RM�����';<��Rއ^���EkdF1����������}��z� �;My���%��\�������T^�d�Q�f��~穝�ȏhU��1�"�jv$&��h��!0H^���/�v��Z¯���&�"(��AG�	`X1���W���B�� g\���Ly�*O"(�!�*`4q3^ń7�͹g?�:�^�|Ê�g_}v�E���t�B_q~q		&8Տm�R��+�Gk�'�:DG,�d� g�����o_���w�b����_��?��pz�P�:
���\���_�_��'aw@E�Cx���*�seՌ�`@h:��Ba�� `��
i��� �-�;�J��]�c]����?�7��������p9կ/×_~����?[F��a�yH�P�%����" ����8�x�2����/»���p �\��?�a��T%%�/귔�@�d���`�<�{�Q����ްT�c�� ���4�w��+T$�m�XB1.~��Qi�먖�hWT�����5��ʏ����U��'u���Ӑno-s�k�AA���@%�j�+���e}/|��矇��\y��U�<�¥�x჈ʍ�~Z��s�E�[� x�@�e�����*��E�繛"���	k:�U�G����k��o����9���p���S�'�0^O���e��߿Կ��'
�O���+S�g|!عX.�o�|����
U�z���kxo�=��A�N��]�2�<[����2a8�����^޽�k��:�?�{�W�{��Qx�w�<�UH:+�e�"s�w������S왨�>ߟÛ��_��^��'��^?'�"�r:��Ã��ނ���I���=�dN��}�@��z�o^<���;�&zU�߽y����>���u �H ��-��<�W��==���Z�E�l���E��yI p�	dYsև��Ě���e��?�#�>����/��<|��/I�tN��~�����·W��Т �;�ß������Gu�~���Ić+�� �5u���)����ـ��NyE���GzNFK�6�U�b?�vCP��U�ۄA
� a��u���/R�ѿ�����>�s}�8X������hkK����ZS=��_qMY�Nf�T����U��:k2�I�a��T��̮�ّ�^_����+��Me����+�|��F>�r�
~1By;�x�wJ�h=wE�i-+^@��߉4��U=�)/r���s��X��L��+,n�ǃHd~-bGSX�o�K� �Y@��P��5E�a��w��qO�h��K(����41����F��cu �#a�?�n��-+�v؅��펽Ժc��	��P̲lV��8�>S,����Q�Q]Fgڍb��;`���>��P���.)�&�bvk[��ֶ�]k���mmk[�ִ?��?�������G�����ͻ�Y������v�;�P� Q/b�JJV�)�`�?�����YB��l� �����Z Q5&�䱗(��000�ì<��I��ycF�� ��D ��e��A�%��蛷��';d]Ů*�A^�����m�@����|�����?�=7��
�Q���G>�Qٙ/��	��=�
���b84��r�~���U���:�ޓ��� ��4��Ʉ9t�R=�솸T_:�χh<�h���\r����-��'�8X�"�\�؇��)��?��ͯ�~�}�����)7 �uS'�f��j���׹h�d�\����۔T9�����lMڭw����h_}����O����$�ȫ猪�;Tp�/��Nw����YIk2������-jN
cF����n#\ڈ?*R:U��zV�V�*M;��;o����_~^�~Y���@����v�%���\���d�ބ}�+����}��|��'���_��}�P�򓟇���?�_��*�W~KPΐ�a5?Y}�(�4�+�/�!T��n��p�ρ'���|�
��\3�S�,�mZ�N{U�<���ʋ�\��B>�C�XQ�뫯��?��~x�����0��&,*������g#?�� �ai�J�!��ٗ_��8��u��疫ԩ̜ks�����js�s��Q���so��9�>gu����T2�{��{4���1m�Ꞅ�s웇:�׳�P ������j^gI8 kUǳ�b�fU����wf@qj�mCT;����gS�`/�ܘL"��5',�����?�<L��#�[�6������R�I����M=�{��o�:y��Yx���I�ao�H�r�� VX���٬$��pz�A^�����+@�«g_��/^p��4^!̦���xq�H���P����3�(�u,^�|�}6v7�}x��E�pv�;��<���ӑ� Tb�Ù�,/�����fS����^RQb����I,�]6"0Ɓ���:gCꐮ��}��O?_���>�-ə��Z��Zk/X@���ӻ�~n��R��駟�/�:����+��B��]����JԠ<�b�"�����I^�8Y��+El��s6�������5f��m������JK#��~�ޟA� ���ɟ�/���Юe����}#���5O�9&�Ċ�1�-��	�,��{�����e�%5Y>-/!>���%�tI�R.YL��Y�]`�{S3�Inܥ8S�CG�6~���ViѬ 9��r���_pr�a�(EI��Y2\?�! |h���F~����&ar�n�ڳy����U�ɲ�@��Ҳ����\ia����uL�T̴�K6�p���0sήq�!�H�ي�p���{���H�F���[&Sfke���M�?`��cw���=���^Xlӫ�j�����mmk[��E۶��mmk[�ڷ��S~6w�8�?����7�{>�B�`��������yzs���U���5��=zn�����#����?���<X�*DA�A������� 	y�'=@��z�P�~�z̴7(�B �u�l �Zc�f���)8���*Wx��g���������x���w��y'�j���G�7Aia64xg�{���N���4����=+�g���/S�����)�����y����!�3��_ ���4��ɲ�r" ��:�
���D�\'�rO Z�-2�@C6�H!��d
�f ��
�<�S!����]���8|���p8��'O»�G�N�LQ��g %·��zoe���K���.�I�m��F"a<=, ����,�d��IR�A0��ݙ��/��������,���i�{���������T|����3�*��S���� ����5����@��t�}�����v-c�V"�u��������.\�OMm�&�3�J8?L50�9z��,��g�iu�+����W_*$��͛7����}���S�7�*�>�Z�
	�FV�p{s��٢���*kb��]��%<�~��[5�m���横j ��~�1�WV��<�3Iz�c�aF]��^�'���r��̗_|>���Y���{�O��p�4��
�n`1�����Y���s��X �/��J��Y� �؏���}���WFD��߮}��R���|��ܼއ�����	c-ж�jW�`wBs�R���܄r$�D�K��}�hx��%�X��Z���b�@�B!+3/��!
�{��e�C�� ��>�y��{��Ԯ�s �z�S����:'��
�`�,TJUG�c~�H���g(�l��__>�2ܽz>�{^=;�Oj�����u��=�MkxOڡ��c�N�k(����!���~I�<�=���b�̞������F�7�Z��,UC�d����U|�Ӌ��ExQ����?�cϿ���������u=�7Е��]����@��+,_�� )��~�T�7�ف{Mgm�F!�c�̰��t��^*�%��^D(	nC���C�D�@����Ϩ4�^�j8�}�m�L����^��솃��Y���\XA ��t�$#���("ͱΡ=�:|fgฮ�� �hi��à5K�QSd@	���8|�ŗ\��N�&�����)��;C-X?��'X�"�;���R��DVJ�#U�/��7B�6R��Ţ4ڵr�%�|���`��G�w��� +<�J�o�9��S�զg����"��dN>S�F��ߔ��Ev~�w՞(�ȞWʄ���M����%�:�hZ�(#@r�n�oW���� |�kO�>�Yx��*�ڤ�	׏�?���ks���f��X ?��}��ZvF�j�.�}��TD������,X�$ML}�i�Z��Ge����2���g/�ܸ�8H1��
�],�)(*94��oS	����SSW����R`�/X�v(������/2�:��ֶ���m��6dk[��ֶ��j���ӏ����o��?���~}^��p����g�����7�7�X!	�	V�]e$V�(�Y�0�`j�% Q?	@��,����k*"�����`�������c��Z�A#E���iՂ��5uZ���.W��}��C�Y���B\q�-��M�0�J�C}β�jU�I�Df�My\A`8�ИR4������o��0և[ ~s�0�ǖTn�s��f<+�U;�D�*��,+������~��Ȣ�,t��rѸ��0ڋ]"N��zV	��p��a_�/ ��XHgᲘc�t}��>\���o(�{�>W(��1
\��B4��"���,l0;gv{��dV`P� PA��$��J�jfNw�9�`4^`6W��v�c8 0 X6N-��>?؄g��t!��>��~O+���6����#���Ͽ:���0��}ȴd�`�P1����m.�p�,�H��w� �$�@U�P�uP��
|���~dK��g�������E�J��9\Ƌ�]��Ǿ�{#� k% *����@`3����x�[�6,u��|�i��,��3�v	ݞ-CE��3�ӥ�x^�c����c��>|������{,�c�b��/W�/�!X����z��ZhR����YsT��r�������o���}�sΓ��/�G}T��'�� �r��wQH-ƨw��{���?և��Ǽ5k@��t���Yw��������Ë���~��Z�A�165�TXS#�@j����@�=lq�p�]%�+f����j�Su4��v�k�4I�GO�jh�\��ܞ�d�>@V1s>f���$��0��{����p�?S��i�v��Gک!��Zωy-u���T��~��V~���MB류2�^$u$j�����7���� rB�Q!� (�@�Z�uś�/�y�|�?�����x�0�]�����έ�͢e�ص��fP��AU)6���@l[��B��IY��A�D1K����1���|�k��Ae"�3b�T1�,�m@�$�����j��d��r����� KX�V�����/ڇm���3�B�Pi�G���`6D�N�h1�(��[��^�X����5RJ�|����j*;#{��I砬�8N����'��rV��RX�LQi�ڹ��o�MQE]��?&݇Mn�� �ƅ�Oɔ�2r��TA6�ň�LR�N;��ZSA��M��}��Wjɯ���֋����V01'�b��lJ�P��B%�L�6`K5�*�}�H�z��W����Mt�2H��93�x�-��2^*X�M݄5;��*R��!�*PI�	ޱ(���j{��ς�n���VD�kmG�[v���q��omk[��־Cm#@����mmkߺ�Ry����8�ߏs�~}�y��w?��?�/g<�S��F
7 �����^"���@�GuV�5�R�>�%5���6��uK�\� �%�C*�K�lV	���.\K! �^�vWٲ�J%�T���,�v\K���*�n��C����[k]����.�o�:�W(��]ߍ�0/�YH�b������^�T`�%���e#9�MF6��f��T~ ��A6��y�z�Ϧ�hhL(��>a���!����'�`DQ����EB�t����l
 Z ���-�p\]=�[ڮ]��q1��N�?n����9��I����h���FO)l��0���+/�W�
T n Y �nl0�ށ*T��&���RH�-'E��~�S���a�(f�z}
�遯�q���J�4Sᡰ�`yD�ƀ
՘��*�vtW8�P��*}KX���� �*�gڜ8($��$
^@�"�(� �����w�*P�2�@!U��䩟U%
?���=W�ú�T/[�p�Z~��d��B���nGU��-}.����3�&4���Lb ��!ڬ��B������"����J:e{��*�����7�x���#�8^�= ��Ľ���zX�K�My5 �O���찾�կh��օ���f_�D�6��тq��*6_/#�^�YdB��>m�-�˯_����d�=�l�z�^�
�6��?�a�N�Z���]��O�^����>��*v�<�[�e߈"@��B0k�BP}�;] �`f�H�2D2�5��QkU������ lbO�xºj�O��ӧ��/�7��zyJ���.�_X/P]�^@�_��-��*�Ik�(E��_L��jj�� �ҺKD������.u�S�7�p��Sx]��p����p,APbM�߯ G	Λ%T/%K�I�D�=[��z�7�	��$2!p�s+�ɔE�Ѭ)�6=�Zg���Ԕ ~���������k)ʭ��T0�e>�ӱ�hJ��[�L�ݒh��h�|I�$¾<�½}����+!d����)��OF�F�{���{8NU-�{e��:V�7Fb�\�IVPa�F��B>�uӣ�`p��Ҕan[�V�HXx8:l��3=RU���M�W'��|�i����U��]�-Xhz׈'��9K���J����
7fO��h���Xڸ���L�AkO�6���v�%o�@LV�#�/���UVzP#�|�.Ys�3A��/�y��T�Mv�Xl��Q�¹���*����2�d���/�heU�Dn��w�<n,���e��f��i�Ǣ�6�@�˺*���
�t%麁=�󂼑�bz��D����mmk[��w�m�ֶ���m�[�����'���ͧ���r���}�a��m}P.�+��P��
4VO�%;��ԗk}�ڱ�U�|P�/����|V�lH�V<x����\�*���1+=-�2���Eo>�^��㴄�粀�h���C�Ev,
 ��逽��ln�aͭc�㳠��R��@�*؀�	��a�c�?,˲j������K������4qہhy�?�v����쁂���F��m��|�]�>�A����9"��0$�/ 2��I����P���*a��D�3��Z}m�V���*q�������m �%�R�����G>�M��Ϣ��a&��-����wm.�%@�����a�=��Qљ |�sh�Y51@���L�q���z��k2���^�N�˖��˦iTEi�GV�sN]����x�0�"� �wH�\��{:��0P6��r�F�e$hA6Q ��))��
����R%�EH�� ~w��,����iˣbޖ��%�|G�܆�3X:#���R�r�z�9���)�W�T]ك*Z�� v
�Q҅a�u�� @b�]+�%���I���e`�L%Ց�1��򩜵���k��KTe�\�?���tQ�q�0{c���2���_|na�uZ�W�Ͳ�!�iv+˓�d, ����A\�%Y�]�M��] UX��!��~�W�:��#��y%�|A��
����H-�}r�Rh��>��yRXg��r,�IɄq}���eM�e���[���硿w���u%Jpv�3kA�n$�:{���-Ŭ�P��¸��Fq�ض��j>q�\� ҭ4�`�c��i��_NʸB^&��D�婟U'��	�d��
܇�I=�}e�<.�]�4-��(��^,L0��Nf&^DZ/b�(�ܪ�'�ɔTo���ʋ�f�&����)#3�Q/��F8��ƁkD�a/;B�D||�V�H�����k#�G�w���/R�Q�������$���o2t�jI��l��nEnȾ��)哩�:��Ƿ�����d���XZ����1Z���)ע��D� ���r��F3Քl�f�a���B��ۄ�օ>��m�����ηHL����z�s���Q!�㴨h��������Ϟi�v�B5���W�".v�BU�>=��F��孥��a)�V�7�F!O"%��1��A�eX���ڵ�dx�'�)��)�Ƌ]���gs\���p=�:M��A�x��)���0�u���w�ǵ���{��eE*J�(�����yS��(�c,���[��{���c���D�^���T��$���=͛�ֶ���}��F�lmk[��־�����������w�a�A}Ry��w�����榯}7wwgUw�d�$Vs����1 �<�艌�� ���8n�j�+��4}Fr'�Ŷ
`X�UT��˅r�ka7$�P x5^g� $�s�{(T_�P܎"�%c��Pb�֦�W���KU2_����yG��0Φ<1�_?��{��a�U�����{Y�(�`��*|P�s���sL� �+v� ��-I2��U��,pr(��O}j��GU>O7+�Y�yȊ��{u~}�a���^�'H��%���!eիY��?����o|�>_��f�HJ� إ�_Z���Rea��ȏ�@/t�W����U��=��l�9��(2l��{��	$�<�� -gR���H�4���"���tx7�z����W�����Y�w�,ňi ����������BH1�c�(���c�d�L��8�����[��U?a�hW�4� �
[�>�TNt16��D�����Y� ��_�7!wu\.�<D��R�y�S��G
,o�rl��Q��e�z,�3R-��o�%��3	8�}�;Η��܇�M f��I�%�r4���U&���,����BU�3+�{Z�a�0�@�%<_ �A�}�e��L{-�W@����}�nؙ7Kg�&-�~<S����A� ������?�7y[��m�aЮ-��U�v����H�9��s@qWz��X��;m��"�sy҂�b$Ivp[��#�2oBz�Ta�T���87�����̟P������m��k_(���� &va磽;7%��:*}F����}Mi�D����ӻ�������B�R�E�(�Y$�!�������U��r��it�$]]͙�[���[�'2Z�����K#7x����دf�9P�u�8�b��kU���^�1?��ZD�15�h��5���>H$A�͒�C��|
϶r�<�+�V�֊�6%�츾����3Ŧ6{L~t����~�W1�KRh�#ef�R�E]s���bq��w�Z	��x/�O�6��ƌDH���b���sG�X�X+�g�9(��`�Y�>�}���}�O�C�}:Q%%;9�<r������/�, 7�g�܇u�2�h)����:k��ĕʀ�BE�rZ_�$R��T�f��d�	�����z�>���8~�߾�0& �a�������������}-���m��x�P�y4���7T��Ee����������# �{#r�SݣA&uVt�m�H��{�p4r2�>AsJ����Tu�dDn{�dd�T�{X��n�}�6��� �%洌��{9.$Re��~@�*(O*v߼fomk[��־[m#@����mmk��K�r������߫�g��˴{8]��(�g
 �Q��I���?-�y  �d�d��FJd�p��ՠ���6X�o���;{�.N�bXT�fŁ�-�A��-�R�2o�m�Z�c���?(��
��W���Y[��jZU���
��w��*'��`Ӊ�A?��T ���������^��z?�Oz>�ĸ���}��΢Pp���yX�9�ڏ���W�+�+�,Y*��@�)Q�Y$Pº�5Hǃ�;n�F��?��$ �Ω�Bp j=K`������T�<�b`^���p(X��R։lG�A\U�FB%�Ȍ,�Y҈jMuܥ��f*l��<0�4o@"  *r�g������+�[�"�t�⤇��^��*+砜�$�I��x��5��FU�yz��3$�9���k C�'�;�H�a��|	�e���@�!��o��y�8���X\�ʥ�IK2�(��%��	T�}�Џ77��$[�H`�2�*h����3�-�o��� V��;[+����F�
@Y2˖��=V��~&���MeT�pߑ� �Y�?3D��H�jwM�{5K5������)߫�2e�^��P��m�bed.��@ Vy<Om�
ƾ?]����^����	6G P�*�U�>K/{ڶMa��o꼹L�Ͷ�e�B�&*��d���urEA���Q���:�˹����K���O��D����E����TS#i�]-Y^��T;
k��u�]E��	�*�{Y���ʔ�eI��p�`�Q~���i�z~�����>�7����]��E-[,F��
�X�F?�3N"� ���3Ua�j��N��l�/T/��B*��[�D[�)[.E�u}r�\Š�+bǳbuV2˦��p�~A;ߝ���1 =� 
kq h|���������kF��
�DS�)_��>��`90$I����3��{S��:R? ��+���碠��x&1��^��~,9P>'�d��!���9#T��r��Vx�*5�^�ȵ���DdeS����	n	蟅}׮�����K�=$ȼ�s��2Cݡu KDZP��l-�݈��i�V����6�wp�_�`�~������@�smd�R�^C[+;���s��M�N'Չ���"���7���R�u�zn��"�(F���2/�g�]���Z�Ih������O�[(c�Z$�+�ҍ���'�����eeɲY����-���j�~^�.p�ߙ�3�Mh�۸���f�����o1�04�D���0����/�0�oF�����R�b�g�&��o7�����ֶ����&�� ��ֶ���}k����������ۛ��e��ק�wn��w��>4�?��+=��J ��^6�a��Tv�m��a�D:h�ϵ�f�`ʨ ��{�('���A5 �k�,Hm�ul.���[Jɚ�Z���@ ������.Z`�uO�����Nk���x��J#�w;�����A�-��3�	U|�Ag �X���F~�8����$6ڛ%#w
a���q\�����׈���]�[�F�E�p8�� ��\��,ӽh�(����D���U�gv��B�Hx�l&�,����y�o��VPS�d�q�ݢ�Ò�MVs����C��s����x{o:�ѳ�B�ڽD�C
P�R{��V��SLk��gQ�[W�%��F#�XU]�0� *a�aPUz��A��0�٪�;� A�d��A�6����tޭ*^>��+l�Ft��q�u!$ʝ;cPt���������!���il�C�1e���:�骎�lZ��������"Z�ǰx؍�<�B�v��|�Tpq&1$��XR:�8�|T�Fٹ�2}6+��t�-I/<R��Dba������J�	�b!�)����#R�fʢ 	� .�T����p�	7�J��C?���[(� 3��Q
��O�*���e=�x$(6�D����(�w6fN��,��b�����I�}��L�,��7q�5���VB2�T��:�6���y.�@Q��$���T$�f�̐,d����K�0'�}�Q'KN:X`ɖi����o̯�Zo펅�6���添�2�bص�`����Z���Pr�F�tSˬ�xn��(Ȫ�e�$"�"��n4��!���/N՟�zWsj�a.����|� kw�{f�
�Zŵ�Vh�{��s��mo�/�iМ��	��Qv���c�����l�a�Z8� &U����FR9��-�ә̮ܲ�؉*#�Z�Q��I<�|��MŴ޷�k"ȮS�X�
kǆ����ޏ�h�\�Έ�����_����B����ID�;�%'X����s��Zȏ`s��t�~�L��=��b����on��ӷ��kS����U�1Q��$��e!J��\J
"�o���|�1�h�i_��T����`u�ڳAV�{�<HU�YJ;��X�Z�>g�����gcD������8�y�B�c������EASoeH�c��q9��,)�*Z�)yob
-����*�Z����� �����#��ɮB.6{�}j�F]�#��>vu+��n�z�Hr��ֶ���}��F�lmk[��־����������߼��O��ɓ��v���~W�����iC�f�EQ�`e��~�L��	�m��-|(bU@���>�C`%)<��Y����q�d{�C��ż�Mj���܆h�K����� F�
��eG�A�L�V��Tg0�o?Ov�j�'� $K�	�ꁤ��A�`����P~��o�S�L3-��,�A��NЏ��V�(#�1
�)�z���U��Y�?���y�+���^)e�hU�&�c�A���HI��h��Y�������*�i��8�reF#?�͈+*;�P1�B�wP*���~G��qh���Bˈ�U*�:��Є/"@ю��<[F	+���ñ���aP�?(��p�����1������������ y��Nf���EK�l��]�Vd8�@�Fil�����/�b�g���������ܡl
���@rr4 �Ｓ9	+5T�w�9�����@��O����Se��U(��6i�@Mg'�����"<�P�%[G �\�A��p��V�f��n^�V���d���-aꟇ�_�	3r0�A6�<v���:!��k�z(%h�%2T (�;����U�H���^����nL��O ׄ��t`_5>�=Ht�:��E����l��uss�OEvm��#����,rx���^��$bH��Dhv��4 ��/�Kp���/Ȃ�J�/�R���}g�Ri9��
氌�W��a�ws��W��1\��>���-�tƋ��݀ԛ[r�à3�@q�������y��;ml�Ǣ�,�=J�;�z��:H��ň�%�A$�Ύ-�o��v�Rx����l��H#��T�{#=�\J�(0�%*�p~s������=;�n}��*��4��c�Q{fa�*�9 K�kt�֍�WS����,}^�f)��4��_�x��`�
tf����u���P�Qp��X�P+Y�E�s�>��Z]�z�!�9D ׋ID��Z�cˋ: ��n�l��>G�S�F��v�-4�/�M�0��-��֙_�&]�_�� ��]\[����5{<��#Ke(�E��R@��'?����}���Ok�����=#k��N6�ID��^�Y��z(�>��=�#��0�񲂀�{!*7�a.�Cr
��G�"��1�`����é�z�r�c�\��e@�O*J����u�����us���G�&vX<G�/YVu�r��JT(\��R;ރ4B���=T�ǰ�]i�$�ml��	�<4�M��S0��j�P��m:���q1�V$��'���1�Z����d�߶'�ŝ!�����v�y�屯�ֶ���m�;�6dk[��ֶ��o��~�c:o���O>�Óq���u�y�wV�� ��P�;�¹>@F��G��P�_�UQ��B���ED���]�%~c�G
nU���<�U$ �������2%S��,����w}`'?ɣ�3�������HFO`v���
��{} <=�yW�!T��<���~ �H�D����.<�Na��� �@}-���a�{��OdE�_�Ozx�nE7'/@(Pz�U��
�D��0� �J%y(����V=+�Y	�*����ύTB�?|��p��R�� r��C�.��Y����DѪ��MG��Cȋzb����-���>�*�d}`$��k|���!8Oz� &fA����������бk���b	��A��.L�0��+IcTvȬ�JYBdW��֟ �4/T��
P���eDf�$�(aw�`o�=�6��x���.����r�<ZEm�J`��F��j����s���T�e!��<v�0ؙ��Y%Y�j�gV�L���$yp2P�hMU��z"a��k ���DH!�z�+���WU�F)?����N�1�ٵ|���X��V�M@�Z�V*���Hs%�`_�c���0�$!fbW��� ���ב �awS��K(����P�^IeQ���ڃ�	�aM\�����9қW�Ū����&��f��?��{�H����3�3�� ��/�B`�u���~���;Y��_�3����>Ηa{���weI�;�y�O�]a0�a�����mTo���*��6�ǎ��~�7�*���P��Birp�7e�Y_�����y~:��>}�G�~2�;� nJd���!4��'��	&g�oYT�X_y�_0�f�صҭ�J�MŷTK�a�Q���� �r4k2'=\�3��l�H�����އ	&(*�ǃ�JR��T�o��b^EY!˽`>��$����|'"1/]��t wf��]���{r�emm�Y��'�pwB�<�&�a
UU�'<滻�p��XuO�Tc�=f����8`=�&������\�yZK�=�ddIR#�}M�;�F�[~�>S�+�^�u\u:ڨ9I�_A�/e��=���k��d�?�G��}][���2��"�꿡���j0^�l�F��m��Fl�8���!�HP�Ҫ���e���wr��w'��*P#1�F^��.v�F���;��h��~,�=�޺��L)T�9���R�����5�k���4O�F�&9�]�ű�_�]7З ��	Qr�9��/� ���8�5��"��@z�6Aʺ�L���=$T�1�w������\s;X�������CGU��UԵ���k�Nn�Uk=�ˠ} $:o�����Bk*��(!�j ������Af�Y��Y{�˺d#Y�AQ���\T8M�K88)�}�C%K|S��Y}�g��^�yl�ޭmmk[��w�m�ֶ���m�[�~��������[HY}�>E}tss������Ws_�Do��Y����5��l^�M/cZ���AVVê:���JW<<��YmYp�_�h�L�[՗���={>��G̡����:��T��;?{F���T,��=�f~�.�B1g��+k��@ U�9/�On����Ջ-i�1:��*m<�T-kU86�e܂ai����z�.����T��r��J�*r�m5zAY}\��$o���슥�U���eY��Yv�f��|<'B(��]ꓩ�h�"c�� &-���Q��)�FB�57;�h�9Kn�S�D��}�R�MTG�[*�L �3˕��|� �'\��'��u-̢Z����]�,��",�� ��C	�}<���ch}���~/ri�c� � %�O�v7�~�+^-� ����t��3�e��G��pK%Ι$+��ԇ)-YBP�a~��-��t�!�4���>>��_���bVr�sqK-��_*�CrAB�fI$"Ê�����Y�p��ݛ;9����Ñm��+�%Y�y食Aba�Z0Kv>�dF�Փ�:O#�m�����m����O�e��9����SM�l�q�8�,��M�S�8���hk!�,}���A`\ϣ��MyA�`���Sz<f��>��� ��۹072�r9��^K�_�H*�g�܁��VD��,�vig`6��s�ȱ< *({a>ϼn�98��p�9>���cՉ�\��^c���\�� ��| 0"k�Q�����GO�㉦���ǋSi����Ŕ�Z��W6h$��$F�`��!,�~�4U���s���-�����w��ҫ9�L�\�y��$�F�G�į�z(
Rs#���� ��
���s�7b߮�~�묡B�wм�^��*�`��J-�*5����秸
��>�'�:q�>��y��D���o��siV�~\N�x��D�&��+|��>��߇�{���M�Sx���Z&���n�"��,�Z2�H44[I/�7�����iպ�@%�T�����`�iK��9��Ů��H��l�6�V�2���A�𦈴�3;���6�)��)�OZ��^�(~���ʤ���O�\Sf����}���t�>�������-�k�>��6��?�<eAba'y.Ѧ�EV�Q�{[�M��Jf���7�i&��� ��@��m�0쇇��wu�����������=����O����mmk߹� [��ֶ��߈�O�ɿ��������4�/���8�S}H�񺿜��Xy^�������@E�'��H��r 5��� <�Xzd�����(�A́�B���j�r�x�:�&̯y�.VE�]EǪ�2�fMP� ˷��j8$"�I���ru{�IY���P������e�N�"��70r&@�l'Q��UW	G ��_o*
<�G�+S�ܔ%TϠU �z�-V���^:ޥob��������Zx9ǘ6d��Q�v�g�3
-&� �Ja�沀A���£�Q����
�vT�ч��f���t�C����V������0O͟ǖ.�0��DVuhg�I�C�A�Y���0TJ��-����	�`�m�ڰ��5���x�t����p�ڔ��"����B'@9�V��LK%{7�?��1� ���L2U�l�T�m��;^*"��K;/��ur�Z��#�8/$��3mD�X!�eT.���լ,��(�ֱO�k�3=L����r\�fF\���Kv+�*fY�n�B e�5�#	MT�f�D$ܯ��R�,(^U�q�[`-�v�M��� Z�-q���gT���kT�nmM�������}��[g*W��q�:"�=fP���
�mT�6,˸�=���h�R��p�_�D�����54v�݁�}̖7��\#"�"��tsr`0I�:����Δ2;�+�=���6���i"cF��~��:>�pP��K���y����.]������o��b�eM��Ս@ց}��@��,�5->�� ��f��l/����@�p[Y�Qu`�`���q�yn�l�:�"�eH�����h��"��o�������Jm�{��G�A���#Ŏ�Nn���q�gp����Nxb�h/����;��Z��e��.�Ś�]��R�I3Y��IK��qL>V�n�w��rkȴX�²g��J��;漼�nek)���b��$��ɺo�y%"mG�j�T��c0���;�ٙa����Ί��h���|j���������x���U�Y]]��%#!k�Zym$-M�S���-;�����Ǹ<:�i��G���͒�hR+���
N�<�l��x�q��t�֛���⚶��ڐ�c�O�ϫ������[Q��ԲtH\Ң*-�[�ݣ�ϔd9���l�ߢEcb>˘r[�RIrj.���ݰ����ċ����������:n/��>�����'����ֶ���m�;�6dk[��ֶ�ӆ�{����>L>���SL>y�Ρ�O�傪ZU�(�|	����jj��4"���\A�����H�ax�[�AK�n�+H�kZF,�6S�=Ǟv;٪�G#��"eJY��l�p���(f�T���0@�UԽ�]��U�pT�1����ar0'.��u�@X���W}V�4J�� ��"o�;|��X�ࡵ�I�	`�s}���5���%�ì"����ԎOc\�� ���<+���  3 &Lztyҗ�'���~�%-a����`t���𼑾��5Nd�Pv�i�\�A�,�p�<���+&< vn��j�$��%��4��L��'yg`��L���$��Eǥ���'����_�8P������}���x�S�`�6j�ZrՁ�-��G ,[t�Z��d'r>_�~��ӂ���q�����扔G^��W �}X�U$�	�Nf����d��?��`��L`2A��|�8e�:�d�d���[�~��B?��J<�a�/�ץr�)7)ez���)��,�B���;oOn�4+3ꠉ ��4b�=��,sb�g`�?/zen�`�����s��V_�}#�- ^�3��@�qݫ���sn�M%���jsM��b�Cګq]�W�[s�D���Y� ����S�L��Q�2F ���]J��		3S�PIbǱ�H
�x���p�vP�ISW;�{��RfHlsm�׀zY����/��W�v��=޻K������L�1B�;���E���	� zX��vm���-ZH��^:>'~m}����8���Ot]�<�1:	�d׬���Z���+S6"�<��w�)۴v;)R�%��d9ج����
Dc��G�s�|�=*h�Ҹ��x�}������xϐ�>�p{�$��
η����v��%���J\��y�LAd�l�N�xs��y�83�C��T1�[���M)�r�D�"���,�@����?ΰУ�&�����mhX�^t�_�*��I�`��-�,*�js�i�"A�*;���c\):�]������b�D�D�%��������2LEQl?'���Hi�����o+�Y�+����_ʫ��E%6�b�d��؀$���,��6�x��+��G�,�'�Jɡ�E>�i�a���t���t��~e$	o��`tY��ܤ:������r�0uXh�K�X�����W�~Y��u}�/���}����mmk�ɶ [��ֶ��ߘ6u����y��/�ʗ����P���}r(���#������C�f�B��~U
�v�R�;X�@ʞ �=HfU<����T����ڦ�+��H�N�3:ѣ�v �H��h �������uY�WQ�C43J܃�ѱ�V���d�Nl�@�v^�DX����'��y.���O?g�PR�Y��N� �J�ØM�0��I��*��|�~��R���<~0��Z��
�� ��J:	�ͪ�N�B�����Ǹ� 栒�0��,�B� �
�sa����^��r^L�#"j!;VE���VI�n7XJ$']�rC:Y�hx�
��ȵ�L�)7�T���DPg�7 ,DT�lv� 0�[0	:
xKVQ�s�@��d�\���0u�
M��p�dV �{P6� Bǳ"�5+BvE��/ngB`)+��Ċ�O�*?]y d)1C�J!BY`�����^
�h��[�@zw]S����u#�>
��;����Q^۞5�������5��Tt�f�m��b}`I�<���� �����2M���)x���V������*�;�9�/\G���*�b�h�Wvn+��9�.LVY��������7����1��p{)9Թb.6rJ�����*�-�D�*� ����ͮ����elI$Wx X=��pY�l���H�`c�do`��-?_���e����}��$ ����R~5���>��Y*�M)�U>׉!�%�C�"�� t�#�'�n��jnY�=�`���^>�͢�v�Ȑ�^�����%;�hd��~��SZ�G�� %Glk��Wx�7?
ޞ��/fK��P�2�i;�,�$���m} ��˼�ؼ����~ZYԩN��yh�ؿ�,��ʮ�Ӹ0�g.�֕�����'�r/��]΋��䧝�A�aꢖedk�?�[*Q5�m�o]�dc��Nt�\#�p�<^ܿ���|"�������d�r�\9�p�����:?e�# ��e�%'h�@{�>��U�Øf���<��U*��J�f�Ӡ���;�buQ+3Yݣ�d��-
JJ� E���n6u��	�7H����v���Ȓ6�r2���]�$�Ď�[�̳9�e,`���i ��>|��3_
��r&��k>����2�e}힡��]�{�Y̻v~�:�ɝ�HQ��;�����o󱀸��j�~/�`��H������>�/��.�_t1~Zo	^��mmk[��w�m�ֶ���m�7�������~���>�Շ��a)�6���E ���@��T �R_$�,�
ִ�ߨ�[�z��?��PuÚ�2�޾e%�������
�h�Yx?���6MP�|
��l>ǐ�CQ��{�t� �� @3(Lq�sZ�$�NQ�-�ŝ\�ԩZ�o�<TU�}�t��pk����Q1v���Ӓ�`&������$���$�M7+�;
 .��HWZ�����z�������zf '�ᕿ6�/���~OH�	0knd��ۭajK�.��w���y�,�t�-O�g(������X�\�*Z���+iW�1���`��:G/�s�8~A�A���.r1��`��U�ӂ�,��~�oIV�c�
���ʫo~�k+#���� �F�'��NT1x�Ș��.��J��j�.)Uh��(�����c�+4���kkӃ�]Es=_-Wd0�{�TT��G���B�;�RNx�Eh�G�ǜ�z Ϣ�X�M"@�*|�� ��IQӵ<�Y�hJ�1){�>v�\���jl($dg6r����ϕ����!#�{	�{�}Pk�\p������_siʟ�e�gw��O�|o,�?)�� ~X M��TW��Q��d9F'�x�ih�ܱu��^�"1��z�G��u�ú�/"���Ւ�� O�i�+���ה)�kC�K�-�y7�x�w�+�@�b��5i}��m��fQZ�q�M��G��o�x��2��!�ԔU��W&�|�>N�"o�V�#R�rFu Y�lCyZ�'�|?[�*K������{�
�=��ɦH�f�w�87��Y�q��å"���k}�|�v2t�:Yr?�����oS�������^���SZ�k��o�|q�v�u/hZ�9�vo47����U�ַ|�����g8a�X0��9�<�vM����SR���5�H�)&�A�K��"YYZP�����Uq��dEтץ�$�������g�XB�ԒÑ�;%���m��q�=)�oE�g��,�9D�H��R��w�F���x_�w�<�h�N�)���2��T�E�$GY���q�,��d
\K'���SO�n���P�䊣�Vq���m\��Cq�&)1>y�l?Siex������ ʸ~~�(y��b�h�����4�wdIK/�@ `���ñ�c~8�N77O�ח����s��n�_�����>	[��ֶ���l���mmk[��oT��_��|\�r��Cb9,������ׅ4z����T��S��^��]�R��ɺ��H~p0�_�f���A�am�#�7)��DA��tۧ��}7���EP:/vG�p"0b��EgU�h�����YUp��{����i�e�ӳ�a׫��٫3C��*eeAI��r�cP5T� .b�
�N����P�w�.Oʑ��^�t~�~�eU�M�|��Vj�"YP�,�c����	rC���T	)�G�$ȣ�E%yN��G�����s��x����3���y�Á�K_~�{.q�ބѼ����|�Ki`��Z����5 L�8�ffxH�Q�B���2��T�N�x��JfQ�/���	ڍ�Y~�J��Z��Q��d�|�۲�|�}�4q�XU�A
�q��^#R̰׺'吼u���V>n�6/U�J���j�
��WK����FDh��V��P��_Z�����H���b��-�G��q�&=߃F��*��U(rSY췜$a~��^K����
�q\���\#�� 1Ǿo`*�t���D\I�̑i&�ԈY#�0^ �������͊l���z)�+=���uG2+�؈,������m�����1O_�q1g)�T���r�Ir��Z��vKT����/���a���;���f��rk�̾��^�`���Zy��~S&P�F�M{	�k��o���Hc�Y��{�n��k�4�ү���,�D���b*/U���v�hc�,��is�-��B��:lvZY}���S{���C#?\���t;N��H�ވ<[܋��QY��,�a\悓�Ӵ�a�sX��h�mO�L.*<W�$g�����}8ɸ�����zb�ܦ��5-�ao�Y��V���.(�I}A[N溄HN��m�C�a��5ǃeH-�X`��Ո���cN�������i���R�Φ�,E�����`R����X�~qЄ��[`l؇�2�=�䠽O�g𼺅������N��U��YV��iQƇ�1{S�q?�y����2T��f�J��5#����D��R�:TV�=s>J�R�Zئޔ*�p�Y��d��
2���6����Ԙ�h�s+e��j3�]����RP]�"�m�B����
�nj�ڔu�$칸��>4aN�z_�5���x|v�������O�g����?���㰵�mmk[�N�� ��ֶ����F�����_�ÿ�����>�����/�����������^=�2%zEhZ4�W����_��P�����C�!�K��� '9t4�zX$l�B"<� ����=`�C��������=��U�z��T)���(j�YE{�����V���4X��-y���;�nX��D����y���)���p>Ng>��>�ȁQYmG%�����K��ڣs5Ȥ��X~�?i� ���YrV�+��>��*�1�a�PQ��٫O�"����1�)(:*CX��*XZ�'�_�壀lY[�ՇUņ�c\�'PK�&z���f�մ�nnZ�x��~��z��l�{�@�*
#��@��U%��G��CbÂ�a�v--��缇��� P�8�����n�3;:�9��h���Lz�ge-��*D��V������ίx4�hY%/Y chใ��&��=�g���l�ݡ�3@B6�Bsy2��C�@y?�5!1��Q�,�к��4r&�p�W(9���k';��}��^��A��βj�4q[�`�GOvSM��D�5�Q���ue6��1H%#rc���cCb̈/>�2X1l}0�{��4��� ���I6Z�� ���m��u�
�wb$r�� r�2P\Q��˖p"�̊s[�
ZD�$�/�>ֳM!υ��p.�s���;�Sp[/X��O�+�s��+$:�П�p2ܛ����}l�a����\��� 4✜�X�CX)d|!6�h`NDY։�����\�?��Џ������r�0�3n�v
vm|��m���wuVI�}��'/y'�rI���4��W�KF���L��vFn�������r|�����L�B"�ڮw���*;������t�)�D�e��Lb��Yb����2WJ����gm	��]��y��h��%u�B�=�Λ�ǔ\���Wv?��
;le��g+�2��Fx���h=�W�f�8��{w1e	��}��P��@||Ea-�Ү�7��"�`#��{+yx8�x�rm ��A�";|�-֖�ȗ!-��F}�E9�ކ���$ʥ>D�G���u%��N�72�m$�+�<�]�dY��Y���Oʲ��
��h�(^��u�ۯ��4 6v�e{���b�������<*XU�Ղ�cw�5�?N��w�n���w���Qa|@�� �ф�?�v$?�4?;�ο�/�����xz���z�_��mmk[��w�m�ֶ���m�7��/��/~����F�4�>Ч�~�������N��� 6�!9��<�<�����%�:��*�ak�a�-�4�fE?���c��� x�4�Y�R_�r\��	�*���<ã�^��R�m��]g�3����D���0�)ܫ=e���]PX�(��>���:X-�|^�\*q A"��L ,`��Ǫ�d���@`���"ߪ�'U'��b2��je˰�ر�O vY�]��;�5i�Q���s��{�ϴ���e�g���g"x"���:���E� �t���藪����d��D�!�H�ý�)H����-�+w��ʽ�Y�n�?��6���U�tk���Q13�{֞�X�MFF�J�k�y� ��2�P5J�D���7��`y�͝<� ��1�P��U����9.��|�e�2 z���jx��������G9�=Ȟ�WI�l�df=�N��}b�F�9������"`s4�fY�.>�U�s��?�n�Z*�.�;ڡ��eXT

ow�4|UG'%�����Z;�y�φ�X�l�s�%���֩X+ړ��y<+��$��nPX��e�����8�����X	�����~�����.R 7Re���%]�s\�Σ���}?��t�р.�p��Y&�{ Y@ �/1'�����#s8ƹ��a77"ƺ���4���CwuoEF�<{�Ȭp�}Or���Eʽ~!}�9�k�
���:�[UΘ�9�O��wf75�77m�2��{�+���R�}�J�p��R6��:�x1k_ѹ�F,{����Q�-�'�+��UaS�1��f�J�D�2j&SR�O76�g�<�ɥ=@�5U2��~6����ײ��2���j�at������"ns#�a�z߾�B1���x��J�^�'�w��V���X��������)\�����#��2�Aܓ�t8A�y�� �]'��[�I�	���~F������R��M��wye����y���\LI��pu�.
]o��]M� �M.��Éw|	zm�]w5��C���T2n��~��-�L[7*���9Q�7�8�Ɩ"�4dc`oD�N1;(Y~E�$G��½�w�yc7�}��a����y���nzֵ�WbC�U)��hy-f�	Ґ��k���>��ܗ�w^���b3�����$���$�|��k�'���Cf}	r�J�4i?���.�,+�9!��o�^]/x-����d~�z�y/��~�\y��uD�p}+��|�mW�嬽l�H8��ә��=����=	"�%܏^.T~�^�5ὧ�D��y������b<�b*�?��Gu?�����'����O?[��ֶ���|���mmk[��od	���ߊ1˔�>G��������k`�Hx8���6� ��bY K	�:ȕx�<�_?��o���֤�� ���W"v��P���5��X��<�B�)�EϢ���1m��jǗ-ܬ�:#�\d)���s�~lUË-B�w�a�����]U��f1ra%�D b�Ǧ"0�L�[	C}�/���m =5%�Y/�����ls���:���pо�1�f�Г�	�^��1���,�eG����K�7o��@� �H�Y {�qw2*���sH��g9�*��Wg>�!Y.��*l'���T�ؾϹ2�B[`��fe�X���l�a���p�d�Rm��b!�*�b�&�������aV��4��K0q6B%S�Jl�;�n̉�P��n��J�^ʦ�X��{3 ؐ`��{�^[��Jh�_{�s�͛Y��Ue@�n�'?�Z ���,��C7�����D�74O��-A,uK�M[��i��ˮ�nWeUe}d��{�9g��X�5Ɯ3"�ɴ�`!|r�Rֽ����bŊ�1�Ƿ�W{�����C��Πb�d�lU\#b��$����Alܬ�IfyàgU�@��6NzX%�ٙPP� y���ᱳ������^G*�e-��Ǥ�x�6[��^�g���g�d�d�s�|�9v�J�f���^H���`�@#Au�V������D6�u!q�
@��F��q.m<J	�s�󰳮��"�jB2�\���.'fٜ�H[5��>��+[2 �+�:�ɖ����ZJ�$t|�.�������k�	gX�n���j�е7���jw�Nq#���f/0eV!Z�PE�vn��	� ��&�ټ�N
�?�8���YE�O6����W��ΰ�϶6&eWc�M�������Έ�J�G�;"٫׾͊��:����Gy��ҵ`9������b�F��(��`P��r��n�*.��V1e����pYv9��v��x�N�U%v�E���ݖ5M�7V��s}l�f��uKLԌ�����c���l�a�[h����$k7?&�վJ�O�u��Y����E�;H���⽐n���mk,ֽ.��:-��\�����*"�\������Ca��l=6:>��s�����6�W㌥6�p5��~5�E]��&��Q��	[W�M��� ���0<�v�>�]�W$�dYi�e�:=��v�I���ҽ�.U���vtH��R��i���/9z��b�,�D@[4���D��.t'o�8ݰ�١K�KJS?�S��w���߼��n�?�����r��������������B����p���/��o|����e�x��^����2^n���OD�R�Nmno:
 ��1�/�p������'H���3,՘�9a�� d���Z�����7���!U�Ө����}�G�':<��Z��_�~ϼl����,���̼��?g�Jo.{7��S�o<��2�p��\��aY�j�e�R�9j2���؆�IHL��j-/�^��nI\X౼K���9�m��Z��Q�1�f(W@t��1r˄���Z1m�����&��#�!}/Y�EA��e1,��\ �����0}
��||��Эd-���<�a�M��s@v�F*��R|ݭ�҈���~���F6�*�"��|�ك	i��ެs$��4xT�Z#e�47k6�#Yɢܬ��~���L�J��o'����	��<)q,�㛭H�ɶM��*k��	x=�HQM�Z�:n(�*!�=���M�ْ� �����ܜv��V}�U��m��i�!d2�Æ�ɴ�I�y��\�W�2LT�`sg�r|�5�.d�7�,�rXr�����I�If��pAt}3�$i���˺�&���V�����8gJY��&$�L3�ւ�s�,�,���ƬH��+�^9���8Al�>цI��5$�'VK�y�V�KދX�`�l�,`]��o`瓅��B�N�4|X�<A|��{)��#�SO}�t[H$r�7J���?�t��*�Q-��uv�� +H�qƝ��<=��<��	�{=��ˤ�?��l��ż��O�;�.�mn�t% o���o7;?;8Zh�p��K���'jiH>v�<���A�uAg�d�l��b�ZJ
��D+�)�2[�[B�q����{;�Ӣ�]Z�=֭�%�/"4��M��Z�q�c��k�ߛV�X�U]�ǝ͖��|M���<N����B����v�/v��ZK��E�\�/͊�s�㠷k&Y2]�y�\_1?ʬ��[c�H�B�<�h�U���-�d����NO�)h�����Wqg<�������H�CRK1�`���֩"����P,�h��w<,�Ôg]3,�n�:��Y�6�Wy=��m��{Y5�oBvFn֢v�<ɴ���RG�,��yۣ3%���l�u=�(�Ij�W��onE���s�ēb��N�<I�����4m
 ����t�d�4E�EP�2=�������oo�n>>�'����?���K~t���p8�`p��p8����������o�e�;�//�e����aF-�i��8�s}`۪�,��?�/䍼4Rr����C~�5L���ݪ%�"~�iL��juv��>Ӣ����Q��D��Y��>�|J��Js�F��g��_!.�Uv�]�Ӊv0 c޾} �g�� J@�IFC�(��)� �yA�
��:���FXc�m�����dȫ-UPk�R�CA�8��:K��x��Z;A�>�7W�	��U�Ġl��[��9�e�
���&m��EZA��}�$�Dz��E%�56]��&�[,����k=�pl��E�e������� ������c�*v���ׄǄ��mB
"A�0a#�A>ۼK�O�f"�%��&"X�G��#n��rfxt�
�$�װ�Z��F�1�|�Y�_��=�K0����h��6��#��34����9�;NܶV:(H��f�����B���L��h=q=d
�&*Hn@�5,��|�>O�f� ��o#5���xkP������y�L1�c4�| ��.�E۶]����� � �M�}]sdl�R=�Ć0�(���x�r�f�<��f��^�
$)��bH��
����E�j���Ϗ�me�c׮�W���&L��u�����X3LX�<�����Q��w�$�]��5L"vL�t��a6m�v��]0Ae�2cyF�:��Fv�l���7��_3�9ylf�\�+�*!vo�K���y��4#�昭[kgV��3K1�6���N1����� t�9d��j��
&Iĥ�NJ���P\ױb�VI��].vlE�+j�T�uyY��]2]�	?�?V!,��CX�!��jkרP��͚�ϖ�b���o��f�P�x=Y/S܎�:'�%�b���G���PA�>��oVv"F\���0�?0t:N�,���u��}��lVo�W\[ F�����`ݬؙN��8�5�HkYEظ$Y"e�X���c(o�+�}b��Uד���m�Oe�8���E�)�l&��s;H���k��u�fJl/��N�:VA'ٿ��t_5I�`�b��(�_������W���=�X�2SH�s]Wh}�u��[]����.�a���_?�2]8.��Կ��~�Jzu�;��r��Wٿ�����q������?������� ����K�_�G��{?�s�>��և�S}���iD��}	�֬��H�JŲLv�wV7�<Nk�_H�Vγ�8�x�`��`���E����b&��o9��!�*hH�e�pּhBk��t�� ��<\�'�7�(*)*Ĳ��c_�M�U��d����w�o�{�j'&!=��է���з�_��t1k<CBI8JG�|n���U��OK��_�1�J�2�~�ǢoIeV�R�֪�}>�ˎ�1E�exI��c��u�$tU*������t�6�P�}�s�r�^��T����Aw$�j��V�O���Y�MXC�j״y��y'��Z�İ�[���[g �5Ӻ)f��ջ*A��<6�[����[�r��k�6�P&���c8>B0n�a%-���"�&�6����u<�Z��D�Œ��f[C_�hU��ꜘ��X�$#uv:�}�E4��z�Ӏ��0�� Μ�e�Έi�Y���9�j.��~�,�f���	JFn�1�XP�d,P�[	��U{�:3���e绊/\O�Y��y���@_TwZɼY�ɜh�6g��k�^�t�a=�pk�C(q#�Sr��|����fe�N�Ns.�\+k��S�r#��<��XF֛%s% �q=/j7�׵��O�{e�Yj�t�i����
�=�-6rf�ٟm��E�U�Z0�B��Q3:�w���z�����QJ�v���m���M�D��5�Ê�R���#W��^,�&hh�6F�/_�٨��r��y�	I�ϫ���H�q����P�`�R�ޓX��u��>gflm�3�,j�Ȏ��Z�؇�[��Y��J�����������͵�͝`v^�}~7���f�::������:�%Jgm����j$ܞ�L*��a���Y�]�*h��u�3"���E�8�m�l��ɫ�U�&�V,�\�[�t<�i�I���$/�z�c��O(�.���vY�T�S��ށ]zōV��Z����ǭ�ʊ����}VʛU���̵�?��qv�\߮�Ed���|���Q��6�(��s`H��[I��V�Q�t�Zh�h�X��*��@Q����v�e$�,��lKc8�݁�{6���߰~:��z��������X�w�}'��:�~����p8_H� �p8�g�y���mC۶�0�R�ћ�����CW�P���t>��lQ��J��ҥ�Jy@'�0�����׃T���)ˉ�����E��(>��
;�w�0��f�$�*����S����h>������+�8�A�}W����*F�0�n+��ş�pY%`a��%4�wRa\敩R������U"�򚛲��[:���!գF|Ʀ!�" �-�������	�~ֶO���BH�f��B�%����� V���ħ��ݢ 1��3$F��>�*0���A�V~e{T$��A�e���K�k��U7[e���Y��%Al&AE���^�r#��]S��������V\ǵ+F�UԢ����Sj�vd�f5���8�"ܞ����.�s�N��~>���$=�?�P_TF*6�-%s����い!�][t�D������(6R[Xxa��Y�9:#򖼉%]�֌�l�Q��gf���	fL	���[�e�����g�m�k,�ª�"�t,��g�R���У��mnX�P�1�0gTBT��$!� �l�f`mon5$:����:G:�m6F�._�#<�!nIf�&���e�uF�YYř�ݺ(H>òL��Y�q��X�Y'�	�E+�)��d�_ٲ��b����/�����G'p�ouΰۣ���x��8�"���*�S	�r��D�@��=c犉6˲u`��Hq�%����U����-W� ��D�M C�A=�㲮���$Q�N�`S��j��e�4�����*��Z�=�Xd���&~�8p���aU�>���l��]8>������1������	̵�I*&�+���)��zN��n�Q���^B�m}�f_,[�,�x���2y��\7�&��n�-�D>;��d��\�S����F��h��<�;�Dv�Ņ�"����E�	�l�l�]���&7�pnb�[�	a��>��P�Q���Q;4���U�/��[���zL��sXN�u�Ц�ZjYq�#� R�W��I���b]+ws��^`y��a����,D�m1����m���X��$�n�E3N����^C�97��L�`c�U�:ͩQk��a�5�{d�v?2�x���)vσB�yHp��������t<q�G�-%'��'����o�|��O���������Y��J\~��������p8_X� �p8�g����O~����f���t�x�F��C'�_�������i�.��𬞮�<�Q�
�>��.J��v�О oU�x �&�6'y{m/����֜>��c��~!�В�lH�N�Z*�B,�� S��Y�:��IA��)Q�F��
y��ͭ��裿t��b�RQT��Rɿ|R�l�)�e�)�ԦG���/!�q% �*XD�v��tX+iQ!~(��]8�	�$ct☇ɠ�tܢ����OY�ֳPs��VN&~� �#&�s��y�B��k���&n4;K�Q,1�?���z�EA�&%i�T�X��K��smu|��H�9Hq"��j��qe�v�� c���"U�Q�`aM,�TJ���bD���&Fn�`��3}�-�~�����=AH+�'vo&���c7�Z�gv1蘘6�l��ֹ k怠G"I56�ԗ\�r��e8mT���Uf�H�UG�xx�(A P��}U�e5��㱨�!�TP1,��5�d�표����e�XӜ�Y+�Œ%�X���<�U��xK��&H�;��]�fH�Ze+E.�Z����Td͋X�s�$��3���&"@�F�Ǎ��p�鶨8�
��-�=����sm�,����#ѷ��B׌�c�!ް[�Sѳ΁m�>+ފ&#��Y͘�,�3�JA���UJ_��B53JY���^�����|�q����u.(a����c�v�u�I���Fs��ڲ�Ĝ�v�m�z&�Z�q�p=vl�^.&f
�k�^+��2�Ղ��]��s���J-���`��SQ��5D:��:��EkǏv$�\�*��D��&0a	a��
��sbL�4����i����m�v��ca�hۨX�=�Od�C������]w��{��Ѭ&�n5���nRA"i�} Y>���LۣC�Y��ۇ��R>_\���u�����-�#���^��`�T����+e�2��m�`üv���O��ZmmeRq����k��)��y]�v�����l7-��E
WBXo�p���z�l���gq����m��MN?QI�<7�<n�բ�'�kU\]׃��O��~w�)&S�[ ֠�s^�v}0c	b�n+�_á�^˹�������c�o.�R����}t:�������������}�7�V~�n���������p8��p��p8�_�G���������04FT٢Z83�����<���9�Ť�U*U��Ɋ+� K�z墙Y�F>�k�!��v���p��|0 ��!!C�U,}�������Qڔ�oyѰ��h] gVT6�LM�!��BT��$5�|>D�|�	�6����/(�Z�K�?/:m��;+�<)6�B�t�~6	*ge��#B�ki0R-��Bb��U8iL2�՚�$	���261r} �ص�'֕H�x0�cV?��5B>��k��Hb�@,�=8�S�f�l�"��Hl��Hs�G!܌�/J��Qԗ\��1V�m�)Q���~hwi��%N<�Y=�YgZ����P��i��?E`#rqR�L�4���������j�7�^̒���]�7�=�j�AҢM$�fJ�h8�F0g�~h��T?W�f�`~�OC��p���4�`#���vq?4��H�|�>*�
V��s:�m훘Y�S�S1�D�H�Ps�ԑ�ǰ�gC{�ҡ"ǁ�!쐂�����F����Xv��b�4Q�>�c4k%paG�a�i��Jh���m�JZ
�(��UQY�T#,��Z���Ë])�F�Y��0[ 3:�
���fdd�N��2EƦ݉�Q!4��xBx��[����
oK�Z���H�&�YǓ��V�z�o�'6�B��&b�X��
VU��r��䅈�٬D�`%V�Ϙ��OG+�f��2��:?'���C��~�i̓�|�����?�O��}#��y/�@��ф�:���5+!��3�a�N��Qٺ����V��uZ�x@���]����RJ��w������]�`�	�O�wj&�e��[�c����;qUD��^˓�d
+y[$E��e ��𸭻. ������t�ZV�S�Ӝ�E-!����w�Z9���ra�j��"�������l����	"��u�������&]��&e��)p�.#�g4A�\�}Z"=(َ|��K�v?�蟗�s��=�u����ق�Fp�K{!�Iwg=�c#YD����~n�*�(bn��6b?g}Y�6lGJa-6�.���8vr|��k�#	#U�k+ƨ�wE�sТMOV{�:��B��y������aî�E�;�<�]Ϥ݂�覀���9$��iA�<���x��aIm��W�]ˤ����m��5l�"�@E�%hAf߄�_m��~��V�I��>����k�~�Pω"{]l����h?��'?���/��n��o�������o������������p8� ���xf�ů�AZ2Ѵ4@5?��61�e�jb�7%\���Ɉ\.c���	���I��e�j`�Ɛ��\߻Y�`�)��U���}|;
~Q�	�"�հa�h���i	�渑�Y|�a/r����� Hb��c3���4��"��<��x_�gz`� o;������o�� ���A�.��`�=�#�&�Z�Y�!"�(R�:��iHK�v��S�ꘟ��/L�f�㰄e���D�<H�m��M�01���{I�B�.�8�t�C�� T
A4������)Jj's<���N�@B��3o��%���P�El���Bd�d
I=�sYY�D�i#��傱{$p��*��4/Z� ةHf-|�B��q�<9r��qῑ��yޣ���aW�*� ���|RH���6�3Z`�3���3���h����,t`,j�U�����������n��R�� U�Q�J�;˅�X"Uɑ�ݶR��W<l��{�E����J=V�3�ɢ�4�yX��s@���f���8/�j��wv!-B����$��v��U�6�c�ʃk�B��>�ڵ�kEOR��� {��n�($�,|��%+IA�6S�p�DƩC
ºA��gYgpVv �n�ŷ��Q���7��mSkJ��|³��z���q�P`���/C='a�&�S^v��$�x��VeG�DM=?�1����̐g�Ǡ]Z%�D,��q�GѮ�CO!��
�F
l\:
ّ�W>�{]�&�lՂ��>�Q���Yc��5SK�ӌ�g#o���)�q�wC���E7ҢN�X��g~X]�&R�5< |�x�XP?�;?�Q��䧆De_�{�c�n�""�\ZX5����EK��$8sވ_�3H�-�����EY[��vf;�[*�EPʚE��U�5��"d��^�z��pG�M�,%\� ��>a-̹	�vЈ;�t�цjY�m7�t*�cn��n"ȵ�G +%�j��rP��6= �	r^4� H��fم�a<��3+�3;фp����M]�&��e�V1
c���џ�X�����שM'�w�K��D l3�/��M+k4րN��1O r`࿥��sݾK>3+�I���V�T��U��8OiNO�����3��"�W*�`,;�ԿC �.���X���9�56�x9iP{J��e6H�͂�y)�L���kQ;,�I�I�Ϣ\ƥ� �c��	`݆��Yֳ��b��B �_���f!?�c��tH���yT׆D6St���t�����S��u\��I�E�w�%�E��X�3�nRmC�օ����3�o�0����{�:
K�opo�&&���Œ��J��حܴ�)$��"#00ċtt� �4E�D�l?b�s�?�=���=�xt,���[ʽl�������AƖ�XA��f�P��om]�Ѕ��ԗ����ї���������X����w��/�ڷ���p8
@����A�AA�X������K8L��X"�4%�)��ӀB�-dDF�
7�9���j��V��A2�~�l�
��ag��u@H��?�p��q�<���#�9��M���H�(H�;,�R�U��R�y#�A��I
�rhWk��x���m���JB�Z�j%4i@`��X1IU��E:Oֲ�,�:jS!�%�MM�"6V.z�U��0 U�QؕA2|��`6i!y�ύ3Bg�G�i������c�����;�X�Ġ�G�$;f
�b��nv(y#�*���@��Z�Y�(hZ͉1� (.ϗ����q�~Pb�M��rrl�s�̏\Kw�����i��άB������4Es�t=��Z�A	��Ю6a��6j���9/��
%BMӅ��A=ēf�^�:@�J�
��[�F �%��|�>hey�����|��س�T�c0�2��<m66�> ��W�� �5a?:�\$U{���穥��bMW�%�:OI��y[���]�ܖOg�@�wn�NS̗�����9?I2�+K���F;����.����`!y,�
b-�vQ-��L�`��vP�����Gr3s�B�:�kk��$�D�"���Ofn�Òm	��=��Bbs�;
�B��u��U�}k�:j�!4�u�@&C�E�S�>��u{97��E�Y���x8�H�c��EB�CX��r�?��Ztb�X�VO+���w����e�p��n��v���� �,"-b�e����p��y�L"�9��@�f)Z}.�_�n�(v?<��&g�j	tU��#��\�h*��($uy��][ׄ��,�?V�� 6DY�����,]UB��6��?µC�s[�r�N���m�vF�[�{��4�lݝ)n��<��FB��V��GZd��u�_�t/j���.�I�jh�����2dQi�Z��f؋���5"0�j�H�9T���[�G���$�$��7���!�7?8g���D(
5�H����.c��,Q�������۴�C�!�c&��G7fTK�����/q�3��Y6��Q��DG_�7��V�E�[K����I�yn�E3�;�J:�ڠu�R�4f��%��L�}��v)s�4j�ȒE�,^t�F'�R���jq���5�nC8f���j�;���g��^K�C�s�BH�{�؈�g�&Y0梨�q=yİf�8�3Ʃ���LΗE�Y�f�_I�8:i����D�q�ҽfVZz_I�V|V\o딒���uܨ��歮_���V�z��;���C'�<�o+ah0GRx��o�u���W������O�v=:T��[uP?����׿��������p<Kl"�Hۏ���xJ�}K�t/�(a�����z��Vbw����c�n4 p�z�I�t]vwI�':+ڳ��vH���\E�2��>��|xq�N�<<�ؐ��y4�֨" :?BH�͍c�x���β�V3�򜍇g*i�_���i��j��K�m�
�M��u�$�^y�U� �S3�d
��Q4>�W8�G	B�4/B2���Aڥ�jb��0A��3��@,����<4Š9\��D!� ��X�N(j��������V	(-R�(���Q�L5�: �rLmʤ��ܸ�xE����[����e�I�4��ݕ�ͻ��ܗ��پ$:c��`5���N�ky�:\��a6J'vb��@�RZ���#�L�B�V+��Q ��Y% ~��i���M ��d#�"
��3��	(��a�>�9��*�g�f�@�B�-;���K�f���D;��e�)⛥�X���K�+���A�2/5�������)��^���Ď�i�yZ�.�R�l����59ogO����+���nq�+*��%����3?��IE�MZ:Q�ľ��%U�AEF!�iz���j�%�m��6��	���ebR�B�R�"��\�&��ю79���Dpk$����'嵻.I�q+�/�]kP��n��$�:o��i`B�Q�y��CS�F��S�Φ��b�����H��2�\ñ� ��XGK�5�eH2���@Q�v{�d�`OAX�m;�g!X�����b.�b���/��ಇs����a��̸��b�6����g�fKEbx{#��F�°m��-q�;��D�?� u�I����ѩ�����e��ے6n�d�9�S�dmR��(�o�Lh3� jvL�"�'�=)ޠ���j�h-b�G�k�����E�;	�XY�颊�$�վ	]k� �׈m��:M"$���~"��&�2׬;%�ڳ��|t�`�k#�kJD��m��aR�X������=�!p��,N9�3�^���ŗ5/��1:!�µ��T�d���sG�z-�h�� OE�������|�_�&�%э	!Wܐ�z��&�ܘ�}��fv��5�2}]g�ͱ5-�E�
�t{p�8��r�rC�j�r|���Rq<"����A��u결ۊ��X��Lj3g״F��%�\3U�S+-J
"��hgP��^:夵��P�����	�q�k���HW;����ֹ�JY��,<e�Z��6�V|KQ�+ۜ��5�Ք1Y�䚓W�?��4��1\�/W��t��@
�j	b�S�Z��N��ݍ7��9H����z�ԹQ�r��L�0<��~���w�W?��G���wb����?	���p<� ���x��w�$<u�����`5�"�>d�L����C<��&<><�Ƕ���=7"�ӚO���#�� ��z�U�/0��XI�"
�G3����d�H���f5T�;HU�f�1�B�<�'Vg%�h��
 A@�L����}��V�+vq����G�j�l�H���i�'V\�i�%1��]��)�Z�]X-e}�ƯO�!tǞ�T����������d�h�iQ�V*��9����-�-걝&��,R=��~!�]/�ъKP���:9�5�>2�"N��C2]R�]ǦQ�� ��J\�r
�T4��-B
�u\Z�I��b��|
BIN��q��})��F�~9���u���d��B�+x�0u�agM��9.J���aBG;&R4��,����� �+x+*�!��
ZK�J[d��b��&��	tyd	x�`�J�g� o�@s�"��K3k����p>�z�O˅�'���b��e�(
�Ǫy~��o\���iب� b��ǟ�Ӌt�h��Y���q,Q*���]`���I%���*��?T{����!Ni/�1HE}pܷ���$�M�ϣ!�A���>_�����9���J'���X�i�#�3��Ƹ�����㬽J��2OgڏeX��)@�9�6"-�`�HZ6��p(F-z��.���qɋ�ӱK.��O�M��՗(t].��Rd�$O!��)��ޙ"��'�Ɖ"I�D����$�,j��sG��Ѐ7��k[����v���\�6o�1�`�GN��mޒ��9��dK� d8:!�&5�.�l�����.�+!kv�TjOS\�,ĲL�	���kKC��!�ϵ��uH�|Ŋ�m�:|�h���(�Dj$#��;�Ȟ�7j�>�_���,�{����c'Y'3BX�O���=�u|{f�Xɕ�f\��q?������Ș k�@�ǻ�Y26��E�2�̥�~#-�D����f.V�S�]�f�D��\�P� �����-0��v�L/���x�u������"õ�>��6��Z��0���-m�x�#YN�ג��V�	��uF���y"�s��p�T��׸FW6\�3'p��/�duQ�Г�9�L�u-��c�亅����3�ݚ�,6�Cf�,�w8�C+V��=�0c�(jʀ{���B~�B������,�ӡ�k�>i>��R]�Ι�Dq����K�[^Kq6^�3��1\WA6]#�ӱؽ�PH�	ν��Wu��5ͺ�E�����<�q�)�0>+����AW葂�ډ����k���qcNX�5�yEE�V�D���xy��kB�ϬE ,ؘY%��x���y����n��gA��"y?�Y����6x��a:�t��:�)�c��%��e��'�~��t��{߬[��/�׿�{��p8�?.�8��Y�D)����Z��)�f��/ٞ�!����T�.R���R�n���p�<��^���x}}���fi3��*�C����r��{��}�%�?�������EA�JXw��/������`j��!�&�f1+���(�3��N���S{�ʾ(����AѨ'��h�4T"4XHѠ��aj�a�3*K��~�����#��׃d�D%��(R�i�9���+�:��BT�\T-CXB�~��ִFAyz� ᨼA�D�P_���Z!�[e�����*Ƹf	$��]8��P�TQ�t�c���rt�Ƕ�c �x�g
Cm���؉]�8��4�$R<�ԕ��P��c[�H
�$!�s��b+Sh����Y'�,�>������U�UU`7�9��s�@��GQL�����\�T��P�Ԧ�gVD���Y�4�]#�Ӷ��.�-hق��f�ߓ\��~�|�O��M$�f�0b�~��tH�h�9�

2T�y�j�5��xzK2?�
�ڡ�IC�1'Z�8��̳�"�%H�q����%� �p>b�@�QN�*�k#i�A'�Xk�L�e�`q�����l�!X�b�y�mZ@����.+喪c���sE,���
��,��� ��ӈ�k� 
�J�K��VxC�]��!2B�[
6���g�ωB��gf�4zRG!:�t@�~L:���X����</�̇��Ơ�y+�鸣�N��i�<.���<��9�!������N�G�a�� #D������W3���O�J�1Gn�B�X��y�ѵFn[���9�e�	;:�CX�@Bs�l$$�]U�]5'9�2� 9wU���.�cHr'(@Ơ]U�eN�XQ�-�%d�)��8
:ff�r͛՚�(���iaY5���5�:_�"f���P�boA�At	r���縬�L��s���V�QΛ6�"�k�(�5���z��4�~@�5I��Z!�a�GQ����)ۂ�vS�]�A�?C����Q%�ޫp��o�}©�i�S�>�"xs̋
ᘤ�Zx� ֞��'�Q�F23�	r}������H�*�KL}!��i)������q"v���D��u���t��t��Z�3Y��"������ڢd~�>�P�����h�uB:,$ ^��"�ĲF,#!���;\���%u>4�e�U'�?�ۄ��`���'^�Y�!6`&:��g�I�I�v���e�8O�RAn�,ϣv7\WpN����Z�s	oŵ?����U��{��$6��/X�-��wݻQ�Ѻ�?�u�sb,l
'�9�L0Z�a!�J���R<�u�W�X���+���d��Ӑxܛ��u}����	Kn��y<����tz��{��˧�~X�;���V=Ͽ]�������{;w8ǟ	@����a"ȡ>����QC_�z���{��y~����Cf��'T>�V[KȩdY�saUd��*քZ���$@�� �l�J�`�3m����}�`gxѧ ���v��:T<��!B�qP~���k ��II�^�rb0qB�}j�9�և��@���{x{��	�v�`s���L��M|<��!?&�u"� ������<��!�ʌ}��&01zY}����3�qg��*�F����vD!���-4�3@ٱz��0l��B=�E���\���ˇX�_�����0K�B�uɈ��ص�+����x����&NR�0��U$#��v��t_���s���6��$��HS�TSFf"y.Ӭ��F�����'k�m������c�e�"�� �ER��ܘ��C�G�T�t�5 'A�vo����
�bU�(�K4���)Ě���B�� q����U�nį���s��Z��������V�լ5��>gV�n���ξ~���2�	�I�2�0K0�������W?��B&I�����1g:~V1���H��0�Q�&�b�X�()���II�v��I�Ͱ��3j�
�:�P�u�A���YN�"�O]�]#QE�E*�!R�|e�=ǹa�-�8O�>���|���:OA4!t!شڱ���q�.��Y���,�����?����;�����]�ӑ۲��'��<�5�U�*<˚"]T����ct���g�đND�^©~�	E|��|��Է�_p�J�pl�M �q��Vo�q�zV�� D'�i��#|�#;�@ ���=`M�X2%�!����N�����d?�ܔEԡ��(� ����*"��ǋ�O ܥ�_�1�9Q�9�ڶh�;�Ñ�d��ga#��)���"��4��%��� @9�z���K�D%;��q�'���WQҸ��z���$/�vT쨛y��/P�K���u�n�΍	�f�E[�/���Cc��)V��4O�z�U��������r��)R�X�"���Z�5m/ǋt�0#g;�)�b\ x]�u��	�V�/D~ԮH��ՒX˵�y��_�\jꚅ��*IF�v D�yD(5O��"Y"E�~;/E\��K�o����!��_"Y!֝e����/g�Q:����{��?��fɪ�y���Vq.K{)����|E��-�t�"GYˁb'�u��3L[�����Fr����%��P���v�H	֠�ݥ�_b�yۜ�E�s���v��簛�[�*2%)ؐ��\3LLcD_Z��*d�=JL�i!?E��<��`w�X���i^�ն������@�nx��"�Qރ�6��zOZ�9��]�g�7�Ћ}Ϋ�2Ql�!��+�b�
r�����B�1\$��|b��k&��m��h�z��8Ab�?�u�^5Sy�/��6�O��<�?l���Ӝ?���/��_��?	���p�_����p|!`"H&WW��rYJ���8~�>$�W��в1�g�v�Ʀ>��enc)�,E��p�'�@b��v�����<���XX�F����K+vU���u}�� ���ͧ����7ǻp��-	O<$��1��~��~���t�V�oAh���-�J�C2,����\�'XrL1L�,�lS[ ր�<�j^�<Ȱ�(��YmV@�B�aHu-���A���:J���$M$����I 7��9�`���}\�TA0�C��ԓ\�eJ+� +:g�&:]�$nOK�Vl����y"�\%A��Y0k�A�V�S��E�� $��yg�2���"�8h�9˱��&�$0KV���
ڴ�A��9®�EB�c{�� ����+�x(�Dj�Z�hz� d`�Ih�����ة�3f�M�PG�����OunÑ��b)T
T��,�M�0)d�X�~�%������Q��"$>H�	�ǖ�B/�kOP��Aʴ皥:v^�,GT�֭8��4����!˭t�$a����p�a7E���G8������6'M�N��Q(/J�1�&{�ma�x5���͋ڃD��0
�^ �SQ��)�@�	�e,Qh͆��ٱ-A�ᥒ�Aª&H��P��R�VD�{�X��f�b]!�%*�����X�X�*�G�ó�w̕v����A���5!�A�5$��r;䝽���L�����s"㚑�����Z��ΌU�W��ԉ��i�BPn�$�e6�{�Q���IDMɚQK�E�J֬ �%*�6���8�"0��*'f:I��睺-���h��G��F�� ��I�@$�@Ò�����I��'2�j�q��R�+�&-� �I|8�(�aX�R���H�K�EDew���V�$��|���,der���<�ʰ���v,����m�)D4:�b���S�53p,<L\��:�0���^m�γ�"�������m
��:�ύM$jK(VD�@KI;��N��I���~˼�$BR�9K�V��K(�����W���1�?���`���E������5x�p� [A��Y{�!��"�$i�9�7�	(�2�j,d[�͍X�%������D�E��r����5��	���z�qww
�S��\�!l۟X�ϗ�vR�/QE`�����9tK����Q�
�:��|%0�j�RT�� @KV��[,�,qތg
�4���uNj�6\�0��CN7�Ն�?���X��� �V���x߾��Ya��:׹������b����{S?����[m�6�9��\�ږ�[��	*���LCzY�ӑ�z����A��B^sP� �?���Ϝ�2���輁x����I��'�-��ҼMm$�	��8^��S�)fӅ��;�v]�&zvR��Ů��,�rY�zQ��?�p֮8��	�����<o��v�\���<�>�-��u:~Xw�G�C^���~ݧK�^�}��W����p8��M� �p8�/V;�R�Q^�������	����y���Ǯ��2��������>~w9��c�M����y��s��ж�e�kƦ�Fl�c��&���:I�}��x���<�w��w_և���pOr����=p�<�}yjţ��4+�_����;����$��=��Ϲn�2�te)��ۇ��2ڔ��5Ҧ���C�حb�xS�?#h�ɓ�m%�mJ��l�+�����$�	R�]��j��@<
�/��6Ooa��A2U��~�"����r{lE�н�|�%D�H�+/�ǆf%�GiPd��nAč������A�'|�BW�m t�Wj|��|�A���"i�z���2G��~�e}m`���I�HvC�)u�7��th�sHC�ž;`�q��:?�����:��~Ʈ��פ&�ɋ!�٭2���-I�:�1��̒�aX���,}/��m�}:Cl�>&VXk��u�b��y���m��1���<���2�>Փ�Y�Lm�wO!4%�o)eYrJ˒�~ICGΑfJx��CwmBp�%��M��ܭ6&@?dV�r6o�OI��$��7�1�PƁ���Ts�fe�8	3��]�@���- �!��������-M��%�ݨ�%�.lL@gE��9���[;��<��v��1�� �S�핐o�@���,V{&|d�V�S1��>u�4jK3>h]d^~����r��G^�:Z�%��K��?p�L�0$Uۢ����$7EB����4� ��W���e�qz �i��h/�X�ⱨp6��N���J�(�+I���B�ob��U�(�ZІS�'�\G����w�v%�v���.��[n�HG��v��<\���lBKT������)��ƒ9��z�[�
Q��dv���h� ����]Q}��_��R�t��uT���)�I��B���K�$E��5�o�����:�ކ{���8�[d�4$�c[@�~�8��s�b�e)뼁l����335�
�I:�����NO�.�7K�A�hf~�}�$���V���o�JH�9��:?��	1⇊��H�v4yͼB��j�aw��.��h�F���f   UIDAT�0mc�c�]Am"�Eϼ��H�

��ƹ|��fq<�������')�5��BE�4��<^hi�.)t�����G�<���u,��9��ϗ�s�,�u7�^@H��"-?[`uڬւ��ީ��9����X���_�r�4�N��C8�������m�r��;�z��y�f�R����s���&�}+!䷷��ɫ��<?����^���Q��ZE��5�f���Ō��=����2�`���pY�ք��O��#.un�*�c�Kf�a�8*EQ�246�|V���@Q�����q<���Gt�Mr�G!���k�s����p)�}���@�x���S�]��ۻc�~��0.}y]���<�?����t��.��ވ���p_����;����p8�?'\ q8�
"�����K����겯ԇ����֗��;];ܞ��a�s_:��]�lK�\@9��` r�9�1�s}�,�: e��2�(���"c�A���|xl>�nN���-��N}���K��Hq(:'0����Qm�c��)����VS��
)����X6߾}�><�Ǉs}0MH#��Wy�qn��]�{M�� ����?��
��~dP�������O��qZI`�����?��F�>D�Jج<ql����]
X�� .�
��v$k�n � PLx/lT��Cn�dU��a5��I����6����el��AP�^q�u���j��+>U����������t�q�W=�A����p�v۶!�쳃��HeD�� ����Dd��/q	]�X]Ώ�M|�q��k�n�/�y��9�]=� ��R�\�e8〚�ˌ��~��C?�kOǃ��Pȱ���1��eߎ�i.�����Z75]����þ~���6��|~77�ܠ�t��pO�y��q���_�w��1��y��"]��s#�r�s=�/c����0�2�������^�BP��F:�����Hן4t>��z� �;$5,/nӑ�w��c.��Ŏ���/�E"�;�5=��Rw������,���r�:/�t8���+yB�^������ݩ�nH�=`�r�$#߾U 3��Y�d�&8���Z���e��;�]JL,Pa���&{�l���5�bH�}s{��߇:�(�0'E9��=���y:׵�,����
�����Rǥ�q�J���D�@����"-�����0*��Q&	p�_��Wc�7�A4�^~.�eN�&�S��b2I�0�Ȳ{=:!�N�&�)n�IF�6&�v��p-����
5��	��3�g�Ť�y:���Cך����Y��+@��B��B7��nߓ���1o������]���ݛ�����;/p����{�Z
ک��=�����k�|�D�o�)�O�sdY&%��f#Y�#ę�Z�\P[��X�m�/�����Y�� j4҉'�Is�3���Yx-o[�ӝ������/݅v����B���H��ޜ�
/.J�	̎r��hτn}�?ş���uN�Z� �A�_�qG��&̉ k!��G�N,�[����m<�!�1#d���ڃE\��	�l	�	Lg�U��O�+�P0@�D�-���\�Gvs�=�H�Z	K˛;���˻�ӟ���|�ɫ����������(�ys�πM�\�m�]�-Vg�I�;(ZK�<�н�|܋	�G���[��;U��&�;d��_33�E�)Э�N��/�eTx�6����z{�|�uF�'j{9��\�v���vZƺ���	m~���8�&�n1�m�^��>�mKx����]s�7 ��q�q�w���S��ay�?��}78����.�8���_��o�I��O����G�>��(��K�i��9���&�7���<S��w7w7��_����Ԉ�В��!�ݛR���O�1�����	�b>����T�����)�ܗ�t	�4�����Gz����~�j��m|��'��HPl{nNZ�
2i�����VY	<<>��*�ܞ�����~����O�Bw�(���@[����M���4��0����mz���V*Y*�gM�HR�<k5a�����+�&!֬Z�b�Uq�1�����Q�T����C8M���G?����Ϗ�D��_���Po�,b��::�]�tɟ ��Y�4�q��a<?s�<^B7�x���~�A���V�̚��<>yy��=cm���X>C�Ai�����{�ׯ~�O�t�x7�� &�X��P����z<��K���(�N�C_�U��ۀ�x]�c(ǻ��$Fno�Ǐ޼������c�w�a8��R?#6yٔ��ေ[�w��0<,K~�v�C�܏�2�n*i�����Sl��6,�:=�<M(Eɺ��q�.��:�ĶyXƙs)�I���[N��v#3)�����<չxގ���Y���>�}hv�O˞��w���S����W���85��zOz���,Qۜ7����2iT����>^m������4��Ʉ��(��s~ה�I���E��kl=M��ل�F>��;u�ݿ��<��k���ɂ~A"C	!z��Dk�F�j��@�7>�C�����e��S2R�T|�0g�6l�P�_Ϗ����d�6Ql�g�['�Ǣ�_���I��E�V3��u���w��b���"��4/WoX��v;���N3���:d,tڥ������{��5TDȶ?���:���d��~D~�v�|��~n
=D���\=~l��\�W��pC,�;�~�vr��gv���~�c��K\i����/�ڼ%� 6�&N���r�n��E?���5׶�V[�	y������E��e7>�ަ�0��O�0��2�����u�l�^�L!XwM�Y��v�T�y��DZQ��à"H���S���b"�5Q�G���K+,�������涞ܔۗ�B���%�?چR`F��(9 �'?yl���?���2�n���^W���lH��7��1e]`֍a���ʩ)ֈ���17��xk(�T���/z>���לf]���=Y��:q��<����*6�
h�|[���܀^�&Bk,��kǎ�Cwi'��o�m#�Jc]��ֵ���W�>����[����p�����p|a�����������ȱ�K~���E}ʼ��x��㛇7w���e��E��O�B��y�������pI!-�1��ahJ*C�>徬���=C}�o�������r�DkX|\��{��U'l-@(���Æ���_�����E�9h!�N����u�U�}��_?���i������o��2-�ۘ�%���U	��8�n�S��i�)�s�fǌ�Y��S�o�z�o����g�at�J�
�=���L;�*]?���=!�r~{&i����y�z]��o@Y����L+�WbE���w��@۝�j�� O�)�c�;
����f0�q���X��?���J���Է�����4�ѹ-r_J��?�I��k��z^�����(�|[?��<��Ss\���M��ˮM����tlr.tđPW&��P繞NS�������x<t��8�^��J}Osu�K)]�.u�^@����O>z���=(Ӕǹ��|�&�^��r�J�0��)�ڶ~�å=�o�|R?�mA��%�@�&h��l�Z��o�'��F�+�����mR�ݮHr��o;0����&f���J�Rȫ�P��Y!�Y�1r�9��T|,���i���¦ttH�!��o�E{KK��!�O({��i��u�$u��X�	�F���|"���z�X��x
��v��-��a9b5�Nf��jP�`��v�H��fM�F�b��21�5�ò:$��
���\��:�bپ�>{.�2�n��FxE�F�XѶmk|"@	y/�5r�����\!��-�7��a�����������X���<���y|��;��*�]�o�a��g�R
��K��������� �g���^�Q�E��+����|�VŃ�k�!����;Ib��~/��--<fbs$�2.i������]�ٚE�_?O_���wc�9N�$�9m����^`�e�#�gC��UD���}�}�u���x^�G�K)�hWc��s��5�,�8O���~I���3ˇ:��ȉ���m8��'��v�iz~z2��O���{�S�,��p��vЮ��3&�׎�OW��_Y� �$&��
�d{��U�ֵf=�ȝ��_�߰N�uSiɶ\��>���.2�L�Yɒ�6Û+az���M�y�7?�c���v����}�]P}�s=�C��\�豴��������p8��`� �p8�/<���O��?����eY]��c}]�9��]L�1�#܇��,�XJz�Sx��q���by��
�!7�1�%�����2|�za�+�dTwH�����Q��s���N��ӄ��6|�g~��y�v���f�����a8�8��ˇ7�o��>���R�6�,k�'����5�q�oS��:Ӿ�`�kjh/���`$�Ɛe��	;���x��5���ϒ��F�M���������\�9��z[$��8��h��8i������(!r�:F!lO�c��	��G�|<}]�aE'?�˓�M,�j'd����_ӿ����>�p�[y7���0�A�!>�о���@
��_>�M�˱�JH=��R�n�i�I�	��cҗ��3u��K�(�O���O!��]��-��r�5�8]����{�=�|�b����������>�|�3䮾�,�?����1��PRyS���<�4�u��҄�5�<)�B~>�%���n<���t��嫺��k������;�6Z��ϛ�� �N �l�y Ȋ�g^�MB����  �j�����q�]����9l,��1�V�l���e}�5A�t�I?�d�O��	�)��z#ש�;m���Ov[~��X���V��p]ڂ��}r�����A���֭ue;s{M̟�Zw�-��]wƾ����\�'S�O~ik��q�M�티T<Yo����'!�m��mw�8�b�}���ã|�m]���.���}��zv��\�52����u�=yyBP�ۗK\��ۺ��x�ws�xd]��-_�9G��y��8�5;�3�aa7a���^���G{����5j���K���Q����d��ܡ: ��C�NM�G�\�,PvM�qY��>oޮ�un�~7�ל0�mM�^�l�b�}�3�s�~�❟�7�����	�{��z��c{ѵ�	l.�{���/}I���+&F���Ӯ����z���F��[kK�&��f�+��;����-t�S��s.o�M���L�g�O�`�:�AW��sY�1���������p8������p8��/�w?x������e��%徉%-M�s����~�w?��g��|�[ʐK�c����\��p�M����&*�(��Y	���{����_�������]����Ż�'���{e�Ϥ?���W�8�{�/��k������?������?���a�����х�T�8]~���u���zn4�)��-e��m�y��TR�0��1��~�_��ݿ�����;�o5H�t��]��e��b�4} s�c=�.���3�ۍ�\.=����8G�u�yJe\������7|�;����p8_<� �p8ǟ�_����s�����ߐ���Ͽ��H�yı����x�_����/�\qQ��p8���p8�@���p8���p8���p<;� �p8���p8���p8�������p8���p8���p8�.�8���p8���p8���xvp��p8���p8���p8ǳ� ���p8���p8���p8�\ q8���p8���p8��������p8���p8���p8�g@���p8���p8���p<;� �p8���p8���p8�������p8���p8���p8�.�8���p8���p8���xvp��p8���p8���p8ǳ� ���p8���p8���p8�\ q8���p8���p8��������p8���p8���p8�g@���p8���p8���p<;� �p8���p8���p8�������p8���p8���p8�.�8���p8���p8���xvp��p8���p8���p8ǳ� ���p8���p8���p8�\ q8���p8���p8��������p8���p8���p8�g@���p8���p8���p<;� �p8���p8���p8�������p8���p8���p8�.�8���p8���p8���xvp��p8���p8���p8ǳ� ���p8���p8���p8�\ q8���p8���p8��������p8���p8���p8�g@���p8���p8���p<;� �p8���p8���p8�������p8���p8���p8�.�8���p8���p8���xvp��p8���p8���p8ǳ� ���p8���p8���p8�\ q8���p8���p8��������p8���p8���p8�g@���p8���p8���p<;� �p8���p8���p8�������p8���p8���p8�.�8���p8���p8���xvp��p8���p���ف   � �{|�  ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `G�      ;     �      ��      v     �#@     �     �     `'�u��2FNt    IEND�B`�PK
     ˡ�Z,�ln/  n/  /   images/6590c6c2-4084-4043-8677-a67706af7572.png�PNG

   IHDR   d   d   p�T   gAMA  ���a   	pHYs    ��~�  /IDATx��}�egu�w�}9w�a�{�tO�Q@(����0���x1��m�1��e�kmo*c�׬q���B�
���(MN=3=�9w��~9ߴ��z$�Vmm�t�Q��S=�����}�������uM�����u�\c�:C��u�!�غΐkl]g�5��3�[�r������5ǐ��I�Ue��Jr�����\�pq_��_#����(T+�@Q�����`������
�f��å���f��k(�a�
=O?.�U����0�5â#@� �Z��ܾǇ��ܑaG��υ!����M���"R�4��.7�E� "�˄��x�7��/�����2�T�P�}U�zWO;��n?q3KKPuLŦ����i�<����j�r�4b�%?���
��"f�*1�?�EL�@���s
��xQ�*x��$2�2n?�/s�)�3��[��T,��D����nbB���I�����BTeZ.��ۣz}����*�e�y\D�*I���2֒ds�!�J��#,���d�Z���rYmPLb�K^1���s�Ę0C�)<�`�bi��q�,��N�:�`j�K�K��N�s;��0<���gH)�%�y��j(���x���h��2I�.��i��9$SkHgW�4�w0����!����q�; AL�[X���V�2"E,�f��&�}na�E��Ǫj���V��Gb5��/�fK��B���r�,Qk�H��z?����*��1z9�&fQ��~;_��Xq��˪�
/]�Z!&d��*r�=΂��O�Lh��ͪĂ��A������3��v�N��B�D�.�$�Љ�FM%�(1�YmK����B�^z��.E6ȋ`0�P8@��lF�Nq{}(��fz�72s37����N��q�+e�e3\V=�e}�*��[�l��EP�c��*ӈ$BG*�GWW'r�,mJ�Ev����Rk6��/˄�H؆�MAV=|,�����9�O�c�*��Ѫ�<1L�������!��}Ii�$�Tɜ���u��������!2t����0��DL�] ��
}I�� R�����?�����'1����	}ش��$������JL`:�*�R��0���ϱd�U�B	4�Itf۶��a���a�v{��԰�1C}>��r�!Aw����,�f�e%u��TG��#��N�eЮ7�xdh��W�����>�(�(��f(r>�o�Ȓ�����s�Š���aK(�5�*r6J�2]�%�'L�l�J�U1��1_)�,���W��r�!� @�C�ƅى*i7=�җ�`����hAc]~��Uqrt,%V1�1,*K7�Ц�T��6mqaPUנ�.��=�o��yf�a3���m�!��X"!�H���>x�icc�d����j+�Kr3��>�������b�|�Ff���^�3'��+���d���kXIe1�};N�<IG�
S������/aan�F�աP�����6���jʑ������c�Z���#]�b�ĉTY씸�.����j�bD�5��G���x�7~�s�x�����?��C���������m۷�$9�{�IG��8C��[��>O�;h�H�N��{����ԩ�Bl�����8Dؑ�%�8xpF�&���IT�Z2��|�H���*l�}>|��$�C���Z_��g���2�� �������zD�F�+S(Y^�6�7^���R�����5cvv�rA��g�n�@�����遏<���v�>}
͍��GIm���(�w��!	Ɏ�PH�L�)><�����������S��M^QI��l��b��|Y��xu��A����M�ؿ{z��z���6eb��ʟ�C�RD��]a��ax�~�'�yb�Y��HZ<hhl[�ku��=�R�1z9ΐW^|�L+˳(�*عk�kh�lC���i�ֺ�:�J ٢�"Y�n�� J^O*�!;�p�Iv�@�!퇖�V�
u�E�p�m&e)�r> ���ٟ\.KGv��	��m|�8�$�X-!�� �#�x<��@�"���ة�",c㘚�#�aej���Ʃ�8C�ZZP�*ؾ� �V���R�E��n�|����:N?�Ζ:^ş���K89|����Ɩ*�)��:b�	�ŏG<�+��Dĭ#U�/�!��n�ȕ.�U��'�`El��ٙY���g�c��K��	��z��O��s#D�ޖ�[���Eck��z������E��y� J�>fg�p/ِJ��'�~Iډ�_v���4�����CG!�"�Y��޻��'��zq�'?�썟0������m�Г�s	��*b�<�'��-eQ?n�W�ɻ_�+t,��ٴ y��B	�\�h���	���gg?>������b|j
�v�@kc�%N�C�q���\���.����0hg�/�i���(�a��Rl΁EVIC[7�o�5���q��KR�*'�I�$�HG�q��l��btz�zb�J�jaRiyR5a�f�!�1�1L0Bww7V�V�gH��I%6����[o$G�	���lQ	�x����]n�ml��dd{{¤���.���`n~�m�Hg&���;��*`N��w6�{&�K��*I�eE*��0م<ٖ<���*:.������Ebf:c�)�Bq|��
��8#M�'�g<t>r���8L�Eۆ���!�1�sKK����E X��sg�6�������-}�8}�5�!I\� �~�HB��%��`o���������Hj�`�,J,�ǁ�X4�8�|8��Bz-	T�#���e�$���^�D�dw�>7Pb�U�
�i!w~a�J�~4������Թ�H�Ӥ�H-r�����AH�����5\�8�O|�N�u�193C꧊j��zB��L�7s�-6߄�9BLh��Ԉ�c{S*=�"B���hi��^/�����ο0���&��J-9eH����q�8����z�$�����h���ؑ�b���������Z�7X��c�^�����Ѩ,'�IC���Ս�{��::~���(�H9=�*��"©�,�α)-���Je��eB�F�1�XF}(/pyu���̸&���Q�$�؆��P��P ×�q�����$�!���OWG+��,����q���Fcs=Μ9���mJO{����>��#�r�!=p����o.&HsJthh;.�N�*� ����xT�+v��%au��� 9/�.N\5�¸�x��^�"NA�v9g9.�@�]B���S�KE�K,咆PЋ���hȋRoAbR.[ j�;͌� ���.F�وIgI\CS�"�F���Y[H`z�\^�_��/,aaz��nA$!�֔��!����F�b�kIT�v���<o����R���f<��IR_9#~�Sy�'�0!�
�$Q��>��� W�����%6tp������Bss����Ŭ0olj���p��cq9����KQ+nU�S�y�N�K��i�ĥ�H��4�Ņy�����t��P`�L�D�P�����eưT(5��&���q]S܎�rw޺�7����`�Ɔ���t�@�B'ύ�1K�U+�Ph#t�7�c��I��VEjtݒ
K%�YX����oh���
"^���c�r�!���/�����k��QR>2�v8�w2G]Y�47��d!��s&��9l�E\���P��'g��|���d���v|�pG� yT>6غD�1�ё=��^�V��#�T���-p���v�3��.��7H��q�����j��}�x<�������n!-�3�UQImd47nގƦf{�U,-/
Ay���^Q�j4M��j'��Ԧ�Vh�4\U����($FF�%{R�a���u3E����
���?H�jمtl[s�d�I���=v��/�����f�������Iv�v��o���H�C�q���u򻣻�t{ ��w�A]C�++�f�~0�Y*\�m�DX�^��Kݖ]����y/�6�JgQ]!��s֡JF��)�J�G'է+!�Z#�X1�o�ڸ��W��q{��/�|�.�_-���H-�P���-mm2�xC����,�m����P5��ө�/^BSK�)��&���z���͑\�bHqA8H:ݭ������!�"`x�'��i|�4�?��MOLR�\�R*P<A�NQ�DpN��a^}�f����Ӎ`0L��`o
�]՘X���(��Cs�(����\\��r�!��y�=;5F_҇�g/����A��&��*\�A��v��܅�gƱ����nBSC��*]\_��d�u�(�.{P���"t�����&)~0�%",yVFA����8���ۭiq�����|����#[ƿ���"A��U�L���O��*.����!H���̐޾�8qr�z��ݰ/z�6q�G_;"�bt���8z�,��&�GTl�n'Iǻ�HA�V��d�]�$0I��F��ǀt��&u�vK��!I�&���Ԋ�y>:�@NA1�!/m�)F�����rᲠ�xw��6���c��e��w�rITڡ��9B/������ې^Kc��!�oކ$yY㣗$ X)W�T'��m����X\�I�6�J��0��C��l4O:G!���'"��\��]:�,9Z.���e�g�5���IR������6�dC���|� H���"p`�@�jjk�ѻ��"�j�oc�wnfV~ɖDbQ̌^D��r�C}y1DC< )Ѱu�F\�N�c����I�iIү:z��0��'���	4�x��Ȯ�+$o��Ly�v�j	FI���Ru,�$a��?r���><��s��:hC$��e��Yt��t.�	���+�XXZC��vl�*y��ϥ��DjG�@�ӧ���!C_v�$���첖��ߏ?�˿��H�1v�*욡=����صs>���o��zX����`�H3KB��0�ƕ�9T�A��V��Ձ�
ٳ���Ǘ������Z#�=0.-e�}��O�*���$<2�ζV��;�gg^K�s��{���$�E�\��5��H�JHe
�����~bǨ��+B�QR$7l�r*���F�(^b�������[�T���ydW019-�.��D�RI$�Yd�$G�����FHu��b~a�����1|��T/&	��ip,lz|O����r��Z�L��;��k�l6�L:�-�����X!;�L&���9`�+h�j6B�L?��5R6j"�H��+p�J!5Tq�T��☘>G�!uF��A����>�%�e�!Oap�ɳ��? ���M2���q���K����w�q��!�ON��g >nc�L��]G��8Cؘg�c���Up��^��u �vRO<�<�r��NHZ75	_U%�M=ܓÿ9���*yI+$eem
��M��l���aF��x�"X���s!��a*�A�T�����p�?�-;vI r%��S'��{��{.W��IȾ={08�/y��~TK���ͷ)C�C�0�h}�;a�\�/�&hjj\�C\��;������\��g! G~U�D}� �I�%��r�58��y�X����xy�*v�݇��f�M�cۖ������?�b��={w�R��]Cs{���=�	���30>ٶ7f���p{�S�q��k�jݨ���a��0��e��S���,��9lVMm����q	�H�J��Щ"-� �@8Bv��j�+W���^�Q: \K$��&�V�y�n�EL�]I��0Nj*	����T�46mF:�Ҥቧ#W���/���p�"J�\T�t�^px�	�^�<Aī`yq	SXJdE����l�9!��݋��.��K���8y򌨏���#w������]h�oƳ/����46�e�e�$;��a�Ǖ�*;g:m��X!Ɲ=���\u�l{��Nnl6�B*�&��d�C��Dz�d��y�y��8ټ����J�yЯ��T�BS��x.bq~��z�=��bx��B�v �0�("�������y��'PȦQO���}zѻa#戱ym�Z.H*��R9�-5��j$dXH��(��߲�uC��g��v����:�~�]�\�s�.��L�}B��v�7�����ߋr��ϟBG�2yQ�x�UG��|�܆~d�8�:�n���H}���[nó�='�A����2ȧ�bjl���g���C8v���F.����?�ݿm�,���Z�JT?4�.��
{��ڭm�l�������n�� ��Vc�<P��ťb�a,�- J���g�#�c;Ii[7m¦�n4�u#�[��[��Y5��W��z9��}�����_�EgwB�fN�>� 6�Z��7��x�>��~_�r"I;]���֦����-��>��Z��ns���e����]h���"Rv�$��M���y��/��/��<��ϟCo�^i��"�IbR��~qn
'O#i2�=�|��\u2M�/�Mq������[�"]^���(=� ��Uw����2����";�`���U��+��U��6å�w�cN2�"���R녷����8�7��l��`�d��G� �M7�"P���ˣ��7�A�b� ��p��ӌ�t�^�3�������c
�?>��A@�hW+vw�fJ/;��p������>�r�G&'�%t���V6���#{�|<��m���&�q��Z\�6���3
�ً�`rz
���᝷݁Db���=ȗr�J�|WHrn�\6���v�a�֩�����~�-���C�����>,�r�j����3x�;n@[G^{����	X+s�x�R�0���<����Ip=�}��֬uۊr���Zg�z����5�Z��ê�(P�X^N ������f��	��|	ݝM�}x��7���7��~����� g;;����YZY�i�Ȗ�`$���n'��8��s��R\dh��K���>��<R�.P���SjiV�o)/��;K�$����R�O��ضȰzji�D �����U����ގյ"��^������M��n�fr�V��x�z9ΐ��v�^� P�SVk87<B��͍M8q�u�l�T'I^P#y;C���ы4!nX6�ڕ�5k�au�'�q^OZ�c`֪UT���ikJ�j�cJ���=b��^����on�Hm������T�LH{�*Μ=�+Wf�e�J�h��/�q�����	�X^Z%���K/=���:���d~	W�t�ԡB:�s��a�6|�Ͼ$I!����l��iv
j��ƚ�8�%M�eQL^�U��R�v���z+5��������574�}�i���}�0͒tp-������hmm��G����,�n����3�ë�1��}�|�~,�N�.�0=����V�i!lP�v�S�'`T���/�!n�t�0�\�C�Y���gfF�6TF��/K�K��R9�g�p��{]��b�Vqt�`�'�q�R#�83���*斤.��>�]C[Ib;��D8���v|��ns�^�3$���!n��"�0�Vh����}/6�����^��]�͕̜(��2���ftv4�J2e�3�@ӫ�iIu�aG����{I'x=v���߸ȁ�W��ļ��Y�n�#�Ƕ¥�)���ގ]{�p`� ~��#����Bn����~��󥤤�wҗ����f̳M�6���{�f&�15��FB�W���:����"u���������V����֚3��R�m_L<0N y<Lx�Fl�kxŰ�g�gR�Q�ϟ���0x}�����m��$�ŅKW����+�IF.^A![�
��/<�?������r�!L�kJ[B�.���\{ZB\+�uZ�o_Z�V)K-O�y��'�[����@y�_V�0�F��]e��#}j-�x_����TI���>���E^�3S�p�y?z�1����ȅ׼~�}X�X�ǲ�:�é��c$�K	ّ���`P��"�RL�8����cS�a��0��	��Zw���yg�!of��~�1�Gvl�kG���
�&!��ǁ�j��Bسk�M�s�?�����8C2�,B�!��� *�2ؿ���.z�Y��p����Mo���O��(�S|�7���P�zi����0�:q���[W���͇��c�.{ �/6G�x��>Mj�,��������O�'6�{��}8w�m:Z��'^�x�cx��c�E�����>����>L�^��˗q۝w����ˇeǲ����j��JtE�F��]v�W*-\�R� ��b|�l�I,��#�x���y�d�R�U�a,F����xbi�pR]��2,G���lfE'���U:��Ω̪bo�ş�L��@�/���o��'�S��N�=�'�x�$����ބ���[�<�H��}�}�2���kvM�ᖴ����KK��+��yRF�6���6
�x��ll߽���w��.lݱ�������7��#Ĝ%��!m��0wnu�^�3��������0�����]���)��<!�"z:ڱ�LI)�B"�\�B8�?��Ћ/���Q��|� �V*d�C4s�s�0aJ�Q���c8.��I�U��&$Y�O��#?}	���'�
��+�HB�L�?�w/"�q@�#*���ك��~���YE�������J9���(��j�B�B�����w#�؈��2y�Qy{a�������K��Gޖ�l�QE���rD�[�5rA�)�= Vw,95�n��
¤�pr���R���]ظi��_���D#���v��I��1�'��蜍(�U�~�queQ8ӫ�8CI�زkK�W�5�	,r�#@��uu𓫹��,��X4%�n!C���w܊" ��xP*���rª�O�XN"�Ѐ��R.atz	n��ٵg/1���a��*7���a�ҫ*�����G��� ��&t� y{���2��Z�=�L��̽�3��ӎ���bk��B� �,*�b�BA@�֡](fS�HWO�d9�+�kld���(bqaV�>B��XJx�����Re�{q��[ۚ%b|��X\^���ARo)��~,&��ԓ��K��^Q.b {��cn�koiBwg�t����5Jz#��F@_�g���cG~�k��ܨ#��9L��P���w)�+J�Չ��0>5+�p��ēO���f�C^��E	Җ�%l��ơ�'�;nǡÇq�-��"՛�?|w�}N�<���f�hC�BA�{.01t��>,r;6����Tʵ_��ä:����Id�L�	��j,�b�� ?`��E�2�p,I��>V�H�b�z9�1�+�	��D�Jy3�����:ې�N.�oo���p�2����SO�34����T�?�4�:����8{�(*�*�F#����N��C��,1V�J܋��g��=��Q�+2���-��o ��?��O�*��Ã˪�W2� }�@�Ǩ�$~��_v�^�3�R��rrW�Kv.�6�P��=v\��brU|�5+p �#����p��El܆�'N`p�6,�O#ܽ���,��"��(6E���KG�Z�C�{p�ͷ��N���
,r(�3�2�@��c�{��KHW�n�����9nttt`jjZ
+��ߋ+����Io���GZHrg/���{��1$$^���'���VxSn���5��!���U��,Ue�L:_�*����f
��ޝ�;}��P���q�����f/�IJ�)�X"��/��*���讝ֵ�뢯^�kpk7��7��E�?~�Tg��ΜCs}�{���أ?�[+F-bb},��g�nJq�GU�6��]6q-�"�P�
������v&ߊ��s�L���#W�Ð�U��F�e@W���}&������Yx|���-{�67C���-}�2�^��=�ϥ��ǟ�!�Ӥb�����^S���`��3w���QSo9��/��%�餑�H�a�vC7{�4�<n{����p;zˡ2�VE$G+�Y�c9�C',a\��3N�]�G�Y^����˵q�$-<�B`���ӪM"��I�� �P=3�s*<~�G��K#C��b�Ss���y�U ܠpB��	��H���$(�`P�,c.	�o���Q��R���[��V�x�<��V��K�p(E�dN�����[rD-�n�"�.Ipn��;v��=[�函/.Г{��\R���6��~���	m�_>#�D���TU�Pm}��d�[o�_���y��#ݥ}���D�P��R���y�M�S�(lJ�M;�QI^;�����iٵ��ȋ.�ޤRMB�|-�����2�#���o��8�AE���̲;h&j��.V`JH�w�k�HH��M�����ǌ˽?�n;F�[�KW��z�F�!H���l�s{������eW5��q}b��Jy�)��?,�>�S,M<3x��><��[����C\�FĀϾG����ER�벅���v��M�[�������7^1���8&�*�X�k(Vmh�:"d5�|���'��M��MI.{���~�Z�VW�������[���L f�Z���#e��mt�).-�j�'HK
���b#�׸��m�Zc��ٯ�j&�� �>y�0N ��7�Z|�۴�Yに��ǟ�l�fڃ9�29��<��/��vqu:y�"��g��	��%�q+�����[	c���$L�?�'y�ŅE�x��/�;�(!j�����������d6s�����Css3��^A.���5�e�D\0=7?'���nys�YvS����vj�n=����Y�L���f��ٓo9�gH�vg�t��庚}Ujҡ�\W�cq"����	��z�mx�'?�]{�-�����شi�0da~��OK�(N.�D�t�tKb�����/�sh�~�]�������#`����O�����W��탃صg���/38�)6D�cɼ��Ɔ�����e��!{'����h�b�Zi'j��V�׼zS�I�h�v��HZ��q�F���݋@0�Q��O<�<��aff�$�<�s��p��bO6n"`�c\�pA
*z�3�|I�%����kG~�_��151�����\�����{�tU���)��-�wnUоG��ߦ*+�!W��V�����*�.��~u��M'��:*T�D�s"����a���A��q;!����/����e
\oo7w���{
.�OP�����N����h��P]�K�1�<���_��#>��{�`�*`�%�H��dW(���KGȦ�p���%G��|P{#�2E6���C�X/�`=n��c�`����#-��/`��ݢӃA��W�������6ҩ�ģ�WWP��<����-;��م��8�Ŋ0���߉�M[p��1:�9\�xQl���8H�8
�f�����ܡ%�@�e�#u)W�yWՊ�0�e���|K���Vl����#G���LߢTyx��w��|êM�F��[���;v\T�8.ӑ���ğ~^��*���3�-����x��^5�L�o�&x�W�2��vƩ�Ge��}�%��,��%��,ߢ��/!�L���U.��������?/O�{�����Ab%�����rU�W*����v=���z��ZB�@ ��b_0`�����B�B|,m�t�n{�n�B���w�įWuK�'��+\��z��]ʁUb�C#f�sMmmr����e�0%�V�������ͥ��ܢ��6-z���x��7�ܐL.���=�-�.d@!��U ǷXwq<�$��5h�r{�:�9q��U�[����u��6T��r�[�X/��Fu9<"�P�DEr�iqguIT��U]�
�gqaY��R&T���(+�t�nd�{���#���ܜ�'����|�N,�-���^��lXc�V�i�
)Nc77��!��P�5��K�a}S._B��L��1���	]:xy��rUrq�q	���I$!\��m<W��qry���p�s~yT�N�y����U�P��zm	��+Shmn�kg��������{�����kx������*�c�����O.:Sm����������3�[�r������u�\c�:C��u�!�غΐkl]g�5��3�[��Lk��-2z    IEND�B`�PK
     ˡ�ZI�)�V�  V�  /   images/f2dbd413-946a-4dd4-beb8-9b389826ae17.png�PNG

   IHDR  A  �   e~b)   	pHYs  �  ��+  �IDATx���|�u������+{��{OfED@"��"4�k��8��
(hQ�p�P��DV�N��Mw����;99�<���'T��^Q(]I�����Ir�)����-B��#��ea͇�~?꿅�X��8HJ���������Y����{a�X�h�W��������m����pu�����0��_����H_d�k���
�"1��)��`���S�L~�lt�#w�qGS*�`���Դx">Q�,�2@r��VBSA�V �z{gn\���w�LE�H$@Q$��<ᑣF-�:q����喦�}�{0X��I�x��m�6���H��@��Of�]@�a
#������W����{�~MQT���"dY�d2ix}�CS�N}�xt���o�!�̆��í�7��lY$MA���?0�	Bh��B(�'^�,}v鷻:;��B�����4E).,�1nҸ���ޫ��P`�<ܓ�ǥY.���i"���+���d�����0�а�������`�8m�l�4��8N;n���N�u��QgϞ�� o:ra:�e3��6`iSw�4�� L@�a
#[�<��O-�z~��4T�T �4CZC`�����3�-=y�7�tSb��7y�|zS���8a*\v�K%��X!4�a�aɚ ��㏏_��?G�W���� �b1M���O^>fʤ'�Ν�����j��f��Y/uq4�����MBh��BÎu��?�ѥ�/}�.C#f���TU�<��'L~jڄ�ms������PY�P��#9��F�pDKHiS�-s��-�B�FV�x���;�kݺ��)�9��LCӵ������=�O�UU	�Z�X�m��C�lNsS<aҤ�{������ !�F>��������ظ~��V �NP��D�����g\p��C"�,t08:z�eN�J���^C�r�:��� !�F>R�m�j�!I2�0BH$��ܼ�_N�5�T �a�H�p�\g��X�4#���������B�BAh�6A�x�{�Z��'	�!��(������e=p���
 ���ᦳ�;����-�g��ϸ��#�Bh F�j�,��k�4�"�H�64��+).�����yk޼yC*��<�{�֫�I=�a@2,DHc����M@!�wAhH{���ijn������n�ߎ�h�4q�O.3r՜y�db���(�����rUR�"�+�xG' ��;� 4$UWW۷m�tͧ��5E�>��6�	�j���Ə�{��ߞ3���.^,���s����|?$m���'BIQ5 ��Ah�y��g�>Z{���-Y���>D�	�iFJG�>w���?����Hb�r���� @�^����W�#�]�B�`�!��q��9�o��$Y,�֩�	FV~^����|�M1��a]��3��no�:#�S�N� �fֽ���3�:Q0�А��[o���z��������~��G��jJJ26uƌe3'���s���`�+έ�.n�?��Ѯ �� ACN����M�w!�C�#	�2�W���-[~d���� �H�H��8~��������j����.��/?�Ѥ	^ܜ62W�!����BC���;�ڳc�=��pG$	0IB/.)^>e洇����F�;�*)x ��'�܌)��Ԡ0������g!t�`�Am�ʕ��V\�ުU�<��2�
LѵhQqɲ3f�Yu��7w�.���@�K_?+�ǥq�⪞�j !����B���E�������;j����k�P$��'ƌ���s�x��y���(����do��w��0U����
�/��B�υ���C�l޴�>��U���F4���s���3^;e�o���o7�"���]{/csL�s,D���z��z�; !�п�����zÚ53�~��?8l�oXf�F�����ig����_�~�5��P��U��fZھ�٘���~�j��r�.�7O�B�FT� ڶy�Y�~��/tU+s���d2	�}�����Μ�;+�`��~�[پ����A� 	��i鞧�WݷB�[AhP���'���_�# ��dg�I�,0I�9z�Cg�9u�����>��[a��&C����,[2��q	��f���1��!�������O�}�����ǰYN��dY����94v츟�{酯UTT(7�v��;F�}��,�7�4M��L3���̤;�w�B�x�B�Bs}��͛7����u�	��mm��Y�ٿ�z��[���G�5���f�Ev�����ݼ�7}쨭�B��B���+W:��l��mm�m ��x"�s��SΜ�ڼa6	8��;��O\`���*DHC%��̻֗���vH!t�a�Ӛ5�_O>yݡ��y^�W(��3[��#$������u�]w%a��ӟ2l���AAD�A�9w:ˊ�!��B_F:mY�_x���������@SccB3�e�]|���-�L�$޽�Y���f]�A������d­��M!B�x�B��ûw�;Tw�^���gB�?���7y��?��g?k���
��]/� *{���F)R�Y��p�zJsWB�/#���w?�������&5M3���6��8�'������Oߖm�����"4�� C�0Ź��;�V@!��a��N���
�d͝����2�BGsswnA��G�~�n8���sZ���,��S ɐpopeV�]q�!��4� tZ����l�eM�ssrrN���Esx��f_t�Zb�N����,>�<�Aف�Er��*��K��W���B�`�ӆ5�w���No8�p����fffBCs���6�3_���[�n�A�o5��������
h��.��Q�>�Zӓ�W�!��1�B��?<�P��x<��yyD__H���2}ꒂ�#?�/�V����Lp&��:��@�f$!7����\�B�#���+/��?R�u���R�`�3n܇3�O��ˇ�����c-��7�l͂�R@������u�B�+�B�\UUy���u��-��ʶeee���C����5��3��k��k���H7��Ds���36�zh2ix�+D��!��� t�e�b��wV����zKJJ�����q]�\|�"�ǳ���^B{~�O09"�BDWAv��J
?ʝ3G�B_	F:��.]j[����j�<�d�h���zzz`�	��L��a�b��o�b�߿�gR@14(��O-���!��2� tJ�ۺu���o��˵�,�]�FFvֆi�'��⊊ cf�������� �Rq���V1;!��2� t�<ZU����o����r��󡡡���g�wޣ��v[�����՚_?�	n��R�A���E��q�d=�� B��#��>�����˿+K��I�ƃ�HB__���o}�y�F|H��o��G&S���>��)��KK���KGTV�!��q��N���j�v͚y���Y�_ȹlس�NK��\\:nܓs��I�0�s�R[�;]�6�<�� �bMM��p��x!��#� t�%�"�����]��rr�����2mƴ?]v�e�:�,�P(ߌD/q�,)�DH2���|�!��!��� tR�.^̼�uSe���xԈr�6�U��Ǔxf��������p���.�J����N �i��_R�u��� �:n0��Ic�
���{�͛��ty�L�6ﬕ�y���/{��s��Htu����@�v��&5�e[�����B�F:i�}�ټwW��^*u�Qe����1)Q7}�Y��|��8ԓBv���Fc�����C�I3�gg�=b�Eq@!t\a����v1����t��O��MCKG��N�,/,�l|�Egx�YsN��(K���)�BwA�س�(�۾�;>��]\\�m-&���ɓ�.���T/��ݭm3��&	
$��>�kiwT��!t`�Κ��[o�)����C�<^8�o�|d������?� w{�����C���x��w�f���ؽ���7!��	��N��~��n��k.SVT��͚Ak�͘�'C��4O�p��.��(݄a�I;����CB�D�B'�u���Zy�)����c��Xhllj+?�����V@�-�h��@����f+����(��B'F:��\�<s׎]���07>Y��z�I�>������bm���T��Y�D��xzG 7{ �:a0��	�e��Q�)%��D}}=����1�ƾ�
 ��{���9��P��RF�@�Г�q��ͪ��B�0A�y�Gl�V�8��p�y�^ػw����[Sr6`VU�o75������ �����B�
#�0�v��$���J˅�`H��:e�/UTU)�lrg�[��ϳ$Z���Œ��vB�
#�0G����Rk_�OkV�v�k�	#��;�����KE6��h�NP�Ź�B�#�s��:�i���s�
�`O/$�D���3�^1wnn�	�gCa�5��T�H��SK��w�4�	B�pA�[�h������q��ʋKa��M���|e�ygm�}���*�׮um��#X�@1�!+mb~��s��x�:	0��q�o��i��U�����,K{f]p�ss�̑�]��}D@3���<���,Yc+,�	!�N
� t\�e�Ҵ��x�;�cDnn.�yKm�u���/�x� �����s��΍JH�s"���ț���B'F:����un2��t�X�;�~I:�]Z��c�/���M~f� � �	=Jh7YX�B�4A�Y�x1��s��H�W�p�H�F���i���~����������-8�)
���U�	@!t�`��f��-3b��y�99���¡haY�Fg�3���?�������$-r� 
A�mB�TA�xq�"��/�p� �Bvn:x�:<q��5:�������,�c��>#Y��4B��
#���*)�tV`]�!C��1+';���DwG�聽�t���f��|
C��#}eՋ��|��W�<�SPP �--�򸛧�8�)���������nھ����x����i�S�@B�TA�+�]�o�K\����8=n8PH�4i�+7����7�q����l#����X��~%2��2D��#}e��m��&9�@ ��r��?a.����x�tb����@D�C��B�tA�+���~��ʫ�^U^6�fi���raa�J��p��B�fp&Yfc Hd�����@!t�a�c�r�J��?���g�l�0���H�8<v�إ������D�0����M��z$�!�N:� t�v~�aԑ��s��*�A�-��0��݀�)5͚Xw�4� �)F�+�B��B�d�E�3ךּ0?%^�b���8I�G����.��ϡ'����a)�����\�%�\� B��#���`iKS�UQ��<m�F +�)g����"5��4I�b�e�c8�!�N� tLv�n��4�1~����?n�ؿ̞=[�O�.^�y�}7�V���Ap�!�N	� ��=��C��_Zv����v;tvv%e���ǌ�S�����C�^������h��B�S#})�iw��\���Do�$U��"�L�2e�;#��� ڀ�S�&����$E�3�:E0�З���g�����szI�b�/�n�}^Q�j
�גj�wC	qE�0� � �B�F���z�-q��O�UUu���CӬ;A��E�O_r�m���T�D�b�}3�CQA!t�`�/,��?j��7��d���qܚ���?�N_P*|5�=�����7�B��B_X}��K���J��57$I����x���O��H � �4t4E���TuB�A�y����˖,��$I�ZO&L��vM�0�x�`���u�� Ơ��X��B�A�߲V�-���.oljgmK$���̿����)J� �@ C���"�j" �:%0�п���/���n�B�5�s� �2p�4v���s�̑}!�)j@1�f�@�$�$M�$�!�N	� �o���'��7�eY I��������Ϝr��R���T\! �544�$�^SSC��!t�a��7�p��|Ņ�,��������Ӧ=�E�}a�,["v��N�:(��I�j(������!��I����ԋtaKS�l�e9��@�4�E~MFY�N@_ʜ�篜۠�$X��X� 8E�u�	A!t�a��p}�����֊0ki�i���I@_Z�4�1�$��דJhn"��j�B'F�\5K��O�x�F��E�f@WT��ح�&���1��z��3�DR���Lz��>? �:�0���:��jnn�9�aPU5����喖�:&�
�фa���:@Tr�7��!��I��>Wݾ��&ح��X�����J�V_x�	@�DHO�P�B�
���S
FF��3B'F��^z�%�˯.��0em�g򂰶$/��	;vi���x[�X4U�t4�8g��t��>@!t�`����pV_o0�4��n����;ďnX� �e9��6��6N��J���O�hl,� �:�0��?�u��2I���>H��-�'L[��;o:vz��on����R"�$P�?����ӛ !��I����Gy��β��"�LإF춿����9a_є�)��ܳ��'��{đ	9B�Az�O��텳_{r �:)0�����ֲp8r���f���P^R���8�Է�4oL0��^Se\���暽�;y�'�ﾭB�pA�X'�_z����<?�H�iZ6L��I�G�t\�����잷���p�i"� BLe���U��4,Y�D�y �:�0��?x��?wD���S4pL�i���y��_�����ku�������^�ؾ�ٟ�<�H�P���%j�;��>�}@!tBa�����)���������/9~/���{�������n����x[@N���$sb�������C�w�m �B'F����j��?<q%I�w�R��������N@�]vi��;�6o�
��!V%�2!��I�=xG����̻"!�N� �wm�����X�A�4����|���Bt�y���Y����pr������t�V5�p˭�VW?ꭨ��B��B�����~{j"�Lw:��P��񭥓�킷�������߸����A�<�k'�#�CS��#���r�Y]�$�!�B�F����ֶ)I8h����+�(�����s�N��1cZ���IĢgN*<�u �A��)����ď��D�v��eS�l1�:�0�Ѐ�MMe���gQ$M���x����t�j�����痿\�q�qM9���?��
�ݴq�o�Ψ��ŕ��n��ǖ ��q�����;w�a�<� �q�
��u:᮹隃��{�7[֮���sm4�`M�V�.���;�ݍ?�����%Ջ��U�Du�:0��X�����M�$��$.��>��'�$c���(�>Ѱ���n�v�t�2
2(2-���eU��G�y���[q�<B}EAvo�Z��1M������c�n-I8�r��.�-��f�b�#�7���(F  �HH�����qW:���[���?����}�VQ�B�#����M$.�a����tx�1q"���������O_�����?OReN� 	���H���e�rmݞ'�?���[���tY ���0���%�=�~����W<.������(���Iw��gw���G�y��ӓ�viL���Ȧ�^l �G ���N�sCR��=�oN��'�����B�/#h�۹��$5�Lhl6�5F�.�B8�&@�ĥW����/o㖍1ɸag0�ԝ�fm�A�A:MEsQ��7zV�̪�����Ϟ�{�-A@!�`cK�,�?x���dY�[Ca�4�Q#G�̞=O1?���k۫���պm[����.s�L�EILp��L����;\�`W������̧�B�[A�X��/���w��i��=0�M���/� 蔫�����7=���P��Ɠ���`:m�&K+d��� p���V̛û��^{�O�J��x��B}.��a������>-�NN�!�m��!�� ���}�k̀N\0���������6�����&&��3����`��Ij@�*p'p�1�F�^>Ҳp�7���=a�ʴ���9sd@!�0��)ko�ֶ�dYq�a�.PR�:�J�V:�X�J�����O7���sIw(xEPNL���24(p�� �a	hY&<G9��ٯ�$��ڋ�m�>l��ᝮ����WvZ��!�F�p��ߟ/I�es:��@&�1[�2�p>�i�{�����n�^W�����֎�tSBQI�L +C�������MH�� ��F\�ܳyw����ؽ��t���G���!��@�a#h�N����'WJ�x��`�ۭUa�¢�#�q�i���BI=������#�J8��E^qоN� WR�t��<� OBO�m'ų�� �o��Yukko����{~�d����DM�4�Dx��0�4麞~����,�(�M����7M�27HRd��>��c?ljhY�}��!��nS�(�@%�W6@L$�IP�d9�OQ�����ȹ���9%��= ��u`�KYi��_tQBh���Z�׏��#eI��nEQL�a�
��p��A���vTWW?�v�Ν����N�Jey{P֠I�!�d� -!C�b��0�����Yp��=���޴qt׺7zǔ�h]���d��M�H�0�����.���q��d"�&C['�k��;]����wEРst�l}UUUmKG��H2�]�#'�5�2�ˑ �604�8�1�b4�(���jqrO}QGK��Z�{ö�~�T��^��jϸoL�dj��P�4̴���w������h��p$�8~�Z@�Z*��z����6:|�O^��s%M��� ���N�_5��T +�8�"ds�AĢq[�����#g�n���p}sG��#˖�)��.@�!#h���o��q]��#S�6�TU�"j3�
�_Xّ��~��������Y�H_��sc��ѫ��)�Ipt'�3dp��H�~N04^�ՙ-��M��C�)�Y�������`�F@�! #hY�z5���~Y$p4�(B,K��R�'�)G��ڭ����fSS�D�k��Ү�]���;�t�NzS!l�p�d(
�SxS�
�|��Φ��~YI���pnߞ#wr�M��J^����4[7%���
Bh��FZZZ��H�lUU	� �u^���O?�`	���hY�d�>������I�ŀ����A��^������8�J:���T��/m�N 4G%4�����[��ݲ}{�V�����hcCu�Ƃ��]��Bh0�FZ��D�i���	���i����v@C�cwݕL=�UUU���721�4͙��<�_���t;m�h��&�����qp:�	>�	9�D�dI�9X��G�3u�un�����d/�� �ֹ�B�9��a�����/�����Gc�pyi�ꠦ᪰a�곻5��ivUT��qe�x:	���ƥq �w�R~�ir^�t���� ��CG8B��(����Zz�:e�$$}T߾���Ŷܼ�cwn��tZ`W"`��lB�V0����}G�z&s4<ˁ���a@˸I��|����P��wo��z�Ϊ��{[;�k{�F�g�4��h�H�yPd��M����h���A!Â��Ap
�8�-:�l]����{zg�tm�.��/�g����;��G !�NA�Dsk��D"�c��Y�dPe2������xUU�4�.����h_!'S{Uu2�:F�&��uGK$�94��"����@G2DO�2���(�@�����{��z��ڛ?���M\F�����K��:�0�����]�_�Y��$I��4^�4ݟ�����/�BG�;d�n������޾$�����2J��	��g�01�ʹG�����L�.��΄
=�QpuE!�����+�C{	##&%2����pC˭�����o߾�����}�@���{�qcF��I�4�uw��t�LM�c�
�&FG"��#Gl �>�ѹC�՟�֥��p�������6j%�&Gecb����Ȫ�f2t��aFu�ޤBR�V�8y�9�6��+ϡRNA�?CK&����$��m�޽
M}ڵi��C�x������� !�N ��!�� �w�9&�>�7�&���󌴴F@�:E����>�_Y��+��|�m�N��U�~C/?b��@���Y�G^.���:a�š��n� i>/�Yi�V��H�r(<5�NR#���ߩ*j�+onem�ݬ��Vq�����#h��6Hlmi;_�$�5��<Ȳ��]�7����X��t*]೫5G�h�)=YBѼ�4t�G1mv99*��M��F�Ǡ�.�eB烲Dַ4 �r�iN�����̢�`\�� )�$�4CS��?����|��{b�YCz<{�9�0�����Td+@'�#��F�W�e�?���i��1�@"�5n�@�3S��g�j���o�|��d�u��j+hYn�,v��4V��8�$&���P{7i��B��nA��	Z	0�6�4�$�����y��O(}�}��{��g�$�;xdAUHp9$��sW�t�}��uNg��ٳ5@�#h�;x����$�"h`(�����l(/)i�N�7��gk½u�]}������&�ljӜ�����,/DP7�nE6����y����!H`L�&%�@�E�jay�NȺF���ӣFTY�Ե�°QS��+���e�!F(^�cD���C$�7�$ёu`G�!4|aao�����+��D"�5�����<^߇���À�I�b�
k�j ����766>�S-��vF9Kc)��I�F�HQIs6ݠxI&����
N�$�I g�x��P��u��iJdh�ER���I�*k�v��A�N���F*�̸nh�a�	Z�(v����`â˱���'���%КN�Z�d�1J���T:g��!#hk��)���(S7�:0��y3	��)�U����S����߆��Y�%w޹�J�&=� ��7�|'Cx>�'��`ڜ�r��(�&����Q�
��1HC�RI�0#)�S��
"k88� >u�IXRE���M�H=o�Bɐ�.+`����\�5�.	ȄD���0q��<"��4[��W�t��$�i�dCWD�=o��A	#h�J�ؐ-��#�p��*�!:�$I�0����E���ib��[wW�����С>{����e'9R`�Α��M�ϧJI�I�#�t�4�$I"�R�2 �W!Ӯ���ԁ�t�R�À��H�H�T�X�@P0p��%�J=A l*�l`='B*rD��D���rPɕz�Αv1e�f��I��*uك�?�]�r
݌�Ѡ۸��&�̪�,��F�5�����w�9#�ۭ��I�IE6<^�'��8�NKG�PF�^��z���ܼw/a}`tO����(�\�!�m�az9�)��8�f�&�9��괛6'ijv�0y�4��t���2�)j �R=d%0��&� ]Q�0�(|$E�ɓ����1(�X�@RWͨ��2a��*����ϪæC�N�<k)�P�rB\�p���Dm�NACTO0����3AUU�
�"(���G��$���Z��;I���X������!	�F S����J}���-�b	��b$G�,EӦYL��)��5��� 	-D�ui��8���4�,�%��X���ͦ�J��R� i�E�4A�4�$��
f+T��Rg�$Ê���^����?.��a��"�a"�N-��!�� ����(�HdY�6��o�����-? G�*YCm�G����ϧ!
.NS�XS��HrkB	C@�Q,I|�A80�:(֚[D�.��Lŏ��
&B�RqD�q�
#��$R�DMYw�Hpr<���GQ���	�wu_�KA�e�؍���~�[�������I�4Y$vvwOV�����t]7A|�ܹq@hx2�~�i�Q�ѫ�ꫯ�8#�A˴L�D�0s��ZN��t�6�x�ͥ#�1IÒ��� 	N7AV	^U�ME�zU�X��$��КkaIS��c2L�"I�LL�����t[��o~gM�Ȳ��KsvDX�����x�B'F���������J$4�0����9�!�wG���m�ik2�G;�ϟ�Zo�ed�&UH�F�Zz�ћ���E��5M��5�6���&a�CHE#jiSM�5�T1��z[.n ���"ȁ��8���&%f���	]�\�z��a*�_s���u��xaS��7�[�N ��!HO깡Pd�,�����a8��-cƍj �пu�Q��kk�"���j�eY�$<���H{R���4r�(ayb�-xx��8LҞ
!ZTt��TɩJ%�8u	`��H����a)�gB)����=ׄd���M�o�X��v�9�8��#hjnk�i�� H�ж�){�Ҋ{ !t,�+V(�G��?+�R�D��3h��3j"A��U(�s��i�:j��^4�!� ���XYV'��r �	kn�dy�_�k�ʔ�𡛶�߼m�/^��
>��qB5B�F����T��*AQ�@)�O����y"�:���1�������Z�ϟ��_1V�Tc
M������$����� M�-��[%��B*�4�+I�'U�cX��0�?'r�㬾��M9��myj��9��Q���j0�������?�1/�H�A֩�d��n�難�P !t�V�_UUu��%�2b�s�3&1�!ș�I���>���%T�epj�����*A��[X	Ag/��k�.��_����r���˲*+qcF��F��{���i��h��͚�iF�hkɨR�`��)rt�~к����l�к��;\�=��I���M�� �Hi��$NQH>�l����>�t_<�T��p�����l����;k��3�З�4��mj
�I)K�}�e�4�.���B�\EE�5l�<zu��#��s�z{'G��3;%i�������d^a �X�B1�	~� ���nA%~q�Ɲ����O4<���B���0������9!9��@ǁ$I�ru.���.@�^��%j���K���oߑ�`Wǔ^Y�ç��m���.?M�fe@�_���dF�D���T����<�[��tn������w B��B�c�|��\�eG*|>F��,�]q%B������UWWh�F_�ߵ�\��;e�1Y.�h1+বu���A,�!���l�M6����{�D��[Q����}�п�4�$�I������,:x�xÈ���������ESז�/7[#��
ň�ѯ+gFhyZ���	|	�x%�v�PB�;����hk�O��W��ͽc�ρ4�Dzz2$)9�"I�:.ð�d��?{�g��WBh�9:\�3���n�W�7��h��U�)9nN�����8L�!�"g%���D�[k{��k/^:��R��?�"�CS�������p!�x�Z�Q�	Dh�;C��Ǖ\�Sg[۬�`��~7un��q�h�:#����f?��&Zz�E�9�
���K��6j$>�� � #h�X�b����P(�v���2L���p��Аq4�����Xx���=m���4��L�7('��K��� �p'�ޮ����#����yw�F�3ACD]]�
�ц�q,���%��ǌ� �А�؃����EU=m��HR�L#z�� ��:$��6(�J���L0^�۟L�����RQ��9��!"
��nN�4�8��-�4t�����!4����=��yjˮﴵ�Խ�+����DY�7!ڟ ���K���ғ��&#Y3�-Y�ˑ��5B�F��y�HI2�(4Ms�.E�CӇ�m�8 ����G�^�h�Ozzjߨoj���s\�_MFXV�@�b�K����9*ų�/^��Y���B�F�K&��&Z�Y�$�$�4���\B�s���u<�hc˞C[�~��(�J�IH=�R4�u�@J�^ ��?l|�şMo�ߌ��p�4TWWS����S��(A��YS��^�� ������jK�\X�n���m��3��ϋ�>�%2�
<8e�"�<�h��u�w��K�c� B�F��}�v��*��,���`��z��BhX::D�塇}�e߮;4��HW.�I�A˃-�8Ӝ����������(���@h������HW<v����D�3���B��=�,h}lɒ�Z7oh ��APVJ�2XG(N�P��1G%W�޲�����U�а�4�B�������?A��*�f�rB���y�B�����m�����6���% "�_��H�w���#��/�ݥ�p�4���eS���6�f>�$�0t�gwϮ���@���X�Y����̾�}w�q�=���>�"a�˺�c��� �ؕ��w�a #h��@���ʧ��a@V�iw7B�UD����iS޸�����5iy��f{(	f"
^ޞ�Qw��]��{�� 4�ar���.� ��8e�l�D�%=��7 B�/ֱ�i�����o�֝��g�F��U�G ��߶��O���toZ�����4��A�����x�p�6k�DkNP����B蟰UN9�hѓ�ظ�7b@<�!M��6��{U{��~x�1@h���B��_���uh������۟�mWx �>�B555;���/{7;xÜ�@K*��s(���Үm���!#hK�&G̙sQ���kL�H$f�=�B����juu��������3N����;B�0�<�@���{;~�hk�}z �!#h[�bI�F���:A֝����0M�; !�����
}��şj��EQ*�cS7|F[�L�2S�����?>_��� �!#h����h�)��I�:/��tA��6�]�z@�/���R}��^9�f�8��i*�@����4��:]]�K�>�1w.Ȍ���A�����H�4��,�' �N�7!�%\yÕ���t>йeG�;�nO0
��
���ރ��R��	B0��xo�7�P��:�l6H&���z$�'�n��/Ś(�z�ꗏ>Ը}瘜4����
m.�Ijnoݾ�ͪ�k�*<�A�XL��uMs�a���X,f���X�G�:#Μ�v}s��Q��%ҟB�^�����3�NM}�@h���4�(Uc	K�q;!�k&A���ݸ<!tLfϞ{k��g���jJf�oFoc;A�� �Ew��}��.^\�g���#hc	�<���I@Nz|Z�V3I=�`�]�:fI�ܗ7����u#��+�F���q��k�#'�BCF� UUU��ߺ#��t�(��A7͠ɾ~�#!t̬�V�x�7Z��ף1�2�a�� ���'|v�����n
0�)Y�]�af��)�`	��'mG������J@�cu���v=��?ǿ�i>�)��km��>��ԧ�B�F� ��ї�
�LI���r���MMJJ����ޣ�<B�+��������w͉�wY @��{&��F0���xԫ(���ip��@�$��'����:�l[T�;^�ťi�� .o�b����ӟ B�F� ��R�f�A ��v�F��A��� ��q0p��/^��ٳ��g'�{	��KL��)�uF�F� TUUEo�ݙk/�
4m��������!���4WG���L��3uX�4 �B#���ԳxD�0����L�in/е��ޛ@Yr^e���c{{fVf֪�ʒ-�+��ŀ-7�=��0���3� �Ŝa��Lq8>����>-z�Y�L�0�xa���m��Y���$�j��=�{̽���x�^�̬�l�,ŕ^E��?"��#^�����&N�R�V����Z��b�̔�}J)������}���'�|���ޱ��lGP�����B	�J��R��=(���u�u��t;��%����UA��O?�t ��RJ)_'!�����z>�����t6�b�qV��r�R���A�I_�$���,E ����>~�x
��RJ)_Gi��q͖χ�uc��.��cPJ){\J�%�3i��e�6r+��$M���2�RJ)�|������?T�ӑ+!IdI$�~��Ƚ�:e��R��� h�	����Z	�Htl�EQ65�(#�J)�����v�]�����R˂D� 2)�0��33�CJTʞ��1����1��iZ���'h��'I�h�+AP)����Z��J���,G
H�� �?��R��� h��;��N��ｗ�@.~���1�
�ZS�˨�RJ����y>� �
H�� ۍjJ)eK	���,--�� ؟�)�|xf� H�;U���RJ)� a�Z��AT����r��+��=-%�c���d�Sz ِB��Ä\��Z�+��R�!"��vR,Ta�f��֞*]a��q)A����5Q��[+�AH���t=Ȥu�[n�@)��R�7@�����(L�2UͼZu��j@)��a)A���$�������O���;�3�RJ)����P(��_�-��u:� oJ)e�K	���T�j����I�����U�����R��](-ǃ����.��[.y	j.l�Yz�Mڏ�3G.����~����zJٓR��=&}�� �.Y�(Y"-�;�}	J)��Rv�Gy�	_
�%oɮ���`0���fE3vW�$��qVI��������_o�K�;���K� Da۩$��m<�п�፷������XlY_����(��=$%�c��gY���!�Ķ�v��RJ�UBV�7���孷�����y^6�M^���K�l4��^�$N����}_"X����߯�4md��'�d6��z%�$*A�T�$�&i�Yb�I�q��v+�������(�eiR�Ӹ$q-�6Y��V[gv�FV���5��7��=z����
��tz!��K��V�u�.]�}��7����G?����G~��R���1��!���	� ��n_J)����O�2��N��	��������tĺm�B�xwNۑm��D �8��0�x�������e�$b'���`�~�v�
)Dj��'ʱ���4��8u$��+�<S��xi�UP��oωm27I�
.+Y�V(!�̠�}r�c�t�I���}m��'p�L8i���=�y|�0bs����,"����Hd�}��X���6�Y�X0+J � �ì�1,��jMh���k�l��'�����u�ӏ<�ȏ�q�e�|){BJ��A�,S�^p�BS/�,�\/�RJم�?.��VqtmM.^���A��}����W�|�Gy��T���]���/ڑ�C�&m�=F�z4�<˲d��aI��Uq=����A�¶�,�� ��8�qY��
��J��������n�/V��jU-iو�HSDjҊ�\��RZ.�7K��a5��Vf!,��]jD��	� �O�����(�D�����80��	�P�T�;}p���E���2�F@Mʙ���*bU���on�Đ����V�Ѧ�3�A�m�+mHT+U\+`�ہ��̩@d8s`��A�^�^��k�g�x❟��G�	tJ)eH	����aڠ�&����_�1���Ȱ=.E��6�������]+E!7�m�|J'w���loT*�Z��۵p6/7�؎��J�V�
���/-��Wp�/+�G�[FIhe)j�8��`PEp�@%jۨ=q)	�L�z���~�����8OY�A��x������ܿ|˛[�^Ͽ�ė;�<'�z=��z��3Y�֬v�-�����jraaA�{�����ؕZ��%�o��O\�
���j�[V/e`Kٖl��'/-�J�ת��8ek�1�����ߘ
>P�`�]�����Ȍ��C�2э����M)����4�!�CÜ�~��b�L-c����~�x�	:O�2�?x2>���+���8
�Pl`�8a�mQ����Bm����]<��S/�E��!�q@V*x~�χ�hтh0 ĎP�ס�L=����%*e�H	�����]�ˇ � C��cۯ�|Ǐ�?z��+����ߟv:�lii)+�1 ���BU�/�6�O=�h	*X�y��w:�S�C������I�̊����@А��@��I���?a��;T�c�ͧ��&����*��d0j�0�8�߸���4�m4b<W�����iL.��\!.�?Ҥ��ؙ��$��(u�$���%�4v@z2��0����'���Fm�	Gԓ �#ba��J�r\��t6�RM���Ɋ%���ih//��Z*�*L�$�LOA� 0<��&��q�d�0M��U�N1��g�>T�k�ئC�6�R��n@���։4����"A��s=�mt�o�q���C�0���2X��\J��%������gN�v�<ؗ���"�jD1����Q`�"��_��r�	�$�x�#��� �,(
�~�n%D��Ȩ��g؇4&�A�7��T��F��l����bT�����U����R�ŏ�:>e@�9��h}�P�>�9�-^*�O����%��K(��lĸ>�>�x]�O�f�ނ�~<GZ񠏀��{��X'�Z���1�jT<kmq��>���;����J)e�K	����B%���7��.@zyV��JN�8Q}����������AT�4W�*�ZX�xz��3S_�b�bʯ�Z���U�d&,�Q��0,T��-�"@c�2�):&NR������� ���k����m�� P�TSF�Ҕ��rnHe��?r#�&��z�� }%�}b�#�Vh���q#j��licVz	�LɆn�B� �M
ʬ'�E�K�oj"�V�0��@�V��`�"h9XoBxq��6�ml����nn�	��5p"TҨP� ;D���y�VJ<��`'�#�p��J�55� (��u:� `����Y�g}}�֪�\U��)�����
8�Okj?+��r��V�<��3�� ��  ����-� "`�E$�jӅ>�߫��[���x�3�cC$���[��wG�G cj�3�g�}%�)��Y}�5�K�Jq���$1��~�to����'9`!`a@���+У�E[��В9=�X���3.4��-|�<�.���k�U�u� R�7�_o��6X�i>��G���/!���1=]��M�5cpH��v$4E*���G�m�^x���PJ)�\J�Ǆ"�2e7�AP���4J=xɧ?����>�_�t���~���^��>j�`���=�]w����i8}���P�6�S��ȷ�<48�QR*o�Ϙ/��e��(��$0ԂC���!^7��^*����M��0����.D8'�J��
��xnV��"���3�T�6�/Be��}>t�(聃��~ M���F�OM�K`�;�F]�cl$�\���I9��*p��l�pHQ�x�>+xo�,7d�±IL5|+���F��`��g�6��nTCޗ�+\1�3]���:7*����E��q\�����0ˀ�o�݇A�Rw.���>4�M��}i�5(A�"���r7	�������R(���t/R@=\z!�g�2.m���t]t�i]) i����������&��35|V�ޮ���a`F����(+Yf��>W�n<xn��F�af?�t�~��jNC����$؂�ed���jF�Gj=��O����x�/
�L,���!%�cB�|1f�"�Y�V�v��Ux��#��D�3=���<����0pTT��I؝�
�A�~��qV����8�Pq�U(�!x)�S�2q
3�L�A��B�F&I�W�=R�V��cs���r��"�rw�Z�D�@C���V��*��5��� R+�I@���1��֓�T�ѵ�t���8&TQ��:@,	*n/����8z�:��j!�@�V���8nA�����(�L��,���;�R�L�i\��w<�`�1a��m����{�[<�Т��a�bh������Y9�N�hh����W+k��^��zn����x�ᇠq���S��W�|�����lн�дGv9�Y������זc)��[��'�P���l��7r��]��˱�y&�D�h��]�:?v=���Bn�g/��h5����YN6,�&4+5�x�o��s��?kQ =g�� 5���ul��i����?G@����~�����L�Xʮ��1!6���[RZ���
��9q�����7'|��	��^"��;8c�à�_���LåK�Pu3���)s7T�ĒB+$Rt��Qt�}1������:ӊۈ��A�
�,�<5�#ȱx�o�
ەX�%
D��t``_���t���c��$���2�`#[c>N�A	����d���g���׋�B`#�{��	��6TP��[��4hLcu�z�%ϐ\/6sN�|���x,T�d����r,���m@��}S@�֬�А�(�Re�����Z"��8�򏈗"4������O�Q��
*�,�����tk`O#��qX��\���u��.XY_��N� �rZ�
T�]>b���psa��ߖ�{��ϫЕ���l���~��\/����q%[��٬Wk��,j�]�%m�R���[�~>���X&D'�q���#��L7�0Um�K��H���
�Io�,�z;��c�0�9�,  J}\�Y=�*0�����;�A��j)A��DZ]�2ϊ��Y������'�|��}�W/]�t�`�.�D�6�hB��l��4,/^�ӧ���_�ςWVV��h��ƫ�!�ȍa1@ɒ4��sځlh�a@�*%b����@H�˸ �uAQ2g�Ef騝4� +���D�]��De/8&��� 2"�st,�($�� Wy� �B�a���v��H�2�sq���p	�Xѓ��N����k0Uk�ט�ԏ����S3��o�v80=�n1+̘|k���[:���T�TT��(���]|� �@\���K��W[�V�>�]��_C�An@�� |e�DvIe�"#���h�$S�'`D��qj��%�̥�
�I�DY��1i P�p��\���n�ѹC����:DOx�+���RY��b��I$���nS~�@�V!3~�B�ϔN�!���8��54��ϡ����v���5�Wc����o�f �(�rǰ�@��n��'�)�8������V���@� ���x��8��+�_�ۣ���ٳ5(��].%�cR�Ȟe[>�И�J_^^���*�����{������[h�YE��Z��������W��_ZZ�:*R �@qh�b|�����1����,aA)sR&�=ak�d:xY+t����@R���x[�Ak��O`YAeiJ�r��eR���+C��%Y��-BV�4Np�^S.���*l����u���.O�����j,�l�%��!������_���]{=�զ��ϗK ��(A���)`�4 1���ܒ�±��R�t]�w���+%�VA@B.��V�e��"`�x��;�O�fR��Y
��+PGX���D*�̳��X��O�ؔ�Q�7`�K/"SC\�ިW�;��/r��z�oQ O�\@V�&X��,�->��C`����QKd\ G|�1�n���9�g�Ѱbq��O�*�qL\_�0�=P�����o���C��z��$`+Y�9S6���[P��7�^�C)��r)A��q"ǱC�(u#��d�Ƈ�*
��ң_�W���[.^� v& ���լ�C��g���I����Cs�D7?���"Y?���(�-���w�a��B �
$*\�2hb-pԓ��6��sÁ`<��
%.�h�P$��86G��"�9ǈ�S��c�69��z���g��!wE:�ՊB�I����2
��ꨨs��ڑ����0��4^�\Kd	!���9"x��#Gaz�Š��G�*=�2	-�u����+�E.��g¤l/#��RC�I|s�� x��[���;�TVؗ(��V�k��R���9K��5��x�u��3Y<K�bJ�D�c��h�qL.:MB'Ax�ƙ܄8�Ԗ�"cX�Xe��G\)�?@���k!��dn��)_��v�	'Aq�Uhz�� �[�#��3�7�)�Ȑ?�=�8bBsl���%h886�H���xce*�⒣֨�f�-�Of�څ�\V���U��:�����~(SGLc��������z�N#"����˥A{Lp&?rI�e�ig�6����{�׹��t���zk�O����*@���@��/�fŅ�g��4j/+���o~3��۠�^�^��/�^p�]Z����,,�����<���*8�33Ӭ�ȂT�c�A�J���|Tjͫq^reqs��@�Hu�B���m��T���9�ړk�"�*���!Y�\�vg��v��
,��p�=�����*�.WbH�͕kAd�*`�$�Z`1ŵ=q�}���J(��r�(J
�#�뎓*돲t�� �ی|X�����y�(O������/��v���=���d(}m��ڵdk�� G7�~:.>C8fxI�BnhI�y�I9�]���Pq{�8[�ǥh}�P,|Q���=� �ltu�Ʋ��cv��g��?�ꪼBA�����k��,B�Fn��A��K�}\�!$�<Id��I�+E-��PJ)�\J���q_�4{�W��bDqt�\�6��.�U(kkֻ��4��!��P::C~���46����\����2�rطM�cHi�4��<Ԡ�I`}e��μ�r���*0-\���	7��f���!�?=�C�!�G�Ew����\9�Z�F3�%Is��hx3�*2m!/�L�9㤐�Ȧ"`R�&e�`˕�n�:Q�1��HѲ`@Ȅ�9ya)��+�n5�X�� �8�I���#n����s�]�:s�!7dm�����o���D��㧚sdr�v�f�鱈�o���9��"Rt ���V6K���c�7��vx��YE�#��8���8�xf�老���A{L��������H�ė�l;�����9}ng�-��)~��/������*���c0?3sSX�|XY�C�9��K���5w�N��ǐ��@
��ߦN�d��^��8��:�"��1�4W�;�;LA���;yt�Xk  "e��D|F�x"&��Hd�T*���9�C�/Z�F ��"��WS<��W��m���M#ۯ KPQv�E�K���%��(��{��c�Q\
sL("�D"ī�xh�Pט����R�Ծ6��(�5�!��JG!8wɝ+��0�$G3�1n��6p��� ��A��19�"�Ie9|yq5��Rv�� h�	������8���&?�"߿�=W��,/M���n"~<59����f��@����y�=x�ŗ8���E_�ĥ!>΁���U������:t���@���m�\	�u�B0txz�k-��"�G������r�1r*[��Db�.�z�B�
Wx^��*Z�`���8� kX-|8F�2�@��"�d�}�`���cmw��eC��q����t�Wx̬hc��%�,�-YIF@���me>2�f�ɭ{�Z���5��7����d�c^P��1�HIΩ�>B�HD}�%�z��3p�����%�uh��F�RL�"�)(��].%�cr��A���.Q����3!�v�s\��]_��m���"�Z���[5���X�"�bh�.���g[07?	��&Q�A�r����@�:3�*���BR�5Yg�t�=���O21x�Z�٩}\*5��&��0�D6
p\r�⾀q)wsw�G1	_��V���8\8Vn)���&��N����@,9�N�'_o���L��n/����V�cR�֦�o��8��m����V�Rdc߇���L1��	4�%H�~f*R���F�w�D�]�V���i�H�*s6�֢�����	A"SEY�{F�$P<'�S4X���Rv�� h����|�y��(�#�!'����K+�(�
?)\Er��	���'����\X��P�4�tņ���ЬVt�u���)�-Yx�%M��8��nT�
g��������pM�,�`��2N`��,�S�iWZ.XԀ�ob��l�yg8o�d�<GP�yҸ��<W���%Gtg^N�X|���*6)�,�4l"[������K6(@%�+�+�eBN�p�dA���ܕmwu<�--^��bg�
1�{nΙ<[�v��7�7.�ǡ�B�]��rd�q��tb�Ps�8��)j��c��9��m�%���@��6VuVlH��� �᭷��n�C�}c��)2��m9�PJ)�\J���s��\�h��0
]׭�a	���X,�����o��!6��H�A�;���Ɗ�a!�!���t6V��AN`ey�!��T��aW��w:ENv��ρ� H��I�j҄��PE uzc|��2�]+�92g���B �L���O�3��D	�)'(c8t�L(������`�4��Cp!�Jv"�Ȳa�~LR�r;(g9گ�d�c0¶�z�\�@ְ/�"7� Lts}]0�]�܃�R��\8�6`�P�)��o��J�sE�R�%^%���,�ߒ~ V�ʑa4Pn�m]��w�ր���������&�6=�
�&�����A{L���s?��m��G45B]�A�A��>�k�U���fu0�K��UyeR�;�O9g�娩S�;G�v��S�k�몂���C����hH��nU`fzĔ��כ����,[%̣RT�4�U��
�]]Fѩ��v�&��އ��/s�V�n�������Z#v��Z�+�q�����[��ʒy��<�ܜ�t��G,;Yj��z_��þ�b�U#��^��
�t�����^�8�*>'�q.��ٗ~�P�����u�I)�y���r锌���ao<r-<|�E�:�~U��
�CJ)e�K	���LO7��_�ЩV���A��_P/-��R/�U$�N�A2��B��⦌�d���T�2���v\���r��h�����!��
��>���m�O`��UB�2K���"b�y 6�Ƣā��Yr�g+��& Bـ99���d0*��1Ҋܬ�8�J��� `T!�焜�1�]5�V�C�3ޭ���h;.�����b'�1~�I]+���^^�aw��rI�.7_��ϟ�m�Q3�c1l��u�M�6	�Mf�{6��Lѹ�rU�+V��j���*N,�������q
G���#,�]DIJ����J)e�J	����Z��~q�V�e����R��D�;h���x�%(�}�J����<�Hԫ=�<9�� *���D��n��֛�O}3�j-�64X�t�^��U=X�X�
����nw��i�{b��I�� ,&�8ӖC��<}�k�*��6n��2�)a"�igv+ZpF�7ֱ"�آ��c�\�
@��waξ��`i�*��r�b�ӋqkJ��B�=���k.ߖ�?X���l%���E:�$Gt�[Wsڌu�R���E�Kgٰ�,���:|T󎬱\�Y�$�2+�K)�^ʇt��|k_4/V��;R��^\�Ng����U&Y?�� �S��Ze7���+���Ĭ��s���r�	���+D*�Y�5��`W�*ޏ`~�*����s�|�W�$�
��LafS�(oñ���D����;�9U�/�,G�8%91d��M�,ۤgG]L������}�"!���G��%�jd�sWb6,n�s�a�t�k:w�Ị+7�1�5M��,^,j;.EʇO�����T�H%GNf�����z���9�*�;	��rR�DJ�I!��Ǐ����2B�R�7PJ�����mǲ�q]7h4v���,�q5����'N�w�uWW�t⎃ ��U�)|4�_��+k�]_Q�� >r-DI.\��֡�^:͠�]�z�p�Qx�ɧ��g�����7ӄ���oV��d��X�:� �#�q��.���oV}�"1
�H�5�d+�#`4�M�f ��������d R\�M��%��L\n��O�*��W
~&ɫ�.��Ѧc�Ā��}��,^cn�q�ʂg2F0<n4����Mr���@�`��f0=53��i���z,S��I�� pt��i�1%*e�J	�����=�	~�g��(��gff���u��ٶ][XX����Q���m�J]�RN�R�5��'��u�g ���~����F������!���I�5hθp�� D0;5Q�^AH�*U]�rB��i�L�T?,�ʓ�}0j1�L���$���.�N��U�\�6*I�� �#&��O�l����@l��X�:�&��1B�Խ���X�$�.���
A��x����Z�J�h2V�}���f]n�b�Q��;�@ہ��)X[��7�J�%��	��Z��1��j)�=*G�xb���s���ש��q<9�o=��i��X��D�x8�Eę��L����C��x�kt�Y\Z�q�@k�
�n���C��� N>�e8{�<>r�8��O�KU��[�����}O�>��N���u��@��)� �����%�4H��;̑	_�ņ4��;�p��.���SZn�~�lD���h[�L�M����*���*���y���9�Q{�4p�]�5�%�����yXbe�d�������n7����A��e�fDIBuq�<
R˾�H��1����8psԪ�����)eWK���Q��o[�'m�~7q`6�k�ǉ��g_�*R=W� r�$r,�� ��uqa�����5=�/�8
aie<σ�o8
/��2T�u�58s�:8K�.��XA�J�A ��YX�����*	�vyQ4��QB���q�ɭ��f�Hd���cۄ�.�}�5�>ۘlq��@�U�w�����y�##����b�i��Y��	�_���]v��F�4��$�<5',-XM.G�lk�7������g��nu�-��t�l�����Q�;�������{�i�ٕ���x).RF�d��e�K)�GJ�G���;�������3�F�Y�X�y��<s��[��cp�Hԏ,��J�r���:'?��|P��ʵ[���X]]��݄�I@�����@l"ʋS��U�r=ܶ�H}�/��#�Bs�4���)�����%2�@�іͥ(�F�M�f̊��V�M=�I�b�$�'5u����]2)��5U\R���L՛dͽ����cn��f+K� %�~K!�o4�@����o��b�.�0z%r���I�W��n���i<�9��#˫��f�l��~\s��s\�1Q���9BL+Vv�RJٵR��=,o~�>���Ǟ@t��d�GaE�z��������}�u) ߨ� GZ�x)�#e�����Zp��:�xõ��'�"����^ aþ�}0��=��=��5XXX�ť���L�B�<uۆ��RZE����R
��q��%)��X�G�i�Ř۠�<O'S.<K��Jg�Zq�x�����BY!h��+1�|M٭�Y{����!�X9��

��LcGi�{:ct���g�+6�F��5�X��B�MX�~��������$'�U��gG36���L�C[��-';Z���l��`I�t�[���ig���'���30���Q|V.���q�`F"NY�9m�TDw�[��\'qq�ͯ;3S-�uC�{��R�B������RJ��R��=,a�ei��J���Z�^!L�B�����W�~7���J�W��;d�*iL1��@���'_�d�L�Y�~A΍��G��V�������E����@���˕B�YCEB���TQ���
�8�:s�| �~u�N���7�!��a͊�a�[)����4p��!����]]l|�(dE��h���
�6�8d�Yl"e>W2h#`S���rK�9$^�H�5B�s 1Q���lQ��ז�%!'���U&%�@�;1�|0�� �4���d��)�fZ�g^�f�k�4��a���D��T��_Ct�$2�N�-'�r�?W���#(h�]:��>��9f�4�:Q �$�,X�$�CV ۑ�E� r�s%I�RV��Rv�� h����~�g��6~�^��Da�.ͮ�t��_������l���a(Q��z��×I����4kU���Moz|���@��2K��6o}���cG��Q2��t7��碄oI�����KYZ���ʀ�JM)5Ҝ�Z������?�=�:�r�5�&LV �|Ǆ�S�#�e,
ў��`a�"e���@rt\���V�� �tT�ZOQ<�T�L��L��8/�Q�(MN���6+E�^	�#!wr)#�p��1^tNlO���\��
�Te$1$�"�)
�`�(�ޔf�@�h�2�`;%��N�%�ɶ�M���I�0<�H�1�c,Nf�U�m��[�6s�&�����������2���I N?AN_�*$x� !�;�SJ)eK	�����M�<���}��]_�*.���%&}?���z����g��5�V|�Z�����,�:�����<�~ny��pۭo���U�&!  P�m�#�	 �Pq�N�ه��/��VI�!��f4�v��r��g�-n,�\=9*F��yY�0;�r�Y��c^9q�`nSF.%)�F ��,�y�������NW�/c�7l���U��pߺ�������R"�D����C��2c���WeA�x��d�;H2	>�K������W�8��M�_�䊬4�����ɻ&�����5��u��L�$���d�]�ى$<QƹDy?�թ�]�n7 c�y/���	�d�o��7rW~��8��#N���+� �D���:��Rʷ�����HX�D�!��	�4��PJ)�XJ���~�6�|�����?<??w`��EV��:�����#��Cج{XR��G�b��T悰� �*�����,-B;d��g|���8Tށ߅��1sb�W!��+��Mu��f�']T����%��j��F%`�s:r·`�N�T����RE��⥚gA`�l5de���D�j�ٜ�:E��5�R�jܩ)���P�yv�
MD�Z�^��'���jt"%Y�¯�7��P��\�l�I�|	���(w�C� 3-�4>��,D �ڜ'���A���Bem����ј%�"$�w�}�d!�1$��� Y��˖���,��XN.�U�l��v�#�
�d��h�>���a3�1�e�:(�8۹�
�' �qΕ�G�Kd�?YE����:���	���(P���a�^�u(��],%��BV�~������8;@� **�/�������>�;
{X� p,˒��Va�#E��X[�Ua�c��&CE/��C�g�UG},�� ��X�����h��:�I�G�Y�ExS3ybFe߷/���,�Q	�4Гe)Տ�81dY"+���D�W4ǅ84B� ʈ���A`��$��
�3Ӥi /��1_�Rw�_��=:�&�X�5$ϟB%�5��`��Dx��w���T��}��j��!�:T�\&x�A��ssj�	I���E�@��?��}��$e��e9�,�R�eI3D�M��+��l�6>[���:n1�ϕf�޶����Je{�YiK����yqi:t���JO���`���2��d�VSܠ4QدA)��b)A�U ��sυ����A8��f�Iu�p'���Ƨ���?~�)�|�����P�4�$U����Ϧ� �^u�C�0=U�8@��P��P�P�;.�$��T¨�۩
��X�+m�azj��/pr�5j�?�QT�M2�b>�qh�L�=S6�*Qe���)Ї4h����J�\!�=lCl)49;������ eF�bLVM��2̒*��tl���&�`'R�< x����'�3����K�l�8T�n���ǄR!�c��qL�ƅB$n�@��k��I���JJlN5�����q��D�"7�� ,X6E{:vY��4oNb�{�����ˣjk19��}3��u�&c���d�Y~�2��:���| 'S.1|6��\!���qYI��]-%�J�kj0����o9}�4=�v���O<��������{TP�i� &l���Ds�b|{-��O�ZŁ����Dq �S�>_�,LMx�[�/����k�e�f�Dv\	�]w�p�PA �"��$���ϙ�dbk
����J �,<�]��2j
��c�,�V�*P��� 9�����	ܰ��� �t[��=`�U�S �7��_Vk��+Y��ik���}h{���~��n0�T��<a�� cEL�Dw�q=���(0�\l\/��i��(w�2(YLt�	��%�Q��U$��3E6�I2�� K��]��7!�C�s�W8W�Gu8sY�%C�8J��=Yc����I�u9Kr������!+��د����e�1׳]�Z�e�y[��6slӄ�R�7��F����OG����wC�u)+RJ)�`)A�U"�V�b�95�<67�Ͻpa�gdk�αO��~������w�y�^-dI)�4����^@_�&�
��ۿ��5x����#�C.�c�nۭ���=��rZ�:����e��}��ߟ}��P��˛f�d	����H+���!�P�I�(d��e:����\�I&Qs>��r7��
�2|�兀��F$^[���C �����܏x_��$uȍ��#`�v.�"���MQX�7ǧkIu��>�N��E�*���V���)�G+pJ+`�:L�UddL��Y�0I�l3k��Q�cd��&�I��3r_؞�۸Y�ѡ���r��3(�*�f�Ly�f�H�"��d4��]l�~�O��wݯ�&Y�T�@U�;%Jdk'?g�ܼE��>���r�/ǎ�������3wE��RJ���]%B���{��>r���w�"��Z�
�Ż��p��8y��?`�'`��\Ҕ�I�V,hY��a���p���ْC�tΞ?o�����e�?p�-G�v�
���p�5𶷽���w���}�AO���+��܏�e�^s[��ori�فRM�͔����V������=W+�g��RK�9�b�/N��]%	�V���":�B"�tb/1زD��J�,V�*,���	����B&�
��Sԛ�y����r��F�����i��؂/��R��h��$�[��͊�H\�Iɋ14�-{K>m�����T�B��_[�o���#�\�"�z����!F���um�3߉8O���pjD (S�B�#�2-MFeٌRv�� �*��o���ӧ?�����[76:u��n۶���/��w}����;���u$�4��l��  ���ɇ��C���env�={��t3�n�!.�V; m,�~AQ��3���U=�x�"���U�N3~n�a�D�)+�T[
�lX�+.�ȑ�ʡA�0 IgL6n��d�� (��Xj�� �����(2a� lmm2�UsWP���η�B��\�q+΂,!�ЌKXȂ�tҮ�e,d��a7�vn�t{4�m:�f�U�v��#�Zɭ&���Mc��g���(�� ٪[c ���|	��r�t�h�gTi�9Ƣ�@>�-yģkw�|O�T�J��z���NJ���Tʮ�]Er��w����{�񟚛�cDJ�R��N��ʏ<��ß�f��=&��yb�$�n߇g�y?��Y8��9���&�N��^��V�l�"=z�]X�gO>��4P�d-����"��I�́���`G��� 	� 
���r�,XyF\1��"5�� ����x�������k�g��s&7��Lt\S?Mqh�^��,>� �Ǯj�'�t��T���h�����)��̅�I&�MDf56����*����O�r���2��$��%�tnY<v�[��\s�e��][��M%��N&��M�3�H/M��_x�n[�#c�ǨXS,�K���r��u6 �k�n�v�{]~^�rᖵ�J��R���Ln���'��xa�f����gp�_�������������/��R!.S�f�K�8v���PkLA���F�_\�'�z����4�v)d7���U��@�>��'avV����[���Ws�E.2�~ҳ_'��K
��qo���H/-����0AG��rt��7���,7�$bX��H�������eH��+^w�e&��Ь=��a�	`�h�1%�&ro���à  ��JX�A&�v� ��(�ȕ��-���8��r�'�Xz&,�e�]��!>�5#e=��f�r�Y���]�����[��֛�ϕ��#>k�S1'���t�j��9���JwX)�ZJt��]wݵ��������_|���������w1�������~�C�?�g|��xRR�~-��CuY�SN��
^�"1o��rDعs�М���KKP�ln�AS�O�$p����mw0�8��QX=���(����dI�]Y��P"�V�
�M
m'��7�ĂcJqX ^pBH�yspN�^�U��2�X�'�>S��v�d�;�bM�� �hL���b_���ti�oݓܘ49Y���f;�2ґ禰=�P�j�=�6 E���p���]h7L>=�ް�F��	��B��X92�C:y���Qj�Bt����Р�SQ��]͊-�+WX�1���Q:��T�.�]��o_��׿����S?Y�V���e�ի��_���}�//�8q�����B�AYRX�R3S�V�!��$p#�W�����s)i[�֡F}�:����8AS3Ӑ�v����~A���v�B���T88q0��E� ax)bs�΂�/��K���C�E�!5�8z�Ŗ0��\s�8�Δ�hD�R��L���[!Ya��`k��&{��1
�HLc�t�@V b�ʓ���h#�Z� 󢝓�\ɦ�A��#�b�9jl]#�yw0Emg���lV��=�kE��&���d#K�4�~{!���"?+6��-o�u���i�ru�>����
	��6D�f�YPKKP)�\Jt
�������;g^9sݡ�����		E����W��+������;��^v�8N=�e^aA%8Ro4`G���t9�� A���+�	�*���o��ZZS�����k�քv anf�fz�U�!��!;���v�����Db�-,ŚW,cyk��d-�"˴f�DB�*�\���2�J�Qmif�E��C��Գ�o�2�8S}����d-`s�f����{q[~���͌�¾�z_���,e�`qɡ�B-��/\��Q]�l���H��Z�u�ID�$P��ڦE)V�/F�`�mr�a�_���!��,�
��Џq���<�4R��Z�>�����\�R���Tjӵg��{����/>q �M���`0ah~����|�u?����n����#|��q2AehV�ף�f�xma�ߗ�V��V��0� |�gaz�>X�m�t%X��Ϝ���ph��6llt����+���ŕ5z>��8���6��Be͐���lf�BG��ù�S#��^ ���Qل�)�T�R֖���3n(�=_���I�Cy��)�ct�C"Q��9�\�ә>M1EkO~�����1��s�*�ILG�gl9�F�\:��b@��G��3њ#uʃ,���X�[ 9��ej�%��$�sN�|۔CiL��V���:OS��ג0�Lz�ID�Ϻ�20�K�ԙ�0�돤J�)�Y��U���u��4^J)�UJt��]wݕ|�ӟ���o��7����w�B��(�f��~��G�m�ۛ:q�?���6`�J��L%� 33M��D�*����]_���7{]��}�^-[��:������6`yc�����E%9�1N�vW_�V�c��6')������*Jim=�w��-fm2\fť��[,G-#b\S��a:¾�-�ϖ,9��nT'`b���m)����s<g�Kn�N���K�q.��M9��dv�{�.�
�~�	`��U&
��5�\[q��d�Iu��t�8F�N�Z��^Ŭ͓@P� ��L���R����H�Ë%��lzI��3 ������R�a*MS�*T��R�����R�?�� �*����=�����1˲�O���Ç����OUVV���)�Qr�駟��?
����~����r��;��u�}�Z��Y�f��h����rg�ǢYg��#O�������=����3�K������G�O��}�Y����5B&VSJ�z���G�HQ�g)5�F92'�4,�  ��_���,�m���l�OL���'���mڢ�u(�f@v�2Tȣ��v��}��#|oq��@�6ܘQ.�������i��!���B%��d�;m��)�<%�m��f���<0���R)$lYc�#��JU)� Z���s�)�t���7�R5�}U�9s��!�3���W��Rv�� �**�q�ĉ���|���=z��,--5��֨ԆH�x��N��G�����?��?����=+v�/�m���
脀"�a�j�y�˹��!�#|�Dmh4���g��F��Q`YŃN��k���٬s)� �7�t.���,{�a }��sT,�C�AMD��9ig����l�}����lX��2�;U\_�<&	b^�A:��Q7ʓ2.���L�yu��I����t]l�s��(� &ԧډ���C�l�;k����� w)&�re��F����� D�[�����9f����	�Hx!�O:%?�F=N�	�#d+���:�d	��
3.����/�\�����5hV-��.�\�.'&u�w�^�^-�S�kDJ�r���+��~�s�ncff�-K�v�]��[gΟ���>�go��w|�w�� pz ���j�Iᴳ$��8��c|��;�r�5��T""ƙ�����-�u{h*t��jHe������N�o;T4U0�A"πW��}�\����Xg�����m��L^`s��;-s��P^~"�@�`��!���6����RE7��g��"���}=dcXn��r�
y�g,qk3^@tD���2���vG�>�
�& Uq|Mm�qp2i9	����f	2�,}y��>��{�c��nu>��xV\�?>�T}ŉ3���ww�߁/�z.D]��
DA1N>BN~���)�R��+7�R�?�� �5$��k�v���o~�>555��3g�����lRvA�����_��_�˳�ξ���m���>��?����w����sIضs)����MV�$�oc��{�� P�(�bX[݀��76,�����,G��;=���V`���zp���Ckj
�8n�{�y�v���<���şX�%�g˜a9�tr�+�0b�9�9׸ fF�kw�xك�����CƉI
�"��)c�1ٯ�P�$�
�����U�u!Xk,t+�
m���V�����ё0z�I
�r��}c4k�l'9OF�\}�4�t��(�"!c����$�Վ��Ju���YG��`���V"�Q*.��4IZb���$�&.)����R:��ť�����ogP��8!	�9"�\��@t-<�pA)��b)A�kL����������O��xwûs}}�N	g��h0��3O=u��/���7����{���p��w�}�?��,��K��='Jb6���Jq�|�2�����d�����A�Z����H.�
��A8w����S��µ����)?D�&�u����".��*8�J�.XY@[t.�+qw����(�qw�vBm��$]/L���x��r��dZ1��l��'�J�̍�������XEj7+�+?u~oy|9E ðy�x��S -aƢ56̒@J^#n������:����ϝn�ր�In�ܒ$��qę��?��Dy���h|����2<~�\
z��$!�ES�n�%	q>2����M&���R�.��A�9�����_�����{=�}����Azy�K�,�+��O?������x��������?��{~�'��������>��)z����S�\��3U7aw��:m��yp��a���O>�nǶ���b�4?3���" ��F��c@n����0�9�'h̆�L�ȋ�꾊��;-�+ ����X�	
�����q��Y���X��d��V��srv�	�t�2����	ݔmѶ�n|[���Eb�ɴ%���=��H�q����е�c�����)������q�n7>����f,RE����i4��-b�p_�-K��6��� �y:O�-�s�_���8q��7Br�*��o�&�N��t�L:�*�R�.�����w��������'}�����ӿ����I5��t-�8��p����_��w>{�����������yl�5�,�������}�u���vvn�z	H�,��֛_��K��-�E܇�����2+��T�(�F�u8�Z<�*���`.*���g��Z6�*.p��g�1�A���̕c�%WwpHl�U��P\?�����}т��]:���&Rw�\s����5���Llg>�.+�����SF&���πQkS{^���#��/t��#WV�� �DL���*���X�F���[��Mc�mX�e�u��O>5@��� �m���>5t��`��lu}���o�d^O��-�j�A����������p�P�v�?��|h6j��4�x�П=p�4�R�.����~��M������ɓ��oO�p�'���F|Uګ��0=մ��޾/?��<��Sw���Ͽ���?y����P�.�S������w�����$�.fJ� "�Rh/��a�� *ຩ�&�p�:��@\��cǂ���!��\�T�ʑr�N-����K@@���Cщ|�����̀gM$�;s[L�^\�����9��-'㙉��He�v��2��Cј5i��#�-^o�V��,:Ɲ���ҽ�u�7�i|�82�A��DE���%y����1w�̄*2��2V��nS	DkK�VחN����ei@!o�>E�f��ʒy���c�ŜLR�o!#�C�	���[~Z��bE ���E�r��F�	�t,
�����}��k��!�J�_s��+�� ���[�A���s��s'N���ӏ<�O>�?\<��j�����eER����r��~��w:r�ѣ7���������{����F��;��yBhy֊}��"��p&pl|��ߍV���||�����`�u���������VP9U<� �s8
�9Be����|?|�S������ʜW��n!�&�cX�\.*���� 2�n�	�/
�o7��E�Z4X�HM�0�_�v�.e4�9wm���`�T�*ۼ� D�2� �✊�\���%�,Z�^�E��!F9Z��e�S�o#gT�e��B��2���&^��<t������Yu�n2s�|�8p)�fz�q�k�����YA��Bpz�z�e8�p��1*�t�D>%v�����^X��~7�X��������Rv�� ��\tA�G��ާ�<��Gx��_q<�[���:d�р}�-_�:��{����~������������{��ܛ��/Wm��=?��z�˚�F�/��L����^�T�����5�S�s|�9�Μ;A�/fTPۅ[n:
˂�f�N,E���\a>��E$�m(���U�W�������H�(`#�%����B����V��wƀRbE�Bߋ۷[�vfY/�(ee,-E���H��IY#�|��8���/��b[�۬�{0���>�C�ٸ��]������*7Yִ��|Pa d�������� ��\l5ʆ�r�$�d�Ѹ�Ȑc�L�M�D�4���}`�G�	��<�j�83u�]�\�%c�e&U��Ĝ_��8o�_� �>��a'�#ʺ�]�0�?�p,����߹�$t��ȃs+�pacV�IF��<�ڃ�hNMq!\d�]X^�j�����R�.���I��n*�����z�K���W^��/���f�5"&{05ݒ�8X�0>�Hq��_��y����_����N������^�v�ᶖ��'��j-Ep�$��jkE�P�Z2�o��q��v��/s����ZU�{�9~����|A�qf���w��Y�֑�`�d�`qد�@�H�+���@����C�[C@,��nMr5�6'$��Is<�\�b�A��0���B�{E�������_A���I��L�<q��X1�M���|�R�K�oUI|;P�2��
6����ȓ<���# E�t��Jb��ɂb�zj!�<��]��Ӝ�&kJ0P	3�O��j�����K�&��v����8Pd�!p��X�I�.9ECJ8�ʀ���[��I����c!4 �@�@���E:�3Y����9n""����F���"����8��J��؎��[����߅~��>�z�8YJ�0��;��;z��硔Rv�� ��-�g���/�8q�w�/\�ة�N���g���s��ܱ�ޘ�zrmq�ۿn��u�9R�vۯO��u'?��?��tiej��J�Z{擟<�����88{ڞ:��۳%(	��ɥAď^�����=��K�L�Z��?��a��E��;X�����ۯ�YY�����jW�cw�����8��	�HG1��^za���!&�?@��Bb�\�Tc����ff���ݧ}��uz�=�<�}�ڵ����~��j�޻�[o���Wk=k��C�.�|��3w����%�H����� t��I���&��̦f8ۡ�PJ}w�g�8�N��)��u�ge���=.���� ���Z-�������w��v��s=R�5b� Q��&d�CR�l#�G�����ۜW/����A�۞YU�=G�׬ ��R�g���������j/��--+N{q$��P��C8ڋ�n��=*y�e����K�8�E��y�k�zۓ�k��e/Oy�'ɼ��.^��Qql�T�Xy{́�|^o6�˿�*���T��Q��(�����V~�c	�:�K����_������r�	^���7m�]O����WmO���M�������fgc�n9c7Y�����x����~�O�� ?�A�/5��߼~��k�o��7�~����⯿��7�>q���ߺ�ޅ���ڏ]1o�z%����یBsww��۷o?�����K/��,/��A���w���~gp;non_x��{�����T��#?0/���qQ��̼��7.J���ݲ�J���U����]�?�۱ܯ�>�N��Fc��5���g�yF��k�Y��������3�~���]|����]/'�JäC��8�fxrb�P'+m퇾�.�z8'��7��7�_���n��^Am��N��������N��e1mP9<�r�@p48����^��9�eamu6x����ܜ�Ӟ��CG����<ʦ�Y�S�=jU���V~Ι���D6�ړq2��`��S;D$a`Q���!����u���^��Y��`�.�i�P�i�Y�δ��fg�սP����&���U��t5lz�P��WW3���~����R��0b��Z>ƹ�]�u��L�3�GIs�[���_�<hd7��L?�MW��F�5?��e�����܄���tavvv��ѡ�����/~��g���<��_!�Ҭ-�����O��;�7^yǫ/}�=�o�z����;���K_���$���o�hv6�����=a��	�A�>�?ܾ�{��왡�!��h^{���F3��ze�AI��2����g�7z2��mO'';�`S��߳�i4��2�*�?��z����S�+��K��/ҩ)�Q�&�]e����S����?�����5i �D m{h��]����.���~b�2��,0���WU��-l=�����������`�Iҟq�'h�5~;�VO��ӵ�{kT����@۞�:�Tˢn�MW1^�i�K��b�΅v������-��=8U���iި�J;��2[~Y�RՁ�of4�Q�s[H(��1Eq�R6�:��?9��d:���N���-��z~u�o]��4�+��)�L>Jiϡ����{��&Q��"y�;S�e�Ms�L�X��yM�Ѯ�:կO�EՏ�����1V�}��ZU���������5l&W~oN���,Ow���H��P��'7��=3����$Q�h?�����|m�]3k[f6:�s]����k=S�Y�������?�;ׯ�@���A�_���?~ W�$��u}��^y�k7��������x<��W�>������W^~Eg���``.lm���M��SO�CW���c��~C�Ǉ��@%m�8T�xc����`�΂�o���L��<8�+��NV@�,k�E܍�;�����dak}�?����������?����!���`�����܎��ɑ�T��uO&� dr��Մ�F��6+E��g��a����P���B��JO�jo�m��C[F�S���vGkJrۊ���<�ln�\��k|	�����k�G^���z~�gu;�-�a�^��K��r;1���n�PH#JX��zm]\R���vF��ik�7!�=�3t+�R�m������CT����y�(����x����ŋ���hXW����Z1]�oC~gt����qs��!:p�o��3Ӟy̩\
�9.�E#u���.����ʓ�!���<9wM����������pӣ���ڭvj��l���7OW#�����vvxկ��Й�N�Z>���H뵭6[��oN7hΓ]�A����7�ژ3�I���<}ca4,˹���/_�(ѽ���邈�b��o��S��y�倃$�=N�p����۟~�������h>�I<
A�?iz�v�"����O������n�|���޳�v�<1�L.�O.���#�TG�X�r��5��4�^y˙<����F�+��f�&3��ϓ��w��yj�NO>'�V��,�@��X[����H�ޕ�O���f���.x�S�u
����4���.�(�b.	e=�L�T�~i�3so:2�Ab�Bb�M�禐�ҋ�3��������{�2;M��^����BܶVdn4��m=��l-�Ւs�!�������1h#�=d��aSǢ��>��jn���	������봨��F��@e�J��Ah�۳C��Gvcq�������֢r��@��GZ0�n�jCUs�v��WO���VC�>�T�W?��y��&m��~��M��0�����=��zS��l�\��1�I��>fW���P�t�N��Ϧjf&$f}c��vx���gr�Z=/�.�������-��(������AAۻa�uo-�~]{��ve+��)�g
ޛ��@c�J�|�<�By��c�oɆ� X�$�7c{��yj�����9��~��
����8˚�&���ד:�*ۃ&ߧ�w��ڟջ�+�Z�j��,:I�?����a�a3�H ��M�&��\>/0��|�3�x:�4�Fo��?x�����x4ܙ���E�3���4Ml�n�~�'Q�a,[����웯��ni;v�n�Ӟ}?��)i��Fu�N*��an�<4��،�3���hh{�l�$a�׉Mo�7-��%4��J��Æ0i�s�����A�5�@�%k��<��b.�4"��l�ʫ���3��쬞<+m����"���\ۓ���f��:�S����J�S���0�6�Z���up����~.��3��٥�ֿТd-��߆8�ڟ\���z3� �����9�z��Y�ؐ��0�����p�'F���X�PW�3S�͹^//�!m�?�AJEC�����C�$;ģߛ�1�����z�Mo5��qe&M�Z��S�-��~�n��B�K33��6���l��Z�{�qO���
��֤�acY����T��p�Q^?4=@�}�^V�Z����mjg���5_��:�2gˏ�_gf�5����jW�^Pr���N�˯k(/API0-�^W�mP�5L�e*�$�ʙN��0}�AU�����;I,o	���O��o�x�'����+/���� |O5S㵼�fs�������O&�Y7	��,�z&(⪊|똎��0�FY/Y;���S����������_H��I��������DAeg�\�~��m�\4c	I��Kk9R�&��Cs|26s	*	7������fMB�,�Ϳ�~]扉�z��@���|���+l�R]�۩��p�m4�|t}�_�$m���K�y���B�=�z���ahև���EU/�g�?yn�VW��k-�U�<��i��=>:L�S�u+8Us�y�:G�'^���F_�f����x���:r=�q�c�'�9����������xIb棑]�;���
��X��hl�G�eˡ����egNɹkH�pr4�����'KC��ioV;��n�!Hi�M����q��5���t�4y�R�U�I��H{<�������rl���ci��nL��F{�r��6�ڡ�vej��4�<_��s!��_�G�ko�]�}��_�J_,_y�,a�w4D�Mn�\�I�v��	4���R�/�0ԗ.�=�����Q.?�C��$��<
�q�(���8<��d,�c��I&a)�`�Iziz�+�SnomM/_�6�rႼ��}� �#? ��2��qg2�tu_��͋����W>��}�c3�����_���:sD/�k���}�_�էt��(�C�7���=6��e#��f�[��AQ��d&�ff.]�bf�S.�E�w�����HC�7<1	N:4�:��٠�Ck���6fkr���?�0����&iȱ�i`(�0c�Wlo��$��Σv�1:�_ka�n�:��a�o
�m��__�ZD�6~:|�u-H�~�g[��,5�8���������Z"y|�H�(�u��L��b����M=�ȴ�����[�hM��)='�<5^ح���ʤ��_����H:I1�δ�=�|:�ϊp4�����LY���*���|�/t䮪�䓓�ә����ʩ��,*�,Ţ
�*�H��Zh�T%WU)����%yt��|Q:Z%�5�� �m8����i��EE:�K����2����<�g�Ż�|]N�x[�V�繄�r,�aO��HG%��?�2[Do����,�<�0��C�qzoYHt-$p�DK~�~�����\^��\'��k+��^�1N�Y6��xm��$���U�����}~��}��:EO��}��N�������8Ϋ^O����u��H�D{x��������<��mo{[���g_��_~�^��X����
��B	_��av�ʕ����Jk[��5%�H �I(С�[���[��k�L�x<�ŮiC���Z�N)�@�=�yj�ۺ��x&�c['�%N��t�]���p���ѡ	#Q/�0խW۵3�ښ��Yh���\di=,��v����f;�nu�lgI��zH����ʖ���#����ӱϥ�k�l�Ᵹ�PM�qhҬ���cv�G�QQyf��=[��ճ�<iQ�xV��n����Gw��׎��4�FA��E>��f��Ȏ������0����b�΂��K#=�o�(�VO�j�t~ ��>��sϭ=�uk�x|���xk^L�տk���-9�n����K@��]��U�n�H�~��\C�#A�~�7�h<WA3K���%s����l�2����	4��f��v.]1._1�n�3���GS�]��i�:�,^���a��:b���)ˑ<V�օ�6ؕ�u���������Ng_�V:��5�m�yf�v��J��j�.����jÐ}��H?����Y�-@��b��U��'�����񲾨l�ot�f�⩜�/߸��w���������`��z�K�i~��S|�k_[	4��o����C��������֙�,��ܽ{� ��F�#㩧�~�K_��D�M]�%�� ��p��a��������t42o�v�t7�L�[7&>4�llʸg��gkN���K䗾v�;��S�5&:���᥸YW&�S��*������x��W�?/g��Օ��+E�u!pӓӆ���?m/����Үme�=?zlvƘ��4��rN��f��g�h�;���-I?yn���!�D��7�Z���g�~꓿��ݗ�0GG���e��͛ e� <2�ml�ˠ�����f)vww��涱e�:\kd2	0���`�<�M��m�ӹ���M�%�%��&� ��3%��"w��-�k��u���^[d��u��I�\�����N�K��보�r����V��6?-�͛5z��BC�n� M��Т�u��fj�-�ՠ��v���5*�}$Q��:�L�H���.�&�ګ��ǥ��������K]0�(�Ӳ(feU.�0���(���._������r1 ��G�G^x���>������ן����I�^�͏M�A$��|ڻ��h��҅�f������C^=$�0SU�Ύ����thJ��t1�ҫ���"�e�܍\/6ĬLw7+�]�CW:�����k �*���<�S/g�W����}����"�&�Gq8��痙/ݴ)��5��6��X�H:A�E�Ʋ������<���Άr��ɺq��^�[\β|���]�~=���k �G!������r������=#������eW�^�W,�����xܬ������H���[�]/�g7��w-h
|����Ix��:H{b�����|\�����:�I��rI�k�c�Yx�?�+3�;~Uͪ���uف� ��C�Dk�����۝w�d&�f��{E7I�r}��\].�Ǔb������Vu�����|g�:��Y= ��#ᑲ��c7�{�����o���㟎��������\Q�O�(<�]fzf�p��yQ�/)��Qi1�������2����%�p�zF�/{3�v,��u���3f���HH�r"�j{ᤓ$��KFU����i��I{q��.� ���HX)��$���� �3� <R����s����Hx��㗾��'���"�Eq0��67��0Xܼ��=��ؙ%a8�]��������ߋ%4yA�S�z�"I�<zY��a8�uW��B2T/�t��Дw�ޭ�_A ��C�#�#��\���ן�ڷ^��9�j��]���?8e�" �w��GR�+s�\�>���  ��   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p!  8�  �D  N"  '�  ��A  �I�   �$B  p������>GJ    IEND�B`�PK
     ˡ�Z,*��  �  /   images/685e2fcc-e73c-46e4-a7b3-171ef11b9715.png�PNG

   IHDR   d   K   �"�   	pHYs  �  ��+  �IDATx��	|U�ƿګ;����:��
�P�e��a�
�ʦ�(�D�A���o��" ����@؃�@����[��Z����d|μ&�1_����U�VW����Su�y\%�2YǏ#�|`,�dymIaъN7ހEKז���C��y(�L�p�+YU_q���>� ��c8��"��%���צF��ss��<��~d��Ԗ�x�P*]�`��4�x�;V�4�W�9��O<�̝��pR�NS������)�{��V,�-���ixc��!��#��e��Vu
d�ĉ8�� ��@�� �-g�s���>^TR�a���U�֖�:p$��i�P<-��t.��j�7�v�^�΀躎��I����5�W{����x2/��>�0gѼ��_Μ��WV�\�IR�p^�?Cyuk�����W������c��MT�����߁⋅�����Ɯ7�����)tk�T�6�=m]n����i�z�[PoU'@�>�';�-�,��tm�$I_)�r��B>�O��#��9zZ\|;�����}�U��n�e�Q�uŁBpg��pFDA��{dI�y�ӏ�:��H,Z��Gu�͚���Pu5:�ȝ��I�U�%Z������~����a��`F�0jh����z�|����S���h�� ��_$�$;�Z(�B�e3Q�uŁ�?"%	����n���Eb ���kV_�����K��������?���c�u6�����C�VB�{QvGG�&j��Ƣ���]���G"��
_�=���
+
��8�3��נ+
$��y��Ƃg��:!G=����6��:�3���U�0F�H��YTr*��\�Ztŀ��b~�U^���p�.���V.B�'�%�Z����Ⱥ��-q�>ThPཾP?/]�HWȧ7"�FQ�`�O#��e%����r��>K>Z�/�	��eG��]����.�ߏ�Ə��EWȼ��`����c"��ӹp��#h��Z�����O�h����f�&B_�*] >� ,ˁ/���$��������W���I�g�O�u�>���g��Y��LÕ5i*��9�] �;tđcY�L��M�?����2�|����nA���YQ��X�%��gXɕ�8������d�w�ȄQ�p$+�&�H�y����������p}zן$��A�h�>#�������9�	{`�W���s��
9��90�e��Ѭ����Yg
������Y��n�g�j̞;{ò�����Yw}T��3��Ӽ�y��1�N4{z4�B
ĺn5��@��`�gT��0 ���>����1���xn�dK�ԁJv�~W顖&;j���;�%7�/�0���5�i�횣Ӹq�/
)���Ϣ���]n�8�<2$�O>���V�[ǉ�{3*>�͊K
��l~��N.��k﷧��XfIAX���\r���s �G�D:��uA�q��KVH�l��Gtt��#�������{DĿ}�q���9�QI�G��m��Ʊ�z�{�l��/5)�z)J�6�8nuBc���T����87b<Ķ�wj��I�"g�*4�;f�T�R �]��^��ۻg�l{�ra�IM��c=5v$�R#�rJ0�]�;���I�1q@��q�{~�3�K���mr��X��]�mq,w(�o���W6���CQ���w"���C��+1�NK�_@t�t���M!��_gbۦM��׭�A��7o<�_������cN�i�ͧπ����O���]�\u��Xu["bG������NNx*Vcmq��R��UN���1,�+r\N'�&�p}aּ�3)\�V�ܓ���?D��cak�᠐y�I��[wH�|'ǲ���ѓ���Ly���++�C<
y"��i<zU����8��{sl�x$j��9$I&jZgt��?_�m�O �֟�)ɧ8B6���o������x�?�'d�~-L��VȀ<>f4���N�:�"���y4n���G(����{\FF2O�I��G]'Ё�8ì�Qw�`�`���*�E�4����N��dS�C��I�%��6�t�i��_:'�]$���,ʺ��M���RH�X�e��]�E;즦GrvG�A�����Ƽ�ܢ��M�x_�����Oj
�%~�	UN%�1�E�,NP�}�n}�	���ԥ\_�*�:U���L��~��� ��}8�`���:yNH�6;7m��V'(�>�Tv�a�������Ǎ`�c�Q�8K1r�X�0�����_��1��eʬ�^7�x㽙c�~`���Z
	�g&N�� ��|G�e�w��;F== o�[�p��oծg����\��k���m\�>j���U�M���켗S^������?��y���/�"�}
L�ik��o@�˷�o@�j��AW7����7��V�h�o��s��i_����2���rn!rm�N��|pi�5vY��0�_�}���6sf�	y�~�=�_U�O�*sOI���?�=:Ǽ� 
�k�p-A#�c
��{��q�u��	X���(�*��şo��1u��ۧ\Gs�j�OH�X ZFȱ��*���e�Q7�k���6b4ޘ�$\��h׾���p��ę�#Q֜0z~>�~�MUa��i�%6A��=;��:7F3�h��n�<8��AX�޻�K��_Q�0l�O�V�T�T:8�O�b�ڵhԴ)�����eaM�b�k]66	S"�>�1!��d�q��q"N�ڍ�������I8�t���ǡo��hΗ�w�����Ś�2�_��:��tyxޣH��JNS�Ҭx��Xʥd�je��g�|�#X���xp� ԕB�2���/}~�Lس�_�����LJ���fY.�Khf�j�Ɓee�c%�48���&�2�	�癢i�7YHS��uEfT�7MS���γ���9��hE�B*�MYJKS�&2"R�R{���E|"�F��Ʋ�Fle���]�
]ד�M�Nݼe��CGQ�
	k��A�#N޺��DѸ\��K���A�t&]<urK,��U�n���8��t�g(��
���\0���9��7��Kj+�j�"'X�N92��ӪVO���y�8�w~S��au)4Z��H�9��w6I�,�h���O�=�E�[�$��VSQ�����?Z��RH����a�b�HI��X�(�\�#F�7v�Q^yWkv��7�QZQ%��.ir2�v��A�K������!��J�Ƌ��Ë���</����g��~5�i�m;�g�0�v��TZ�ÃN'�g�AEyE�����	ԥB$2�	gLtyyQ	��5��ʧeLCƴ�*�֛o���a�bJ|�%��ѽe<H
�vL�ơ���&�]zg`H˂$@��2��V'5�L�_	?>�bj>�j��Z7j��e9��e"�aC]*d@�/YX�����ee�����G�2�eB�x�7ף����~��oGr<Gmǃ4& �2h`�#OG 
�rE3��[�$51@C�@��Q^�ԮK�%��/�$5A~�gI���l��������Th�,�ݺ���W3,��7��|0�[W�j���.�-w���E7%G���q��t{ &S N��808u�(�t��$G��t���KE�i��O�Q �����&R#�z
� j��tsi���4rp�"S$YrUҽ�R!�ۅ�k��ߵcϤk۴�7����o����_����V[��VM��m�"q����A=A�sL�=�k�]O]�
�Ą�.Ư���Ԙt�F{�40c�>�O���j{��p��լ�Ia���!�eA�AQ���ߐ �;�M4IN���BoLL쬢���NG�m�Zf�^�ŭ�oBϞ�໳�p8/��$Q�X\����Q\�o�!^��]A�\r�^�!�Vl�v&�A<0F��������z�uR�~h|X�ڞb�ֻ�lzgNY1m4s�bZ�'�.��w���hۦ^x~��k�i�y<�%�m�;o/ԧ7JOF��bv��@�|4�/󡚶�HNEIu�t�\j=M�Y7��ي~��I�7�5xMY����c�����d�F@ Ѭ�F׭������hh.!52��Wu���1�3�-�p ��<+�Y���.����_�ݥK?A�Pf{h�p!+�BE�Ԧ>Y�@ǇDj�Ԅh�(()��j�� �`�w�ź� b�4�K5} ����Y�r�~�O�'��������� �~�������@�惩���H�'ԥB:�d����k~����M�vg�r�oӺU��ʊ�YC[�ܳC;���n境qz�8�D��Su�k��x"3�J[��25j0%`H������y�E���mrР�n�ah�a�E�O7�[Vn�P�E��ļ�tk�	�A:p�GgyNcy�'H��k4O�s+�:��M�e%�K�|*���7`�S�q��!�j�y�'Or,s2�.�'�����fm�춊���Y�U@�.��9��a�07��(��*,���%U�2*ݦss:��\���(V5����)&T���gM'~k���$���S�a]�1Ǥ=Lg�� �`Q�#"Z�4�s��zb�6歷�06O�+

p߰��<���������׮?=f4���CD����R�x�W����2�����ꚦ�
X�s��a���2t�K[���M�����g4��n���&���/bd4��M�4:F(�?/à�K���e�l���M"���&$ ��Hk��[>����ı���.+_{/�2u�+������س&�����[�@j��d�[I��H�j�)]���	���Ԁ��頿47'�o$�m_8pE�{��y�����;���}4gI���@k����]��W,\83g���ѳ�P�T�@f̘u��mކY��į]W��ty5 	35 	35 	35 	35 	35 	35 	35 	35 	35 	35 	35 	35 	35 	35 	35 	35 	35 	35 	35 	35 	35 	35 	35 	3����K��n    IEND�B`�PK
     ˡ�Z>zG�  G�  /   images/7485d96b-ebc9-4409-ad2f-5f0bda14de1d.png�PNG

   IHDR   �   �   4�z�   	pHYs  �  ��+  ��IDATx��	�e�uv���[{���}0�@�	�$\�EES�Ą���rŋ�����N�8v�+r*�eI�%��X��eQ�HB @f��`����������|�_��b��b���C�t������w���w\��隮WuM�n���U^S����z����k�^�55�隮WyM�n���U^S����z����k�^�55�隮WyM�n���U^S����z����k�^�55�隮WyM�n���U^S����z����k�^�55�隮WyM��ZeY:����@o��"˲�2]���YS�{�K��#��M
��(��y�7�Fg���<^�|6�y5�R�k�djt��Rck�y���%��I4�f�vu�j��UX�m�����k5�2]��kjt��*��V��؎|�,�#�e~�_���AV����*n��%/�;�(��Z�vJ��;zM�Ԙ�y�|w)��U3{������"E�����,c��mY������~V֗���]S��OXj(n�.5���8��.�l[�g����Tw�MW�0��|�S��0Sn��(�?�?��L�w��_�Ԁ���x�啥�:��fӿw������ҦslWʗ�:z>58�3�1���/{�̭ʳ���֟�d������^�Ξ-k�d��+˫��O?��px@g����{�v�w �j\��.��I<�?����ߨ,����
5�4)���=y��'O;}�O?{�����Gf���7ܰ��4�����F���������~��'{0K�[��n�����O<5� hB�%�˩��U����y��Ҳ�Or�����ǑH�����^YɅŵ���sϽ����ȡ�;�~��[�SLe���uM]i�+�uI����5��wA N�ƻ�z��?<��s����_SO4#���jt��Y"����6�xPЛ�S/g���f�Ҽ��k���%	�Ζ$.%�\��پm�$Y&Qk��2�o�X���..o���g����[���v��t]S�3�+W�]KK��wii�{?���mY�7�,ru�����2����-g���e�~h�mi��Ķ\q]�F�F�6�r����0��|`4����M�*�,Jf1}��V��k���b��.�z���¦���NQ�Qof�[������\X���K?y`��a��kf]3F�x������+_9�C��ؗ�������@7�z��\e�F�CЯA�.�mI��-S���A���*���$2�͸���j�Zk����o��x��:��0�$)%M-��"ݍ�����Vϊ׷�ȑr��#���η%K�z��w�<������>rp����kb]3F��t��xq��Ӣ&���z�G9�pLjX�Ƒi���c_�[�~��y�H4�e0���0<�<Q���dI�z&��M!�>�T�V N"iRT�:1_S�O4�$+}�����ƨץױ�K��k���ҢS�^[|ϒK���=�_�?_~x�k,���_ׄ�!v��?���R�V���|C���'��Xzݡ$�H<�p��g�>N�Soh���~+���溎X�z���m�o�[Id3]��#��%�W�Y=]����z=�#ÑH�9]qBO6zC5�LAS%	�J��cӮ\��{��^�n}�O�t���5at��=ʅ�{$�k��G�Ԛ�k3�c�rC�b�T��F���w<�G��7�����h4+O$��Sř>�	��u!��s�p�^M�FgU��0S���L�k��r����K�6���U�����z#)j
�OO��� ��Aw1X_�U�FwM�k��Bq���-�3�Գ��ȩ���cҙ��]��˹�g���c�G�:ۑ[�df~�4���H���P�����-����V�7R��RG/eE!_�Jͷ�
��4�;.�%�C�~8K�7PC���j�L�$)���,E�]��0����b�(Y4��2���t�2]�ĺ6�N�p����U���l�Z����|=ָJ=�;�/,�g^���K2�����+��{�\Z�A��v���c����Oa��'t�:1n@Bx��0�յ�dyJ�$�a��,��-I%I�C�����4�<1���kx�����ny�������'�Z�PW�,���ݞ\:��^G��]ӗ�&�5at+���Oփ�Ha`�H��
�r�2����j�d�B9G#'5�,�B!����][D-G�Q��Od<�ح��k���08�쓚����[���^�tnq��Z4�4N��BX|��M��F��J�X	l��L�]�NC<���5$wS�v�d�l���aF�wOG�z,�uM�k��nݚ�ՍQ����j8�����J���T�suC��25�T���s�|���я�_���&���d������U),c��-�_l��Mi7��;���#�̲Hc4}]GmC!�e닸��nH��G��*E�Ю8��n�hP��\��h,�k]Y\�LX�G�����}aV����讑uMݙ���kt�m�Yi�e�����.Q�_o���V��a��aS�sm��YZI�񯞔�O�f��h<�o�ur`�^��|���Q&��XVW����6���z�M}/k�G�R �BI+�-Ә�3ׯ�|ázø/QrF��Q)���~�H�d�1].����c�6ٱc����%�L�5���]�b��G��x-2Yhi��H�˞�������gXV̿��R�Uz�HbYVV�������8�cf�&�D�h�ލ]��D�y]w�n^�K��R�H>����i�'�5�먁�u�L���A]}�/�ڱ,-�dc�+��`��D��`M���*�+�b*���C�$�n*䌢�ģ���c)�~
O� �����@��-[��ז������m�鮑���Ӈ�>�����/|���n��>A�$��c�m;H�d{���E�;)y��+ك�3��-���R�+Ԇ���Ƞ���o~��(��u�9��"���Xl�H�q��]�x�^ٵg�����$��|��^&1y�-dY��r��X�!�y�J
�ے�z�B/e���(��i�V"v�Y�ḟ2�~E��1���z1�>0S�2WO�v�ٞ�@/�p4��yҚQ��i�n`�ځL��Y��ѭ,~����[���B2G��Z��^D��H���`�mW�6#��,�������UV?C,e�!]_�Zd��Y
�F�Hڎ+��c��wt
�̵4�S8�j���g�;s���RC���������Lc)Or��T�(�i$��$�9#��es�m�aFz��w�,B�R��B����,Qx��e�u��u�I�H����uzsB���ԩ����u��3�ƪ-�wBq�h��B��X��ѽxr���O���<��!zZ�[2���=x�mz�c�f�1Xq�2�qt���Mxf���t��k��n��^��-5a�=�k�t��0�co[��Y�O$ԃ��M����1�,'��V���1�ȁ�~�[�*�z�<Q#�'��j ��I��Ҝ�zHƌ#�K�nv戕D�Z�4��h^�:P�Ff2���P���7�5~�^��P�i��\(͖�0�O0���5�-��kd�bF�n����Ǡ��H���5����!=G�z2J2��zM��)&g06+';�e�#���)��X�#���j����-oԓf
S5�L�-5 ��i��x�+�%���
�`���[�BP0Bt_����P�n��Q��.5�
}5b�Dk걚R���fj�i����Xs}�����u�,����qr�|ˆH5��6��fl}Ͼz���F����s�`���7N=�5�^9�,�k|c�ݡ���Zh�4հ���cz4Ժ 9�sč�ؗn.0?1PJV6����UK����p���4�ٺ��l�<x�X!l�0�(��{/e�O����,��\VF����������T���bA|4��p\��Ņzp����5=b���*�z$9����u�����PV�3��z��z��Q��K�����������I�8��� �S�2]��zŌn0D�a�8&OrY[H����'7��v�M�<���?&!��"fC_���n��-��A�+�����Sll�=���FE2S�'�k��xR�5��]2�r�x@<k��I�Oq :�-Y�ָ*T��NU�
����^X�Z�8�ߡG�0F�I�J�`W����ʨ���t0���b�����,�8f���'���t]�3�Ѩ��V��y2@V�C���f��z�%���,HƬb"���R��j���T�
�q�\��ƅ���m~�q���wF���($����
5_=z����Ju���j���Q�0����+X���xP����b@Ӫ�!�� ����l���9M�[�4=o�&�q�Iǡ��H��c �zW0^�Bz���f��jl�SV	%Āv"�uM�W��.]*��ϯOA�R/�T�bLf�7ֺ,��Ci4Z2�Gr��Kr��nJ��ZM��KM���t9��SS�G��x����-�b���s��Yq���d����1BKr���ۨ�zz}�~�@�K�/2c��X��q��j���tW��sz[[=�qDȢ�1+�����.A��ׁd?Z�l��YA�gj� �"�k����C��8^0E�4�x���t]�1�,�23G�YZ'|��Y��^3�.�v,0qǑ4��z�z ��I�^'��;@9|s�j��nW�� 1�Z��R�f����\ K�L��#�f�"���7��yD�X�Il���q.�8�c�U=�D(}b1xf��x���dƱɶ2��ж�f3�jжQ+bh�À�MmV��u����Pް�J]���8K@fS1�F�R�8/��P��Зܐ�&�+bt�a�#N����5u�y~����YG}sP��F
[�P:����ÚB��A�>�͂��^��`ha˼�G}z:��I��I����($�k|_=&����1b-z7K�Y�X�5z�4.�JQ �A���,�X� I��L3*{�X
0���+L�#��U�YI9إ	�JOS�d"��J s�x9��[n�D���A�F�=�ǯ���� �w#/g�3�
���hϴ$Q�=S3sdv�i�#K ��b�(
�\�ʨ+H�4�rG��u5Җ��:7+Zn�}�(%�u���/�����c<�}H�K{<����]
4�*��	<�l��_����^ �
�xS�0.��&��a3 #����X([���V��n@.�T _{Y�T�O���斩M"y�g.�Zݯ��tOL[{����]����WB�̶X�>��3$\0�¢�Y^��fG|����=��Xss�u�{_ ���Xt_��P�L�nZ��Q��b���U5�����9ٺ�%e,a�#!�E�I�Y�`J�3e�^Uz>ą̆^��,I�d�!sSf��V�K�m�mI`�)�%װ= WYU���Z�����v��kb�"FW���������l.�l�`�(b(���er~��*�L�T�e�@7���Wf�`�0�Jx�eR�4�m�z#}�N���F6e �@z�kF����Xd�z�T��"���ų�<z��.���)L4�Ȓ"6�6�>�$�Sɧ;��!aC@��Z�W�|FI1Z����#��ش�{�I���ϐ���32읓�έS��kd�"F��m^鋣�%�����Έ�.j�>���bR[4!�W��<6�4�5b;�Z�a���k�&��@(Nrvv��ȹ(�!|vݢ�Q,��d
I��oI��x�s�m\�hݕVݓz����iYaX545��`Jr"��1f+J�t��5�{���"�\�o��A��r2�.�4�>c�~؋e�FoW�����D�UY<wD�ݡ��2]��zE�.���o��0��ҭ+�h�Z���m4�)�~�J���4�O�ix��1@Lkbpzþ�*A�LԷF���p�'o�/C�0	�m�I��+4��/��RWV	���^� ��5#���a)kW�qg���m��-CBIdG�@�S_2t�+�da�`f��*CIo��V)M�<���Q� �d9��T��F�!hY�z��S���dV2]��r�޷��+���>��>MC�ߒe��M����^,n����-�H0)���<����q�B_|�j^���$�2p��k����]�7�/�총R&CKM:&�A�7(�����D��@O�=�@�X��$@'=5�A)�F���]�K��6�ǌ�r�w+��e���d803
ֻ#���<q�.p���2�BxV��G�JBF��P�KƟ���x���rĤ�B�(浃��~�I:���u��]c�|Kͫ�E��7��t]��ڳ�=E�%I�PXv��ܘ�33	8�K[�QS�!���x�_z��*���������?דf���qM
{H-I;P��#\�*�nH�1������nbt�����k|��XHv$�?�tH\[7�|��>���aؒ�8!��ɓԘ"�e�$L��q��ʕ溬n��P'�M�#�����!��:)Y�V�k�k�-���F�D���蒤 o�R,t�S�hSb�R�~�'�KKb%	k�y%j��5J�޺��u}9~��G����??p��g8��9u���\�᡺B����Zu�5e�x`��#�J{�h������2]��rG��H�:$�Z}v@� ����se����c�[��͐Y�L�Wz�q. ���a-h��Y�t�;���a%m��COG�d9S"�*i��Ă�V�?�͟�h�ב�Oˌ/�Q4&>�����D� :�(e�޾(0ݏ�$��z082�lJo��ig�����Xz�H��HPo����Q
a��=�"�BI<ޜW��<:�����	1��	�ϵ�Y�z
��}��u�:
uqHdzM���"E�X�>w��Wy��/^Z_r\GyQ�=?�rKDh�Dl���@�(w�7W /27o?v�ʕ��ٲ�L�k���}g�Q1�"�)Qh�����EB�m[�tC����*WV����}�gD�@O7XoIkv��2�_��TP'�~���s�v�Mk<���Ma�:��Ϩ�U��T�o�
���zD�!$y�|��3�%�5���s#�æ�k@m���$��B�j�a�ͧ�j��>N���#�g�֖ 2����<d#�Ѣ� �Q�+���-'�pY�2|E�ǁct�s�e��~2V *��l6�@�����=��a��\Y)� j������q)��O�h��98u@$غe^���y|͵;2����*V^��߷�uD����t���E�.e7��.��L �j5_ΝQ���\)o��S}(uw���05��`�`�0ݯ�E7����>��z���}�>�Ĭ�!W����À=��ՑTVŁ�8+�ⵘ���T���� �#eM.�%��ǗR���ɠ�Y%;����
��3��^�$ѧ�P�d�>�x42*_�>'�d�H"^�|@߀^��QtX�t�����@�!d��A16T{�_k��<�xyE.聈@�Vt+d���TvQsE?g^fg��qȁl���f��k�ܼ���&I�V��ɞ=��Y�#����P������_�aF�$Nk+3�S�2F���j�bC����3V�.��~SF6�C"�#�i���T*ȕ�����z0�wy?�� (�y�������j���r�	&Oc�En�]b��0 ��J��2qct�D�g�g�>� �ƚ>�.�U�4`3~o�����PA�^�+L�g��Ʉ�Y2�����A�����
�������R�F�|�2��;�악�}}��	�e9CO�u��|q���7c��t�f�MSoӓ��M*!@����W����0��/�����'�,�V���7�n �PLR��BK�7wB����N7�X�lX�7�&ɔ�����.�r�X� 	qC=�f�ht�Q2�1PR.ʉ���@.&4ͩ�L�I�!V�Jcxe�4a_��H��¤��Wc��HM��K��
�6���*�r�cFtш��Ɠ�Ik�r���z�k8D����/������!a�!3�s����l�΃ca�����qp����%ik3�H�ɦF�.��s�FP�5b�s�\�B#�A͑��{;�>/�3��rbif)����S,Y��
+[�;�RT�9�Ɣ*�A솎�qv�:�)ZT�k�q&%v��񄗹i�1RE�Lәm�J�Z2DdK!e�H�I`.I'��]�Y�FX0:�tINF3+�3�a�X���c�#3T���0M�bHԆ��O����4�׍n��1��Q�c��Y3�a'���F	a�m�
K��lK{�n:9�L��b f!���oV	�ϐhQ�Ҋ�lY����'d�^��8rB���{��۶픰Ѣ�@2���+�Z����6����$BB$��@'8ăB=�5V?�xڇ�@!�%~=`�����%e�$1�u`!��3��g)<RO�.k�c8���qn2�X����9=��YRx����Y���l��y�"�j��E�#<>S�Ϊ�<(
������o����M���Ě5^�SE(�e{˪��*�M�F��w�s��~oF��z��7N��R��ǘ0�1K[�B>��e�\����D��5[�w�;�y�F�\8�(KK�,�f��X�5fh� ��������9��h �4���'��	]�,���;pA�/7���2`���@@�	/������FOa�z��q.3���s�X�H	��2��x2�*����l���#ǎfF�|�E/U�kYUF�p�4��z�L�;����Ax��q@����� �,:l2�=x��bGk��y�#����Oa8���Cb�V���^y�H�@���d�|_�F;���dn���ޏ��re1��~��>�cwe�9��J�)��5Z.��G�X�f]�k�~���,���1g�`̱��jԆ5���Po��/���dތ�<�M�Q K``#6�S�J�����k���b�RwZkf�1$����	�%���!����p+���t�c(=<'��kgYF8gF�X�j��ϐE�� q�=
����)�rJcd8@����H��#���Mư�txϦ[���M]�j�'U����tMg�>OMc䭳s�]����� +�C�iC�}+u9-��ņ�劽u�4e׽f˥ �@8h�^�N�AT(�YЍ���;�b�/���4�A.O�HOݨ?fFE�r�A_z�p�zR�5�C?b��g<Y��	�l�F'�e�;�Y��O�Nf|N��͋"�4\�F���Ùy�FJ3���a�^G�WLiš�~nn�/9D�!PJW�`��K!7�އ������^}��]�-3�5�VV������78��On#XhYC��8�1T�p$W��@�l����z{��q,a;��`������1�,q$�V]����2�Z����<}�u��^o}�L��5[.NF�9�@�Ը��z�_���XEb���`���Z� ��:tb�vՀ�F�����Z�nd�d��Ѩ�w��=J@Hԟr4�����zR4(_"&��95Ƽ.z~������T��q���όM�����bӳ���>�4P
jLd��6f��<�mM[tPB�+��5Xb�YX�4��7[��,*Ƕ�I� �U<[�F؏�7$RRJ��-KxP$����P�.g&d���x���K�޺BN_��ĭ(�#��� .��{��zM����̞E���NX�e����I6z�۸�-��+3Z( 3���,�1E����� �6�T7H���q�
��r����������k��B���ׯ�m��A�0%�d����W1R>��p9�-ҳ�z�E�z�1+u��3Y���p�`��FT�b�;fVR�a�\G4�B6݁��`�N���۠'Ъ�27r�U���l����2�s��������>��%A�7�~w]^8sRz���G6�0a���\�_M��6�O�f�<U�4����(�[_�7d�^��b#��-�����:��R��z��}��������\�u�!��0#�$PhՖ��ش��U���E��2��h��F�W���n��p�|qϕ���~ L{a]�'[o��qZn�aI�����v:�_a��z���L�ڔ	���' ]A��t@<6HΌ��E�d}}�p��j(lV���,pA�o1d�ħVh��XZn�gx&�:�/�v�������jhb��1!�m��_�yz��ٔ�G��^�,k�+*�޵�w�N����ro������^�b��E$��`?��e�^���C6HuЂ�57�Ax+T�f�Ы�Fu��.֊����02y����\��ri�3�=Z����Qo���d튯�֒8Qc͚F:����H2-�I|g��08�ޔZ�R�Rh�
�^�[��Ճ!l�iؼ[�l�6�K��1��O� @�&e��Gh9�7�j�Φ��h()��l��\�+�8�)��[�4QAo�ZR�rs�)���gQ:��:]Y��
���Y	���z��W�~���g���S�iǶ-�o��h?��g�_�#�v� �����2i���
�1��e�`�ղ}ü5��{��zyD���k���U�0���GO�>�XC[l0ن�G�ݒ�K���33�^n��d�yٹcA�z���n��4ج�e<�砾�j6 5]���B�p^]�#Ac�J�����0�
Y@�B\�ԛ ��M�%tw0����E��_ϡX�Ϋ������Ư����_ِ% \�1��i=h�A&x���ծ,�!Rcj�T+ذ*b�'��Kt��:x?hw��Y�׉Wƻ�9
jw�q��u�[�7�%���*Ҹ����ҨZ^��HU G��������J�C05��`�Ǟ���k3k�P����$����1���ukƃ��U��}��� 8��U	����`�W(��)T,)�����V#�F�4�+��DnL0,,��ʺ�l�)eS!f�����x��"�'w�é��wV���a�j u��uirF��`Y���1�`Բ����KN�����c���hə�JSo�T��:e)8<$�*�e��ia93N|,����$gVӮ�����Y��.xE4��p�=t��v�\=oM㶑 ��e��M��4��L�1���5Ba�ٝ�e�^��o�t���u�z�7�I�8����ؑՕ�[:�p����g{��Lb�m���3��2;����kW����c�L�
�ᒛ c�чP+UUu�zR+��s3��י��,��W����;L(P=xYi���k�3S�3�?%�L�*{(U�Ͳ*�Iה"l#�@I"��>f8����	?���v5Lh��yđ��뀎zd�/Ō����tXH�X�g���z�"y�:<��:�dw���҅+�~e�l�(bD>Iז�'^qu�W�#��L�x�6c�R?���C��{�>���t��˅F���F�}0]�L�(d�Ԉ�]�PF�>��D�b�eT��͟�t�t�B�J<�͗�_����~6p��%��p}��<N�+�?G!����Oc�a��ȓF���a='?$ج��bè0��R#9ib(��nr�4,� ��͜P%ڧGB�ͱаt�&V��c*�E���h��:20c�L��!��lY�|Y���MO��9��d�ɚz
eS���H�'������þ��&{�bQϥ���`(�P�&���~��|m`n��ƶ%�8.ة�&�"��K���j�ҟ�� 8�aBW������rW/3�?37���<g�Q�\����T]���M�����'�!{���4����2���ikc��_n%��dEAuU�3�HqQ�6^iyO�yl����l���q�Ԙ�����4�MzL�őT6����n����I��̄џ&(�+��Q&A�7:b~u�Tm��	�M)@��H+�His�	��S��|��v/���F3�͵����8�G��ln�º�-yj���饾�:Gy����T=�����`n�������
�,5Ժ��m���+�ZF��߭�"���d�&�B�I5��xL*�8HtftӋB�(�S��D�X%Sl��;�]�5�J��BP݈��04l��I�}5�8g��+�Ș�b�P4�I�j�3j�zr�DQ��0��40ӆ8,s���)ċ`̨��L<G!�cB�I�Br��LIs3���ԃY�X������f#�nc�ia��B25�uY�0H<�\Nq�ٴ���zX��K.�{_u7f\��*	�/q}A=?������idq_��`����e~S61VY?�A�٪�g�ׇϯ߿,��Y�ڞ�%���,�����l��<�1Fb���Ɉl��Yㆎ�S�`_@~ Ob��;�t+�s���Rk����u�˜�S���6�E�p
�XcI$U|z:��0�����]���d���� ����2��tV��M�O�>�RF!E��aʝ$�ܰ:��M�Z%}ʠ'�03UX��U}c��bC��!.)Cg[e-��	��$q8����8O��"~��?$m���&�,	�#�4�u��,2���@Z�sR�0�
��q��fo�r)�w��s��1��gz��Г;�K�����.�,��!ܘ^�-�F ��'腆ֿ�:��qZ"�G oپ�k���~�[Q7�[%Xčd�q��50Ҿ�P�6���ǂɏ�geV�@X���ek�� ���eE6Ԯ���ªF�4	��&Z%y�x���ʪ:P1�3C����I�]�ۡ��ƅ���]��-=Rnz���*��T�kāR�}�6�6Z�|Bu�6Q��TUL^-��5^c���ڌ��c�(e��2/nf�S��ƫ�̀�[����52*������� g�G�4���c���y2]��r�Z̙إ�TÙU����K�e2��2�k�mbL-�c�D��]���rX���c�nٱk��z�܀=d���ڙ�ЛB-�.� B��a��*I�r]����\Z3JWEg����:�ީ0�G�Ic�*�uW����="IB#W��B,)���:^�0��xl���7=L�/��1���<7�˪wu=ݪ�G-4͍�B2@�0Nc&���$z\�����a.��I "t�E�8�]��� �(P�B�(�_�{P���S��	'��5�|�Ȑ�6~�[2]��r�p�_�����8-�q.5'X=��kY�������fR��n����_\\Z�qP�Y=���n/���+rݍ7���]�����XНk3=[�pL����D������¨.'~��|�c���W@[T�'u7�%����R(DC�<晃ΕcԲzD�=x�T�ZW]�Ф��I��!�r��0⪭�*�.	9�I�9�#��:2��>��H��0�M��LI�`wy�̎���B|i���<}^�]#1BJ�^eey�=���Bc֗���e�ܼtZFjemC�{�>�tE��Ӆ4�AAU3ľrY��5Y�O���S�ly$a�n	�ӿ�� �*�i�JGv?�\7�<��]�<�t���ufK�?j�������?��G=�k��l7�i<UF�*�DV1p��%R�h�u��ĈQ!���M��&VL׵�(V5�c4������!�	'q�#�:ҍ��Bf|U
]z��m$��Q��'���X�ۧ��hv��#�0�����Wv���N�S+F���>�����A�D���r��y��Hhh����u��-�I;rE�1���fq��|�X�J��]wݶ۷m9�%Y������x��UX6�?Ѱ�=?��h��-��Y�U��v���p�=�-�����_��{G���ܡ�bym�^ϕ���\\W��WCsU��CE�j6?����c�����i�Śȫ�~m��eb@����H=�<�Ma#x,lp��j����x)v��.������l�U8Jӌɪ����E�e�.H��H�4�'bq]��}���6jOz]��@V7- ya)t���s{d����pE�Г��Nb�4yx<��3�������e�e��_��P�Ŷ,�����Y/{�d�]h0T�6��Sum_�����x�m�֨]�(���E1Tχ��/ͺ��A0�"7|�'�4}v.;Hs�A��k���L�L��*/��]^n d ���TVa�gjf����0^�f��e%v��Qc�`<HZN^'3���3J�P�Nr=\�̴�7��� l�2���W!�%5��u���
7�������kjp�~�e]`��V^$�F� y!fk�u����~��Xƫ�,_\��o4��	=?��Y"vjԒ�G��</^&$�MmL�F豘O�b+ټ/z�&Na���8��5�xhcBR��Qk��.ؕ8��m�K�/.���EO͓�0V�����WbH�oj`��(b3�$��H,�1�gqոj(f�p�͙z��e������L7��G�4R�����2�a���p 2�¾(�,��Ԃ\ڭP�:�;�����5
��f�'�EΦf!�z���:��*_�1�i��M"�2]���	����0L��l��"���t�U/TV���o�U�70��y�k�ӎ=���ʆ�Ö�zjg�!����t����dֵ&�uM��mtw�t(�J����%4	���Ai�C@���c��/�;�Q|�}̲�q�T*��Ω<�]aIWU��PO�*�תa��,�،Ð��_�R �S���׺U��7B�=�%Fgm�L`RHO����i�f��db����52��;S�T2z��<+���J�줧C�1-kt,������ӑ�&�+��J��L�9�T�r���R�Øl��a;�������~�=�<�G����a�W�a��w�<C}��wUk:�S&Y&B�FQl�Tq+����ҿ�%/3S�M��y͗J�o�ĖE公JK37B�n��g�7�xU]�������<z��n�A~�>*o�wI?}��1��JA��]7�c4(O��2]��zE&�Z�֑�K�F,'��0	R���Ziͧ0j�V�gK��%Ewwifȁ�EmKת������1�Z�u6wR��2�ʉ��M�#055�s\a�����i�)Kv7�jW��|.�e�7���gJ��~�\�t��5�~��<��,���S���J�7lz}���y|n$
A��������:_��gsn�3Ps*bJ�gL>��l��Q�}�u:K4q�Mv~{�Ö@��w�"�1�0b������Tx��tn'���FT��G
 �;�����L�
��Xѻr��L#���,^��B!��cL�W^�j9�ĜW�+���`�Ԗ��ٲu��A��'�:�w��c��Q���i(Y[C�9�fU��u�^�ѹ�r̘�	���j�a��&���Aq8-��8�]H��c���o�n�ǌ���=����K����d0���lI'l�Y�/aPg��I��9�81C"�JnԘ�z��R�@����[�&	�Q��j�zg�	x�~(�}�����ٵ���s�K��aZtI8�ղ��a5S,�\>@ۅ�f�7�%��,��U���<�*S}�����x(�Y}��KG���32]�����.Q׃��urS$�²(#`����:��ll�`�D�������g�t���"�/ȓ�?.��<ٹJ�=�bz�RCȌ(�4�s��m7�9C�+�6��V#�bMM�^z��.4�a�$���ffZ�[�WC?+�/^P�ې�>�O��ߑ/}�+{~E�-l��0�fP�l�Ig�]�e���aC���w��ѐ˗/�`��xQv��!�=��&l-3�"4��P�a�������V�����-�G>-��W,�����z�F�3WQ�Jz7�R�B>xP��I&���#�n&�L�S�����O�;,l�"��y�=��<��c��Si6���wߡx��� ��C55���:��\g����nӛṐſ�7V��B�[W�א3g/���Ң�w`,G��G��0�h�5+��Q<(+�kj@c���M�=��Ğ���a�l�H��&��2����ި��I���1^K�x�2%��k�o�R�!����"V2�-dm�(�79n�Cez�g,��Ge�^W�I�8������d�m������L�ϭ��ؐ4L��Oj����k3�Mz��v����ú��1>��tY�x�m�o~���>��{�>��_�Uy׃ʾ}�d۶-|>�I��>���r��obqR	ǎ</���C2W�(�#,d<��Xغ��g~n��^|q,o��-�����/И����>�I������x�����6�*��p������/Q��,tUȴ���`Z�7�(B�N�i�]�����I1��ɣ�o�G~��ڿh5�^��z]��_2@��t��	7�d�HI��d�����袷˰����k���J:/��B4�ҡ����._{��z;$��|����9��̫Q�n��~Ǎ4�}{d�\����9/������	n��{�|��19t�I���w�M7P����~K�jM|�~y��Snq�e��O���������C���.�����r�ƽ���Ǟ�#G����)��q�<�Ň+�ȅw�*k#j����Ƽ&3Y6S�7�4����b��_�P��Cb�Ϩ'�=T�KLϜ��ͳ��'��{��_���;V{���h9u�T��~aV�r>J��|�FQ�Ecj����G{I�����F~���z��ܖ�f:����X�N���l����t��'��eEU4Y=�XXf�5��Z���A���B5`��M��LDxU�%�m]�x���++K�#�?�'�����I1��-o���ױ�G�?���?�^���� �5���'h�<�vy����?��_T�:��C�Z]_��e����˓����Ɛ��!L�s���{妃{Xy��z��َz³��p��a�瞷�^�p�C?úU�����א�8+�Lc6�����(D�K�0�I4���!�ݗ ��h�Uh٨�o���/Y�����̏Y��Y�<��33��|�{N�<�����[~��ϳI���=��\�x�,�	H��2�U	����r����ܿ^�_~��۳{�n���������k|�%��u�I�c���6J�0��� ��p�e��FD���.�%yD51�r
'�aDu�V�-�Wc�*�\+KK
5kr�-���o��'N����>�)�|��9y�;]y���F1YD�g����|���ozӛ��$�������΋@:���q%���.�vMc������_�'��e��G>��}�χ���_�|��q�ʺ�H�fG�h]��Hi7|�.�F�c�8M��.Y� �u��q&�&�Љ��5V��8����"�ھ=΋�H׾����M_�W`=���[�?u��G��/����x0��k��%�0FF"8�\��'�)�m�e�w�w�_Y�X�{�ԑ#���#w�ޏ�ȩ]{�=|�-�|���o��q_��yn�q,c{YE���I�xnX���i�$�N|'�>$
ǣQĺb'��b�jb��er��)��?$7����nT�!�~�0��-7ߥ�唜R�{�>,gϜ�~/�z�Q�y�l�j�w�x�I����e���e��M|ǻ�ıs�`�����i{�
���y�R�F�L��`N>�^�psM������n��_���O�[��6}�}r�ͷɑ�q`d]���)c�&�5X�dOs�mY�p��2��*����?O�$�d��Ӄ*�C�m���-�o���3���_��f�w^�V��}�3��x����տ�P4�>��HY��^��M[���-�(j�����(^W읔�qksF&�B0=��8�qw����+��>��3?���������������D�����.�l��;���=�'X��͕<�)��@�$�Z@�̱(���FV%�~��HQ�+_��]�M�w:$�n,\/i,���'d4��`tL���ē�����}�sr��yY]����{B��RK������V��1�G����y瘲�kkk���s�|��/�Fo�Z&�1��&�E�r���,Zolz]��{k����Sr�}�ɞ={��?�x�I�V�PTJe��"5d�QoD��(/��'D;��r��v�~�Th�3zM=*@���Y�l�~��>A�ð����,��\=�c���������xbO���u�ҥ;�y��������o�G�P�̒��2��3�]}�	����G��2TJ�A��3�JS���_0��!��!Z�\3�ѓ�p��V�1N3v��a��8���>����'�Σo{���������:_/���J뺑l�T&�r�"��:��I'@E&��b|��U]j���ݤ�<�u�
���;>|X��!�cݬ����y���
9�'�8d��t����IU�3�Ы�л�ևx롇��Q�CR�3��g?S�<�u�uĖf�2�$���d��1m���_�>��pm��"R���u���uP�CV3�d�KK6��n(5FKì	�q���jb$W^BM:W�Tc�9>ϤG�P�1��ޕe��[.�!k�mO���v����<}��ǟ}��$=�����f�כ=w�����r�����(<��8R�a�8�	xc��*�i|�5����J3��E����1_oKT(��2��)!Y�!�F})쁴f�;�|���N�:���3?�����G����}�9y�����Ls����23Iu2��p�D��U�d
Q00$�)���(�ￎ�
�~��,�Z_�d"�P2���jpyiԻ�̀�P��,z�Gβ6�L�D�mfff�M�1��5����0p�։�]^������侓$OQM�1�6c��D:�cU	O�k��-!{faa�����e�T�J~Ne^]�r�\��G=��7��X��.��𳴐��+�w��,����[�ܡ~y�J~�����=��}������A[��T�Q�fMa���n����a%/��F2H.�k�������� MH1���B
��K%�	�,� L�a�($�������"W�A�����@��S�SH�����Y��gO��߿�t����/�ˏ������c����d��ʼ�]#���ʤ�O���l��H��i<tT�ģٙ��X÷̥��b��;�� Fì�\pP�����k4�I�O����Ǟ�����ڠ��]C��^��fg�8'��U'���u��Y��>�|�:�+u}>�R,�������VC!���9~>ƳY��1�T^�3���!"�
z��dUw�bH�$�RFH�!a��!&�A�P0�V?Ó'����=���.��z�T3@�Dar�����K��"��A��[wf��;���F=X�ޙ]ڱu����̆��]�����ڪģu����M�܀h�T��c�&���r��u����X���B�ԱQF�evvN��ҽ�&~��uY�p���g~�ԩS��z��~�%[^�ѕ���^X���f�h��9������͆�f5]�^Սm��.d�|G���w���-����ۙ��ONx�ZТ��d��Rӹ���bT�&iixHx��f�z&�Fx4<�p����4�Ʃכ���v�v������Ϗ�
��"??W	�	g�^�J(�����IY]]��n�<�=6�%��T�	-�4�K�\��H.�p^�ђ�^�V 3�G�0����R�p�ל��r_�~��{��k���$�7o�Q��~����
G��zp�S���5�Pn���o���I���x�v�o�n����/��@�ۀ���1��"���$�g&��F����M�k�B���+=���̧4x%�t�聲:��~
�W�=���[�U/�9�7>�;����_�⏿廾뤼Nַltey�9�^�����_�E�f�zS�_�239�'�)e�A"�c�u�-7��b�HO�P�����c'��o�m[f�E./��]r�[�"�q0ɾ�h ���a�o���X1E�������?������S��	;�;�����q�|��,��f��;QZ�u�`���=��:�!uCv�20բ��ȕ����W�h5���K ͼz.�<5"'w%Qÿ��yq���bH9v3x]FO-`bb�{}0��i]��¤���(�)\�J7��3��Y��:��'-��V��i�)��ݯ>��O���c�i�[�j�w'�߽z�v�^|��kG�^4���"���=�Ǧ-ʭ�TT�����શE$�CF���2�:�g�(�l��%S�)�ƀ��˙�'������3�����z��N��`}�FW��?]D�ϊlms�P����R?͘�6�M��󌝢L�`Cq�k���pGT-���ڕ����8�{�ַ�#����r��3r�7J�U��So8$��x�n۶m�<�m���ƚ�ܹ���s��z��'�6B��~FVW�4��5ɺ�9�l0�	�l�"8��
V��ܹ��}��%ٱc���YY1��u ��,��(�6"��{6cAd�h�ĺ�/����3�+b�2�,]Z�0�+l� �4�
'[Rz��GcY�k��ڕ�zܬ��LtC6q`�����$�PE�ʆ�}������]5tk�Ƥ�����[�nsؽR=Ln���s���VK���%�=a�W�y�zp�rk�-7�"~���l�8�7ү=˶R7)�v�l�d�-���`�ƗԷYS�LC��`���(͌?�}�LF+�ҥ�o��?��o=��C��=�y^��׷dte��*6}��m��g�U���>U��mOT��vQ��TJ�O��M�����&�5v���ڿ�`��:6�z>�4�o��.�����t�/���ߠg��'����_���v�-�j'Nc�x��ٵk���ߕ���U�¢<����������?�5�J�7�}J>���������O����Y���ןxL�r�[9���ɓ|�g�}V:��k����,�'lj��bU��	�Č^�l`�LQI��Y��:f(h��j�)�(�]YW/�rA��5S}���k��j�H�{7�#��+}�B�����ju��!j�zH��i����סޯ^ӟ����l����dY	�o�L��lٹ}�eǞ��߾������>��'���=gy.�r���7�x���tiq�m�BȾ�-�l`������B�	2��Xt̠�Μ��s����9r���v�@��׷���%������f$<b���)C��2&)�xč6�k+�Y�?Tj����������`��A�R��ý�7�W�2�����az@�zïb�B��ey���FX�8Ƅ��u�]�炗{���6�p�MD�PB�������?��O�G>�YZ^�믿��܎��PP��r���>���J�F�� 043<�o�hH)�%Dv���m�\�ҥ���"�7��ܼ.>F��2�Y��1զ����}�x��t�
�	��Eܩ�0š�pF�\���%���8S���&����M�}���s�R�k�!�%�Ʀ�EF��}���X���o�R_])�~*���bן����u�����-e}�c�C.}�S�q�٥C�(�vj]"�2�W�j�.K�hê�
Bk���k����'N|����/�K��ߔo���]��^���l4���U�k8_@�	w���PN��	��3�3�X�l4�(��%v~~���ؑB���7�av���p��t@?<qߓO>��oݺ��Ex׻�K^|�E��&�s��L�c---�!_�� #Ey�[n1������������(�>wL��Nfggy� R�9s�1�w�nZ�Ą_W�xݪ��(���J�e�.�Je^�	�5=�G�i�X/Sȅ����e�`b�/��<"ŉnT�@�9��o�[릅:5��Wl�Q�kk���E�;i+�n��š����8�2�f�I��!�8���3k\�,F������]���?6����^<��������ܶa��U��<4:�m�]��=�>�R���ş�����?�ʏ�Fr��56N9��C��ɰw(�!�9����#��=��/^��ÿ�����~���t����,��d��@��/����U�sj�~j�����٨Z� M��.謦9J�A9����G+����O���}O5F�0K�˚
��Ѝ�G<p�~����/����	�'���5ȭ�2���&�����d� ^?��s~�Tϱ��6���63����V��X�ԩ�sm�
��*R �sad�a��K�q݉R��;�dF���ر�$\�h�5��#ֻ~�4jס�X�΅����ح��P���S�����j��5��!����c�rO'(�#���gS��exg�Ϥ9�8@�r�1��	|�yͤH��}eo�_�;�?��^{n�k9+��'ϧ�ݏ&N�_������'����oزm7�f��'ơ�P�s�حP��b�m�W���na�~����O<�_��}�i�����e���b<�LaM�*ކ�7�͐�2���,V�A���D����do��|�>X��0 �t�tlP�aR5�����ML&r@�W#�+�T���o����K�B8 ��=��#�8~Zv��)WV�*g����,��`����&�R�&<���l^3C6�n(�#E7��2P�&U	�(�E-�Q���В��W>����{x��*m|�zz�����@ ��DQ�b���8�ofĮ����@AD@�"�;DBH�@ғ�[r�=��~��}��Z�978�|C���ޟ�Kn9e�w��=�y�Y�i1ߕ	�C!�Vh�s�xA��H��J�X��C���\��!i2BU�!��Ѱm(K6JT�g�n5I
	L-
a%�@�#FѰB1��&YCbI
�t�	�]�ɖ�����/��/�a$Y@�ZHm���1U%s���-@LC�Z.@���Np�B �:��oქg%�T!�G���K r��2^ߛ�������K�ex��7:?�4����ӂ���%��Γ �$��
21] ��ɔ�����Q/�F��;5�I�.0��}�*P����<RE��E�Q�~S�ͣ ����b�xM�@e"٩��}�\M<����3Oo���o���]�him�{ｏÖK?�o5�LI���-A��yʴ�=�E���`��1�9�$�IE��&\�ok}4;X�>�~�yd�f�<����%y,	'�Gg:�!����rF����y�( 4��L���)-MI�����v�]�ft�x+ѫ��	��r)?KA:�j?I�р-�Qc�%=�	�.7'�103T��{ǜ=�h��Ƭ官�j1�z=*��`P�U`�:��D�2���2�J0�3	�-M��4�؄Ie���|A ��dxm�D߈��I�?F�b�#?�����K���:|��*K�,�����0ULP�$�K��X���]�� AJ$�ҟ��9:�a:��s�A	�ӆ��LP��<�@?��2S%B�ze�詨7G��`=�z�7�^�^��k&�[���8��m��:��PcZ�\�r:6�Z�I��80t�7m|�����=m�0�1�$�]nM�Xb�J��B�E�=>�8������ф�@��{0�sd�#k,V��n4�^��zx1�hl8��a�}m��dk2v>Q?���F�s��C��?�|���)Q�
Y�c�
�44�m-�_t�)��,��]P�ȜnT�6�p:X� 
c���4^
{s&�ȸ��	1�c��0E�G_��F�Ii[6�\s�$h	�[:^?ìQ� �
Q��"�>�b䊢�0]�[3��(�ʝ=�����O�����a5�!ӻ�ǍO��U��l�A ��D�ZP�hU�{�Vc�P zQ��~�F7�D�/&�NڝiI��XJ8��0,����)$�#�)U|п�����C�!�_�:z!O��
exn�fز�ynL�F��+�G������c(�1�5�g��v��#��3�=t���$!a�SSrT��>Cq��Iт/��I'/������4�4�siJ�z�>!�I�!��BUɰ>K��̚9k��%K�l?��-��r:��'HF�<�:c�6�����w`��(g&a4�Gă�𒤑�a����dKCz���r�I��k$$7ط�##=��i�B����~�*�4)���1���I� ;����<�[d��q�*�
橅*�h����Y�A���R����~� �F�b
P��"�((Q4�(|2a<�L�OWk	:��ccco�o����f��n��ӌF�t0P��5i`O�I|I��� E9���1�QIݭ1#ө��_�<�y�ͨ�YR��9C���2
�
4BV��m.[�x<Q+v�it2�xa���\o=�-0��?��<�a}�gw�b(WP�ؒ�i�tA�^�U�г��t�C�t>�U��j-,���3	�!��4��S��<-A���}1ag3�'���sh�0?�B�9BU;��T��D,���ս��e˞:�MglX�x�{c���zxgP���A{��T@��ٔ����&h�l���)0���y�^��Xjűg�~0��:P+S�+Ǟ�/~n����3:9fެN��!L��L�m�������S������;$�0�-�n� :<p���`jЂ�ٳ�y�4j��U��u����H'QP���E�ë�S��ГӁErbzѰ搞��t���P�s�A��|��x�����&�����r+x&��ڎ�Gx$�XN�`^V�����^�d*s=���/�f�l}$��D���.����,�1G�k�hr�6up��Z4�C���J5C�����I�0Q���� \�ȳ�+�M�Ņ��a�2���2��Of�WQ� gpN\���c��2C�VU����Vx��XD*�!H�8	���
S5��\v�$Z��X���۫\E�[#a�?�M�[���gt�/�9�y����������<�뻯������"T&ᒶ&�E �-N���ĹK>;�7"[O�7��c�=��"�_</��l�����{�\�����K���˗�R��7��WG��{ovl�,�\�]��3Ү)|P0KC[*��;���on^8�hZ:o;8j�r����(�<h�*�)1�6e�塕��jl\~�B�2p�%x�r�
�t86�x�P�������7��oY�|Ž�{�.�+��3:Ϟ��Y����AC�2\����;�(�s��[�B��Q�@e^�X��M�:�4�n�#l��)�0���C�jB�B+�!i��g�1�әց���R�P-W��i���7ba���$�m��p���R��r?�չXcr��96���N�" ���'4�U[�� j�G* �yb����C  ����9s�2�EaL!0s����h��+���cr(x���~��/���/�`���/���K޺S�wޣ�ݴ�s�R�G�@�+��'5��W� <l�Y���|��ބ��oL?�e�Y�==ge�GO�XM���&����i|�?3~޺�����^zר��|�e_�������=�s�S��Mkn:p���D��ð��
�-�l��ʳ;{>620�������!�Q����i����g���	�Lau� ��$oG��z_�>�EE�r����Y�ӳ�S_�⿯;y��_����>�uxF�mܛ��w2Z5&qSE"��@^��Z2k��h����!SR(ŗ�ͨ*ahm��O_�ީ�%x�`tc��.�=���>,�fO!������*�C<��S�S.���"iL�yN4�����pɛ��:D+�ak�a�3��peT����o����|��B�t�:��qH�)�������̙�0����kY�x�" !O�Ǚ2��y�)re����K�;����/����^�e���W�����&Չ5AlW�J��
�խ�����G���w���?V�}a�����R�O���f�H��%�r#oܴ9{���}��s��o�⥿kx�������ǯ�?�Y���;�\Ȟ�U
�Z}3ҞJb��ò�c����l���"47�Ȅrv�f�� E�K��12��Q����uzf�>�X�3�N9X=ǯs���������^}�78��Sr�Yg>�j�Cfxt�/�Prp� ��Y����*�P|���C	�T��zC�	����	�4�l�#�ܦ-�N'�z�zߋ
uV���>���$���-m�R�_+�=���r8K���q5QS�t�zz9W$�$�r�@��~�#���7\!��pJ�0�+B4���J�����Qɛ�[.��(
���n,����f),��C�wY뷑���wl;b[�G`��?���-�y����Re�fR(���k�So�_��?��Ǿ���ܯ�����ٻ�m�����٘�6�L�J�����o۵o����Ƨ�uǂ�)�Z���9z7�p`������\�rjGW��y;;�9z����%!l,a^}���*�f�=ö��/��^���Eэ
� �#�-y=�XjcWm>��7?�ЃO���{n{���^�u�F����$���d|�ؐ��74�!�1;���2jc�T
qgy,*
F	�nsU�b�B;�|�����j�h� r�+{~�y^kz��@`�=6���H<B�x�x1�OM��xf��,yP
�k(������O�s�pD�t2��1:8�C�d�*��T��,�P(R�,C���0� ���K�<V�����h�����7>�a��p�@D�䍉�Bc�4��[:ͩ�@z�ȎYSh�תU�����~Su����+�1Etb�.6���c6�qc��w���/�׾���˃߽��o���3q��Y��S����U�"�̒1�O�����N=��٧�� -X@æ��p�{޾���g���p2ͩ��atP�2��,,0�1زu���<-*��5~�aѢ��E+u�`}HYP*���T!������ӗ~��'�<��N[�Dgg���:O��H@C�܀s+j�Q.�����	��0:�ej�b�����"�044�!�yq��K$�7#y5*j>�S��"�)hČ�̵�����ܓ]�b�������7Uᤓ� �>� ��؇?|1ޔ(�r�-�����[�o�9+/z�;��!�D:�b��a�f�p�y�@"%H!��
���w��T���	�D<.zHT'=W@���:ω/&.�qb�<C��5h��4o8�G��b5\�Ĕ�'/N�D�<R7���k`��7};_�͏j��
Jܬ���v(��}�Q���o����<��%�}�o�\���I��Ձ�Zm���y���szz�����?|�E�OZ��� n�<��c[��\_�E׏��E@49Am2�0A�X��c������v�	�p�^S��bЃ'�1\�j5y=�ۙ&��	N�f@��F4�w�u���֮{l��7�p��z�)�T�X�at6�!ƅ�U��7����pj>��iSє���M��hhQ0-�j�&/����j�O��Q�ŉD����S���'�Ę%�0}B��*!N��z�HLc�n��Ê�3S��Tv��4_���w��\�5���'{��d�5����%p����߷J�,s�BY��,x��� o�^�z�iлt6<���L�C�5�m��@K:�Z��{�V��A?Hs�R!2<��ohl�Ss�%q>���674�K�[-GC�쑼�~��{���/�+�k��%�Dlhdx��z�?�H���s͚�;���}{v�w�81o٢c�oX�Ne&g�ݵ{�}���k���;�:�+�Z5�r�iD�n��a��KV<YaRZh�w�NaRЭ��Q�N氝�
U�$�h�:U�4�BFJ��V=���e�%KI؆PE���H��}���v����k����SN:��%K��E��^�at9p�
�b���s�I�|6�r� !*�;U���n.��6Q�+�Qy>�4�&SLK����WI��jA�p�>�P�Q	m���"�<C$���� ,�7�{ѻy��������5RQ��Щt_������09��W��T�"���n���
����\Ő�>f��{�� ��(5���ڔ��xRS���BH
e�Kye<���Qw'��x��ʀOs�!yCoS�ND�!��2�&��Xp�W������H	�/���lnL&�]x�/�^ؿ?�f�M�=��g�m������ˏ]'�p"��hٻs�'z��������>��ￛ�.�ܾ�h;��T�K"�@�j��8�J�� ����)�hh�����)�? ػ�ɤ�GS&�|�+��FBq;ʪr����95qP�i||��L&s���On��5��t�i��r�ҥ98�Ѝΰ|?nR� _�K��c�F#5�X[?xfC&s8�,���c������

9�$Q%�&$�sڬ�y"l��1��H$��,?�� �������5c.RB���ϼ {�leɬŋ��oX[�Z�����jn����p45v������p�3�F�!�q�`�g����.����� d˓09��� 3;��ꮫ�Mtx2�< A��u�.NbS,@GG;䨬���B	�Y���ۚ N�{G�w�6^'�kҤD7О�;0o��c]S8����36��g���)���$�8aHx��U�?=t���m��'��|��s�̘?�(f�<~������}����w�e#����#~�0!��a�(ZZ��Q�Q�� 
R��B���{�ٰ������<5Q��ѿ	O�s�`n��A�k���4|���˞~����ٻ������~�lɒ��S�E��C7��"KEL��J����NI-�7M�b(<=<峬r�s(%��Q�w�a�Fa�$ǅ�=����3��M��@2>�ʘG!#Ug�bL$S���Ή�S\!�Dt8�ē��?����x�>8u��0��w��wp֛V�j�p`�n�b3a�����'������gp���x�lشw �}�i��QX�xLf���p�o�=��b�����Fz@����fm��c7����{�4y�2س�f���I��ɦ&�QhCW$�yC+����"ɾҎ���mM����<��eF�G�qÌ�G���-�G�%�x�/oyۦ'�.�͝1��K�;w6�����qi�4O�B������T��W�@�y^3�a1]�@�Զp��^��>��kO�a���� ��D�A�}���q�H��z�Jp*;�brjrŖ�~꫗����3�x�٫V�~9��0�K��H:�)�SYD�2��H�4��S]�kP-�����I��/�aI�CAP#,B!����=Gm�1����1�T�ͦѩ��nmM|*�-.g�пg,�5津Ѐsp�u?�����������vX�h	��*���렧o
�[-�m�i�ÚatpûX�y���faN��p����I��R`�*�W<D�jS�6M!`n�<�J�H�14���S`�a�{���F*���94
+�JS$�Bp|WUB/+�{�e���o�|np�G���T�(�\���?~�������Sc��h�k=7:v��Q0�3(�T�p�����j$� ?n��`�֪�P����f}����XC�F�(�
���]���(�۷0��V����7�;�YkC�� �����_���|���s���v�����ù�xf�&A�N���Q�Vb�5��	}T�]�kB����C�rV
9�|E0��B���Έ8��%��E�8�Qk8��IΉhĦ:p>�rS�tV��f!��ixj�c`b�ɂ\�64�.�����	�YBT�W���94�
��J��trYvC�1ƪ:�x�ǉ7�1L�E� �<M���kB)��8����3�9Œc�3�<v������v������`X(��T3���#�F7�?{�\B�tQ%���5O=����U�x� >����i����j���s�AC�Lذi3��^����Gvl2G	�Ey������ֵ���"��������g�\��\�ϝ5̝+���y�G`xx��/
U�#��f{�XC�T*�+
_��p�׿q��7���7���C
;��d�[Y�J"5*E�"��qNc�.���WH}��1�RT�Ąח��ˍM�4΁���������5c6���	ӘJ�i	l� ��O!};���
T����NN��&��|��s�
�&)�yq]a�%)i�Ѯ�;���h�T"�y��P���:z���V48=�@ĴDh�U����f&H�+D�-D!��������R���I�#�~םFi)& �<��1DM">K��L=�L'�j�2�G��2����6�o��-p0쥭��7�:�Kq����/�t���o���^;5Q\�}Լ��->88:&
grM^��F�8�Kk���ڤ�x>������i=��`�h�y8�l��H��a�h�Qt$�":H���(E��2�/�����;YsA^�o��/�����������p�)�����é^���T&���I�NѸ���B��������Сs�qgT}0]��]4dVh�*���3�en�Ľ828� g�7]��E=CC5]Fz8��UVd��i�	<\E����ٝQ".�%�I6>�^��3��h�
�.�g�PM�.�U�0�5��FbQ��8ѹ ؼ��%��2�R�ykZQ#�d:��MP ��7Y�=>0(Ĕ��M��
�y|���ԭd4|D��46��Rf�"ٯ�5-A2��d4�93��W��h�|׻���Y�������N�s`�qw�ySyH�V�a�ԧ4h�
PP�{��^���?���A��@_?���PL�������i1(�l�٫kXN�R�K!,�2R��s�?�Ys;QD\��}�C6:I�յ{$M�����â���A7��Tt��hYr$�s�|���/�-DS-�������ԁW�3E!���*��t=%�z6IDU�k�f���9��)��3ЦU�8��h��=2ʒ0�k8�WAB\�t������o���~b����hL���.O,gK<�@�p�ރ��d5��A:t1�@-�	q�]�R~a¦�$l�ʦ���xؔ��H����0.�Mj�WvcSG�Q��ȯ/��z���f*�O�R�����r	��Z|!S�}��k��^���ۛ(p$qfЖD�R���L�GUMʓ�A��!#��<h�1���h�Ȫ�"�b��p�Ϳ��v6T	�B���Vִ�chb��[��0�H�������Kr�K}��<����Ț9C��X�A�e����v(�bՁ�V�XY�oE�1H����Q�����y�I�r��u���|/;߫�#�x+=���&xR�SDc�Y���`(@=���!#���I!o(��t$+E��p�fԆУC3��x7XTB�50څ������#�iU4N�|h(r$��|C�r-��X{�̌��ג,�`|>wR"�O�,Cw"�B�8�V�g���#����}Uf`�fv/H����ٶ
�!�>?�ï�Z���'��W������� ��$t(�	j���H����Lz+���D��+������^����hoo�p_r�L!�ܰ;v��;vA"�´	=W��A��5�ni:jaO��@tT<���n{K��K}��3:+> J� ��� 4
z����*�J�DZZ�c�(N�QS
�h�P�;�!f��6";Ѵ�$��%}H�b@zo���2a�$�F�q����>�s#
���J�����$��	�O��A��KEϖ�$0)��F�7��ۙl��Y���:�h�m��GTWE�I�{���>�I&JjB�T��G6$�B�9j������$Mj�����c(#�x�r�]�܆ L�s�i�_�N3��//*m�\�-�X�P��m�tB`E`�^���V<\��QM{U9�B%CۛB�h4�ך<�������{vs��?�[����h�}��1�s8����0/�xn����3:[q���6 �:���2�fl��{���3�����j�'a���i��K�e^���A$~d�J�jD�p����+xU�hӫ)�55&�P�O`�E�!:̞�c�CP)�w{b���ߨ�I�:�u�m�W��Q5*�{)|� �d,!6�:�\��	u��pcXp���5��(iMì��f����do�HL!G���TlI	���;�`(Q@���� ��h�,9�VF�j��(h�E<�&�����	���n�+4�5CR�)�ILk�!A~��[��^�"Nɱ?��2sj��k2햲`+�Fo^Ι08:*�s^#��w~\��j�_�Q�Tﭽ��,�!�*�39G���@�t ��Ц6R�����u�w@3&g�c���������߱�~�\5yE���$Ϩ�N޶>�qPu� w+M�P��9L"l45�_�wxF�he<z2�b�M�K�Y�&㖔�J.�×�"ZnO�N0�Li���H��g�*~H��B9~�BG��+�����)�����Q��"�&��̥�;��b�b��懆a�닪#�ɩh� �.����%�fb�OD%Z���/:�x�;}��+g|#4�&g�֕�ԁ�`�X%�})���%�.�C��ŃG`�"\ע<;pX�.����5��ͱ��~�}�:vIyr
�)�M:�����0���Аj��c�K<�����j]셼�F�rd�1�W'�s���`BH���!'1�l?q�!Ź]%��
�##p�1����~7���[�(�K��������'��ZXo��[�S��/������@�D#vCC�KB������
�V�p/�V�)h/��.��&�`<���-��W}�G{�Dˈ.��7�X1�I<��'�����W�b	�H�2ga���|��R��"y���,1�(�x��`���5���3�!��&���i`[���O����� K1=Z�؏a8[�����8��WM� W�e����hC<BP�s��$	]%x��ʱ�����=�}�2��4���e<5���n
%�_0%(c�T����Χ�U^S���Z=�����#:��A�&I(A�|!	��
 ]�Ṫ����F(#���!�N�>��)�PuSb��`��K�q���A�s|0]!���օE�n&���K}�ä�k�>�"�8I�cU���r�U��AO�@�(��B��V	�|=AC�2�⎫��إ*�{�	��R��S��]���a6Tj��0�|�P����Qj���� l����DϗH�
++F��9Mo������"'6Ĵ�Ղ�FOOO���}9�xd�.����`��	��7�Em
�|�[0^[�k�"�U-�Z �y��4��Y�X�yȏ��`h2ڀ��}=c0��@���M�
��~��O:��jm�x`||�4���`H����I��N���^1�/����Cg.UQĢ��������~頣I�3�c�k��N�̙],C�p��c�VP%�1�� -�t :�b/I�SR�D���[[ۆ��p�>�a�^�>3��a�i@A1 ��L�tJ� ��:�/t���Y����FF1aG��\�t�&��"�ۦ��4taMGt�V�DX�j?x��f��Z*��z'��^�`�R+�
&."v��7�@�rr�or��>�����f�v���Wct�� a���Q��/n`Pc�����P�Z�,M?P��f�����D:�̡ޟ`�j���R&��ńQȀ�EoKscJ����J� ҍm��#p ��|��֎�ᯰV�����s�G�m���;v3�
�}�U�x���4�$����$����Us'1�"$P�Ҝ%1A�Р7lz�Z|,�SIX�x1W"��K�I�=��Q����_tо��"�(2�Ɔ�=g�}v�>��]KK���r[&]�Xc�0�on�#h�3U6�K�܉E� �/��<O��<2z���^���ѕ\0��qhH��$(�Dsɢ�>�x�;2 p��8��0N�jj��%���T��G�7�2LH Z��xզK�t�xN*�!Y&��E�2+��^,zYGJ0B�Sk���N¤�>	/��1C�{�@�`�[
�a�g[�O�B�)Ij=�s����<�۳���3�,\	��)�rP�ၖ�C��9��{��P�(TKƦ�b18��^����m?�·�U���:��s)���{�g�����C���`座�_C�(���k���0-1P4��y��d�Y����&�)���o~�;p�ʕZ.`��j�R3U�oLag=j����o�4%�p:;;�fޣ���a�dG�?�xΛBZ8��6��	��������`#x��rS�R�����ݷ&�{1�3�Ei���JB��!憑4�F�D��9|���KI^(�,�pћ�D~~/D�[4\�KD��)h�v+�kA{^_R�xbMC�|�>�${��4X`�4��p/��'��*����$W]��&^Fτ6蓴�rD�\|q�iŬ��n(��$;�]��PW)��e�d���c���Ja� 2�����3-ǚ�Ѵ��1�ۦζ)-�U$)c
����C)�!P���?�1�~ѳ��r�a���bކPU���l#E��3��
���Md`�d@��y�_y�|�����������g��O<q������ht��A���W�s�b��`w�W��(q�H�V*�̙�D�E;����*�`��Z��>�8466��E��9�������-/�v�>�w�l�P>�a����=���'җ�S���Dr�J�W��߻X��[-��KfФ���:�h��K�ZÍ0B�08��m��X�+���X�B���N"��`[�3�Vá��bI5�W�XA�#xةD��6�ʞ�g( l/;E����
}ɖ�K�Qb��T��p����M�縉C5z�������V%U�$|_&���<��U�{�/�xt���x������������|�C���X�y��eOU���@s|?����r�G�x�~8�_\jJz_�~l��ʎ�n��Q���r~\2J�P�1WƜFN�u������I-����	�3y�[ڞ�7�� Mo���:�\����~��;�n�zq__�{0T?�h7����t#G-tX�h�=�̙3Y���۳�E(�B>��E��%h�����Q���k��hG<�ִ�T���5z�ѓ4��͛wH��a]�������O;��L�D5��b⟃d��V�Y-�G�~bs�O�ɅD:�M����Ӡ��+��K�΃'7�綏C,��]���!O?.5��|�����{ I�k�����h�7[R�G���)'��,d�3��Р�a.g���*:cȥ����C�X��'��s���{���O��kt}�C�i�|�ڵk�^�y�������V�(qhG�]�0r��i��u�&�ld������)�1��g9�����HG����¿�fi��s��ޟ.���0�P�Q(���C�^~Y��
D�F�c�0��h�#$�T�`4WY�Pʦƞr�1��ΰZ��MG�q,o���04��]{F��ZEMK{����w�����'����Ύ��eQ-x�k�Ν��j2�5o@ԏCȋCq؂��a�L������0��1<JКgL(��w���[�u��g��`�w˓O>�^��.�C�er�7p�%	$Q/R1�jb���0���<�������ox
�{v`+��q��Anߪ���Dym�H��S��C�R*���͵�6�rF'Ǣ[�lyʵ�6����q�46�����͚3l���m5h�D9WyC��3
4�!d�A
yp�q�mF���k�n���78OS��%�����lm��gΚ��D*�m���I4#X�,	YEt7���}��� z�XH:5pSP�-�A��$R�d[�W|�﯅��U��~p�}��tp��{{��13>��j௬K��'!_���6
�$�0�MG㬉@-�r� Sx ��y��#�\ҊT16"�)M��Ȅ���a�:_�hi8�����C�/�����Hz�a8m�x�q�@�zo(Z�V'W:ZUӏ�����X�XS���IE9��<�x$C��,	τ��طg�-�mګ��o���������O��iVc�%���w�����T�&����uK�8����T�e��
��ht�M0lW�wj��%�yɉ����-܋�9�C����w&�>��Ϭ�xe&�ӋS��Ţ ����b̉J��J�̬s�Ȼ�����͛ٛ��;�'�+U&5��*�6JL.c~!�F�����&��#�H���s�P���2:���0~]��'�N��Z!Ɋ�&D@�!Ƿ�N�Yߏ�UʕǛ'�_
�Rz~���@}�z�5���ẃ�ˏ{���w�ў��Tθ�G�߳���W_N�N�?�������i�Yl*�`dds��*�4v �B����&Ѩ����n�r\�l鎙�kt��B��\'��mn���O��g�:Z��vAij���Z����}�|R�/�8�#@M�x��˾�=p��w����܆����˖,�?��N6>B?�!Q�I^̪�+���ػ�.��єFg׌�\p�!�\^��ъ���*��%SYsQ�A�x(��T�-Cc)v��4>����Q~�P�F{�3:R�d$%���H�@|@�Ө9:&�x��NjXzܬս���`I��07��ߺ~^���k?��q��Z�B�7���`AHr�r�1(g�@!M���ULf?A3�!�E2�0�?t]Z��k���
���[`�.�AXM=���r�5w?����TOQ,��T��hJ�F���l�L�a�u��j<��1x�o�z�044�a%y-&>6�Mډ�?M�@FW���k�[�ϝ;R�$�����{}�F'%:2�}=ߖ,�&�ē � F��<$ڛ������{��??��kՌY�����x�B �<��P2L��F ݉&���p��K�6:\��1��(<8�u�ʛ�����p�#��|�kz�ј�����Ƅ��)U�����γ�p�2��0�D5H��3]� ��P�#?Y��Ȏ�@vT�����^���<l�遊�!Q4���n��YW����l���26?uJ��}�(f2Q�A��B�� ��f����x&�H��+��1�ңzRᮻ�$F�x�'
(�c.�A^*���+����\�lkk��쐁/��h5�S(L��
r։6�H$1�I��/�F�M҅�z`���0}�m�-f^ط�%?������\	��o���$�<�! UzR4%�Z9�ÜTD�մ̮�˪%��٩��Yg^�%���Ⱥ�mS�c��˯��O�Wc�y忶���q���0�ԏ���9��:�jzN���A#�J`c�ȕ3�d�׀ �$Q���FR�`b<S%��0��߉FR�I �dq��c8�_�C7^��������.Z���^w�$�W�{��ف��O��OeƦi�Ix�������r˥�{��֕˟�ӓ��f�4kΜ�@��;v�b�bAST�Ԛ^F2��4��{cA%�ǅH�&e��fs��!�EF'������/�U�N��������BCш�Ʋa��o{v�,57V��Ρ��3� �]����HB}�pS��6S�qe�C"	�1�8����I	�[�3.H�����e?�W��˻O;��;�%g�Q�T��x�
2N�-!���;�4�[7�^v�v*豐&�S4�K-��4?UfG#Ҭ�3B��
�B�p�D��@!I媋Fc�~:��M k��DA�b$�������,@1[���<TX8Cr-��րt��Q�q��ݟ�BƱ0�A��eZ�7�xt�o`���z\徾��X�MC���#C��V������3ϼ�5k�w?���l�/[.��K����$Yok<��w���B��u��i̮��Lp��?��+�� t�	�3���l�q�|xY_����{��qʥ�O�P��$H)L`yG�yK�n��]oڿS2�q��9'��𧵳�f&��X�Ǉaj$�i�Y�U(�Ғ4BTD�܏�J ^X��Iߏ�Y��G;�w��1&����ﺣ�{��G�.Y�����x�[�}��+�C��x�񐁊�9K�=P�GV�hH�oE�QU��T]N��'*^B���^41`U%�svJ1�U����3�y����ZT;��_��1%E9W��DJhlf��硛����K8U}�B��b��f�P���F�74ܞn���������6 �;��G��׿���^ȕʐ/�Hlϵ�ϟ��?�����]q��5y��+�l��7 .<�P(_*�q�fքL�	_g����t@0^�P�e&`Μ�eMr��/6:ZR8|��݊�&�d�)I�PQI��<����G/*�sKő���w=�6k����L�o��.XhhIh�<�
�օQȗ*�����hn���h�IJĄ���c	�@�I,a��G���=�V�Z��]Ɯ�1����N1��qy�5���Rm���)t��~W�W�C	��L�⋡\"Z���	�A�I�}1wG�Y�$P\B�+`�,�q3ʘ��PȖ�4�D�C���$TY[=j�5��9�1�>C�Q.T��G��i�d��ni�*u��k����C*_�-�`h_�ܖ9�wzo�>68�Y�����Zn:�3��o��>�W��q��_��羴.j;Y��N46&��˘��Tx�Ȉ�c�q#O�r2����?d��#bt��3G�>arY{.���:�'^*L\U8�#�߷~�����4�u�-�Q�j�A��C��&����x��2KSP��u����4z�]��9�ѫɡוU�7�V3��Y5���ż�tJ�=��I�K�9� ^dC
C���e�z����&�ԸI�^ȧ��ðT�f��E�:V*$@F� ;g�#�?�0�&I$��P���%��T$��Kx�d&a<_ _�L��DJ����4�~�������
v��ݜ�ٹ���FF2L�1��q^,��C��9�ʚ���j
���Y��O�7>�����gp��F&�`,��њ�H�Y�}���T��&3S���!�/G��h�g��_ٳ�{����Z�!D� 1�(�8�6t�@A��)w��붤�l޸��W[�:�W�f�0+�]��+Ƅ�*�*	�5�1�4��f�4���Q"<2�d�u4f�#���8��7RM��Yc�#��t�4\�c�!�Z3L2B�` n��(��<b��Ő*�7���eK�2��e�⎃y?ۆ��OE402��!o)���2DY���r�D�0��̧��=�jdd &�$/���$k�Q�A�V�d*����3~��o���
w�c�^���?c���M�;xa�P��h友�:������
N���ӟ�}����\�]���K�I��L��mW���J&6�~��������$$��#ft����M��ٳ*�0���*�➭���A\��%,8=zJ�s�v��o��M��}�]3�c�Y������T�%�ј�H����(�7+z�"L��D��g =��âD���LA#@��r]�ί��@���xA&y5�6��;�B�����J�A
B��0O`,riU��V.��*����ި`0�
�Ê�CDN� �â��r �^4���ΔE��y����	����p����Jpu��ԱP4������_��[���2�l�����oM�EG`>5	���ޅ�a�z�W�-M�����/s��?�y��z�7���plt�ݸMV��k��C�@I���������r�W|��Z1G����J0:��ܨ�z�<r6:I^5����y��4Ks8'���qϮo�����.�8o��[���;Y>f�����o��9�htYg�'[Dn�=`��-�.f��������B�,��T�Pi`1�L��J��`��lΚ��W2,1��p4�'�5��y��`X�;��bZ�4V'=������NTcplC$)&ީ*K��<��	;��B���~�z��brf*$���K�Dr�z��м����z[ל7^}�u��BI}�=��ѡ˦��djd��G'�`*_�F���E�B�j��M�o����E>��P~v�}��w���g���w��gc.�-��ܹ�}�;��z���9�FGK�����>/e�n�RY��n*�Q��6D1�jU��yyB�����z6�*L�u�p�w'�w=>�zs��G������;v���pvGS���pJ��n��k����r[���#�c��!��UJB��I����h,�P`ZL�r��cH%��T �.
5�T��Y�C�[4w��BTj�		'1��c�ɋj!f!�<*� ��U��+�-&�e�,��9]@���b�'�����Ǣ�+����!���w���}^�+��N@����m�|�41>;�+��x'�-��p�Y��x�ro��SO�"f5|'e�_u��N�?ɶ-̤fl�ꗿ���>�7:Z�9svW���*;7K���ᖇ�T$��C@�irE1';6=���c�����{�{��?��������'�ŧ�b~ݺ��;crd������eן�
ǘ<��v���J���'��
�xH�4ϕ(H��!&��<�[�����2�ǯ[���S8�ؼ�YgF2����ߛV�!�R~�f��J#1��<X�ş
Q�d3g��,��xpX��E]����6�r�n��zr��O\��o������*�lm�Ƈ�07o����:�fG�'`t��E&�VP��?����ս�O=U�Wa}��n�/���s�"FG+�dަ����w�����n$pt���p��34R�6�e��߻��.�Uw��;�dH��NH^xg�i��P(�d|�x���䊾ɩ�(7bе0�f&"a�&�.K�Sۂ���NpH��teAG�F�a�GT��t��L��h�TH���F9t�s������W�DL�c��
��R�x��a�q0�#y��RLt�U|.�=��s�`���BOJHc��&�%٣��-�DjS<�Zw�o~���ׯ�o��G�K����?�����rɲ�SBC&��89��z��_�������K�W��h5,>jKv˶��jp]P%�5L��DE��_�Íۿ1	��lg{[�����{{����y�m�u��7>���h|4$H�_L<�xܶ�y����V��p<3�V��i&4E�*���"�DH�����>MC�B��缍h٨���r8��O�x��U���W� �m�<l�,T����е��Z�H�	05-?�H�So�f�4��RXÀ�*=�y;�Ɲ@���wu�w�[�x��O}�KGD�����m���l����������'+m�<ߵ��]´�lB�p��BfʀU}��U׿�[�{��h�������Kn�ڼ)����aI�>��(	R��a�t9BO���U`���ґ�􍟺lg�*'�U�����O�CjƏw�-�L�'��>o^!$y{}�O���
379)MNNƧ
�#_�ﻲo���{U�H�Ģ����H����<��~`���kC�t q�����3m�9����M�Y�x�$���Ƶj\�U�z�d�U�]6D��<z��+��֣�c�XoKG��3g�}���W0�T�|Ã&�-�Y9ڮ���R۲;l���nk��C�d���w#�"ry<G
�,��pW�p�H9Ɩ+׮}E�h_������N�>�e�sV�����aU�Z��$�����	P�i�b¸M�v�Bn�8j"?x`����ލ��Kn����jnx(7&WY��=O�]�4��]Q����\��?>"�����3ό�q9�yr+�R�cU����~�7��u���h�A=d�,��U��VXRM��;���9f޼�.���,��`�}�IOm�7�zՆ�v�]Ǟ���,|t�ֺ�����%HVV�f�!;�gQ�Ѹ2%�<��x S�I#�Xt�K�y���u�^��հ|�����`U��>LG�iY`ROC	=���F�m�ơ���Hgf��A��&ȎgW�O��O�e�<�z�fI�?��ъ��P�%��$�%�� *���kז�=�?��)�*:zI��}�"��U"�	麗hh�5E"�K���WM~��,
�������C�Kzqq׬De�K��1U�Ec9���?����9v*D�{b�f.RFEWwcQ��A#��G�j��H�����ʀ�^(93�g*�X�j��Uw߽^��U3:Z�'�+۷_2�3��\��hs����*p����O g�0"C��`pΥF�Lh���
v��2Jf�Qq�90��p�dܟ+v�U�/p}�%G�^5���
�k�kb�C��ʚ]QC��6{��8V<�]���wE��1�y#��T�n<�u�-_�����#�	k��	��t2(�=�/:�_M h��ԇ��
�(h�O��.�2Ab�rE�M�D[o���гM��`J�{
�����k�Z��������-i�b*��pd��uc��O�#��{ժlH!K$n��ad�����b 5脛r@Oؠ6됰%h�Ѱ������B1_,�,��j��W6��ߺ�	e�ڳ�V����	�5k��ZB	̨j�1���H���EcIxv�Mg�HM���Ԣ�(��RS���>dn��������4-x�/�k�\�!'�'�}��@���q��w����X�Y  Ʀ��#e%�2�\�(�$�O���`��Ui�Ҷ����i{;,׻�p�۾���;��
����^u����e˞�/��🾕�&��K���v�XQhzc}=�rO��}0���AS#����9�-49����E��_dZ"W��ʓ��?nT��������K +.�U_��Pԕ��$%{ڶ�~���A�Z��φ=#��bԄ�(���eWjD+h�lF���ǝǜ4�;v��TӮo7��S�ĭż����e% ���G�#��U�U���,%"�NU/��$�c^�x���	+²���T�ځ")+��%����������(t������,�d
,|7+��g�ͩ���U�]o;��j?�k�&Y ^���]}�;��v?��'qG�JDc_�G�1�Z�\A���lS8��&��^�i`�b�؆&p0I�:��#�G@d#�0���m͸��c��{�N�8��L�.+���`d�����~6��Ԑ��<��@�
h���L_�{��+qS��s�YU�4>[�?1Dː��e�Ƿ�Ƙ�]U��		m�:�J��	����	8�'�"�E~-�Vm!b���0O?��(
�_�8�!DJ���US�=U�ld�-���Ʉj�F��R�n��I
+E�z�\��<=���l`
W&%R?�UYü����aMQ����K�/�~6�&K��aU_��`z��z�W���Z\u����ӈ_�}=�DT�?�
E��n�
��I�U�yij�<�i���S a����,��4���� @�%v=,�㤠���TP]U̻y0-�����P��e�2�����=�(���4|,��i��#C�< �'Y�>������<��;b�A<�`�
Z��
�/����������Fb��TM�j2P40kUf9�EE'D"e,���=[d�T�`c�H��c�w֙��i�8��h5��xO��_��*�Y÷�5��C�����U�T~-�ׄ��ׂ���O}�?�uҰ�V�����������Qf4�]�0Iu �j�	
��4�!8�r��+��Ԛ��/6z=v� ��X�0�R�_�i�%�1bůM��JVa�U��&!�%f쀵�Ew��C�h�/`�^�{hl�^��>1Ny��͵D������k�����U�ի�n���.D��`a�bd�!1.X��n��ƥ{fł%B����&���>�ç����}��jو	�37�t'���5y��y��s�@���q�r,���7|�t��c]w��k�g+�Fz�ds"
��#�sX��e�!e/���!��V�.��� -h,#=�b�������)�G#����������/�|�5Z�&�aRb�@�xy�>���n�>�U_�w2�ΖY��.Լ������_%8l�9-���G	}F�A��rh�RB�����O>��Ź��R� a��a��E�G�|>ʁPa1-ba��Z�U�4Y���4f.��q3 ^�z�9'��ioc9iݰ�S3½���U�{V9xΈ�'�٤�uY�.A�H�1�T&[g�H�Z����jhg#B��,3�X?x��h�Et��'@N���A@�_�{BI���ɥ�,.����6�>:u�?��ZK1q������ůgΜ{0l��`>�T���:3;��@S5�k�$B�[�z4Y�;�"�	�L�&L}�0i�D'�4�t�����菇` ��E#3ؘ	8c.
�X�>7�Rr���Z)p�E�I���@�yP_@o׿[�:	����1�q��Rޥ�l$���D?	���V#Q,�fmPede�Y���!�pt��6�r>e18�:l3�Z��"�_2����o�B��B���D�d3w��pq���ܜI���Ăn��ߏ��h�|s���O���/���2��)�ݤҒ2A�r�Ԁ���^���#����:*����@';�Q�q��{3�")vN�c鎏:;g5��,S9hjŠ�nbY��M,��q��l��~٬L���"�ل	49�1s�(o�磐1��k�D��u�X1t1�1��Ճr�����h�F(�^M7���K�ĕ�KY���<�#T~/�U^�D��6���c��d=�[L<���γ��g��s+F�T��R�וL�ˋ�MT4tq�3�SIN���%oJ�k8���GgJ��'ed8DGm[��D�2Q>�]W<K�����xw_�v�F�.���2L�x�'��,��6�섽�ad̠�J����`��M�v���Y��I�f���z�+��?��0�z���m�p���
��Jv�&�M-���a427�t��|���̚;�\k�f@�d�9x��8�����ߧ��KZ�ou�bo��^����֝a=�2�L�(l�aS�T��e��<{2��1�9���\S��r)߅&�iq��Gԕ�iK3 ��'9���%�@�K2Qq�>�f���2(}�� 9�;LQ�|��l��qОc~ J�N׍��+u�ܨ���]X6�S�ʄ0=����{�UW{�Ԋ��Q�����g���7�$螌7B)�B{K�=��yޣ�Yv����j&�~��~'Q�)���5�C/�m�f��.����i��B���>��e�9sѰD�,"��OŢ˸H�����hPE�A�mju$7���f,W1Qɯ�P��jM�j�#��o��讶v@{�PW�a�b����`K������.�޽{pp~�%�1ѱ�A�t�=|�������'P�ܢh������r�.��Oz�-��"��):��y�Y8��`]V*s�MK!^ �tMU�<%"�[�YW;�qZ��hb���@�l����[D�~T9�q�� ���ud(���5��+�tda���h�����߁��@��nX���~t~vV�&�d��?�zc]׹!���8K��VK�p�\	��.���g'Z]��~�		��)*&��    IEND�B`�PK
     ˡ�Z��)��7  �7  /   images/544a1249-aa5b-4970-8b42-188baf88f36b.png�PNG

   IHDR   d   N   �ճ   	pHYs  �  ��+  7�IDATx��}��U��������^	!����(��T�cAt@�XpTPGAA��H'�$����o��^�^޷����O��98����{�=e������d��x_���}6�����[@�g�oy����}6�7	�������||UJE�D��@���" A`��y$I>���@`E�D'����\��"a�>��5 ,+\��AfH�� q�NA<��/Ӟ$�	���'��(�J�a��yv�6�ho���&z���T�V(���{o
��A\F�H�2��3L�?';Y�uoo��%�FG��Օ�d2�~������*���h��^T,~E&ѕH��mش����Kt�aӛE�_���|��	g�"� �D�QА?�2Mg�Z����{r��V���=��U�v�0�=��>,�����������	�����w}�|�o]ԫ��{����D.8�=�VA�,X�D�<�&�.���L7���� 
�ј��>�.*~dV��4Bٳ�>�=H0��r�f��Po���=t�tyG�a?�|���s^�	�DU�%���0�HInd�?��=�y�&��h(�:���y�Y�x�����9��_?������>,��p�����vZ3B�)�nE����2j:��p<��iT.�$�ɺ%E�p���"c�,q���k*�*�ɡ(��f������3���܋;��C2���0��hO'[��B@��:�<��m���gR���<��A�!i�u�v�:Ԕ�H����.� +<*�k �
����$�5Ҥ*M�gՅ�/���++���Gԫ>����oc"]��A���0	�S 3S��Pz|�d;DE���֧�"��u�����O�>��P���P�K"U��{�J�F����ۤת"�� K��'I�E��U�eڴ{��`jG�T����w���=��:J%4:팇 %�`�M�:��̫L/i������M�=-�I7���K���n��ShK_��k�RDSG��RR�'�[	!���`���,��YC�CdW<�W�W˔L���e{��]�N�jчe�c@~��t��H���~���rϽ~�pd��t�8H��@��@�@!Z�N��>}(߹��=N�J��
�:u1��s��d9KV�J�2��R�6Y��� 69N�\���b�H��WJ�L�T%�[!:(��Ո�������1 �9�,z�-��;��G��6R U�t+��I!�[^��$�Ey�*i�0��}*�=���I �h*JQ�#�t�m�rK^Y [�\jM�d8Y�B�:2��#	}��(�R:��ĩ�#I��Q/���U�>,�2<:@#U�Ha���A���r��H4N�(B4ED0�H��a���I ]�(��=HW�	/r� ��&;p�ski�R5M�GA�!�?�W�,;.b��5yPV���B6���*��C��̐�s؇d�;����_���g��(�A���*Ռ*E�>���D�4}��"#<G"?��q
���Y��� (
���` Pg[&�����-H����(�>�8  �U� �����9�gea_%����xǀ�X�6����k\�$Q4A04��D���[���-RԀB!� %�2%�*��T/C�U뀼����y��$s�lb%L>ě(C�yܬsO�*$�&@�0��mܳ�s�eY�He� uO���� +|ǚ�ib��Q� �U X�)����OqI��|r[�P�!(2ܶL��%x?Oq��h���0��Z����T� &�qs�>S��4�2��I� ^�8l!+��w����x�0��;wB���i��a��5yڲ���P�^����1蔣ک;��RM���`2lR�!
�E���$5�������&��YDP������2		�S4>��"q�@�d��\�3ܥ3�����_2��&*�I,�S/�S�*D���J���N�#M`�x-�BQ�֮+��Π��f� 9n�sn��p%W7���)=��4h��L#�J�Y�6싣�$�D�%�$�u�|�U���Cax�i�PJ�H�h<H�S��\��!Uէ�(� .!�*F��H��)�aa�EF@� ��ըR*Ü�hbp�\S���IDԓHˁA�S�<�`Ų�$�Ҵ ,Z�q\�zά��M9����_uHN0��ʂ�R�r�l͏Z�i���k��UHb���R�q
�L���5)�!Haܴ4$BF�J��s�C:������A��0�A�:��%�!�u�G�a�y��H�Z�U����g�}c���c����~����i��Кe���v"���DIRdR1�S�wS(אּz�%W'M��W�H���DU
%#�h��ʪ#�#^�Y����Ap����(����9B��8'Ddd��I��G�h����<�+���#��R*�ޗ t�»T�
�G~%)jI�2>K�Q���<W��Sץ�k��d��3K^�fr��$A�O��LSg%��Y�[!r7KAz�Ic)�X���	�L�l�Yf��-<#pRv�Q̦�IxY�=���߻���dED��7��39k���%��=�ühP��i{u(Ez�A�O��N��k��Hp�Ў9��4ߌ�K���l?��:}�<����&��
��­V�j�l��<"�xR7��nB��-k<`7�{���`rB��3°!�1�Lɺ,�H��A%H]`&��Uv����Q�
b��R��=��T L�r�eV��s3�\d8�P�i��g'�:�%��Ja�D���1�F�!����:$���d�}6e����@=�T��|I�Ș_�V�/�$��Ȍ3��3��U�G�UcmE�aQ~����o�a![LRe($�CQ�"�23��2\��>�K
�2��tx�:�%�M�0N�])@n���<��XH�{�?̦Ϟ�����0 b���R1��LI��4��PCQL�NCC�����n�]p�-�̠�1Øi�E0�>�Z*I�LВD <*�jT�T�OIw$��$^r)�����gJ$������6��Z�/�$s��Xe9�w .��`�p�N����uw�PK['�N����[�u26��j���-E50Lס�|����Q��ɨX�/��nhiIP\�҄��y�ީ 8�-NM]S)��u��.b�Y�K�$� -z� ��9a>����0���J��H��^�C��1�*��bN�C+��r���bf�E�l`U� �����XH5�"�t:��)���\�ӪU�ڮ��> C��X�
O�(ʏ����&`���0���Ie��D#��HC	c��s����kB��P[�F�ᜡH/�0јS��e�m0��@�r�t8� YH6!L�5�GT�Ë��w|�A�d&H�	�ܝ�Q�& %��1<��Q�P$������g+Su��`D��(�����⃦ba�Z^L�剘!+�T�R��Pb�{!@EY��<�.Qn�w��`f�c�eSO�)� 2��c.��U!2K$`5{��~�H)6V=�<�:�$��Xl�]bR��x�A���d2�(��cX�we:�Q*Z9����dW��g0��fQ:!�sT1�>��#\�:�_���5#EUϤ��A�IMb�ނ��b�,�,�����L���C��D�A0�W�K/a�,�V�PrE��2�R�Ñ �%2q 8��Q��n_��r��b�5-�"�D0K*T���D���+�|a	���dy�h�M�!'2���H�H���T*^J�fgǆ��C㙚��>�:���
�	�LAa%ڿ %�(�h�Y���;	�
4L6k�?86��xG�WM��{xed� �a%~�r����17�*J}@�� IP[LJ�z��O����P����=]�9I�ı�j�g�B �"�~ʪk�#`z�Q������>w���Ҋ��h��͘!BB��	�sϙ�2����J�o�I1!S+۰�ǩ��'�^l�&������ٖ�ˤ��&?�Z�A3�g-��Q�d"z]�^��
!p6��`Ci�$,��B�l���ۦQ�T���~q�y��O;��1���֋�`�`�Ejj
���(M�~ D�;��BUA%38 ޤ��:����X�U!�d	�J�xij75g�4��U��^�;����2i
�'�{8����$�-^!P�+
�
�
� ����8��c��cE�(�,�
��R-���k&��8��j�����C��;���t��a[
��z]���U���A򜽵?����L�j�ŷ]�"J	L����d�T�c��X�%�B H�ny�C�����V?#�F5	�Fp.I"�}d�MV�����L^`���-^<6L�I�t&.��p���ɤJ�?f6���)�Ao�cȎi��
UV���J0a.+m�hY�6�JP��M
�@��@@ٶ� TdH8o��k m��^	�Ҽ�b���~ʔV<V�a�il4�	v�A��Q7*|��>u�B�$ۭQ�(�*�ө�5�ӿ�uR����.o!5�}P������A^�!�u�� �|�*`E��m9������;b)�\��#� (
%E0��F���d(�+Qv�N�t�>yʑ�k�V��A۶�R_�@��9MM����M�����|�x�*�Xˏ%.3
t��%W^s��5��\}�W���Ƚ���IBl��~�u����g�A��w>mݺ��,��5^{c\�<���n��=u}���O>Iw�_3���7�x9ق�ao0�~9�51�6-�V�ZEst�n�i�=�Q[[+&��Sn2G3gΤ�a�T�4e�H�:��3���y>�����E��R�X&C7T��9�;�㻓��D�P\�t'|�E�]%�.f�������$�o�#mw�E�Ht:y�>������~y�mt��'��]G]���9_�T��k�i� �B04A��@�8��q����;�+��{����M7�����E_�*��O��D,L����M����9`e
p��BDM�g'�t<A��IjoNñ'0&e;A�ELnë��
v_�}���h�u� M��A�����SdG��D���&9�X��w�z�A�8������a��IϏ���4���P(�#�d|�������wk�����ߧ\K����i��5t�7�A�^t�t�0N�ओ�sk/�wX��|V�c�z�d���Ϝ������d&��އ�ڦ7V�[7�A_:�$:d�#�3_�������w��а2J r��� a��wXw����u[hdx�챐6o�Fkזy;P$�6�I#C��a�s���
�����M;it8ˋ�;vц[�� ���t�6mXŃ�L #ݲyqRf]'�_�Vx��|�lFd�A<�s�W�p�+�_��_�ze3]zǭ��dn���3��lٚ�+O�,�)��g�Be*xM����~���MAIըr������w�ɴ����O��w�S�p����K/��dN���ޡ�4!��(o^`{.o�qX�"�c��)�n���"�:��%�ĸ"c�Ƞ�\)�����b�?����_M�L{����KB�$ߣ1��B8�7<����4m�:���m@�%����F��AUY����̢u����]d9���o�㠊���r��[�ԉ�pxC��%Z$u�hք�a��[���kl�1���C��#R�,,��e����:�gʼ��=��k���[t���θ���}@��,�����a�����k6���Y�"�������jŢCٛאJ��֖f�~��0�,������}U���*�+���x����>���`�u	�,��;@���F��U��ǌo�A���O�����E���9���]Y������ޣ�:�5L�L>��x����.:� � �mklq��fHY�ɢ��ݎDe��$DŤoP�P9x��������%_x�G�����k_�o�t�{
O&?@�8zE[F<�c���`Er��0�2͙3���N� ;Ҹ_���Zy0LH�T:�՞�~�^�����6F�͙��g�9-d�:��*�����0^��c�,,�X������n�n��h�$W7)_�i�\��b�*̢(!�k�Y�WWB���L�iWh��$#P�B�U�@�\	&��u���*� L�+ʪ
�hث�����j�8�\e��LD�e�M#�������������=%v̱Ǿ�)��X�I!w�W�zu��PA^А�l7��M�϶e�sǶyB[{ 3���!K=`+s�q��a<lV�
ia��@5�W�B,���)=S�������yA����1a��6@2'.Y>M�XY�:^�&�`H|�+RhZ[��5kԊ�a{9aL(@C���ԁ�!���b2v�O�oJ�W��Ne��M_��uU��~��S�Y>D�@��Ǉ�Fo�6ޡ�sC�V�F���'	�uLN`�W����J	��_힯4�>� �����p4J�����\�@�I���q1 I
����ً��0yMT)���ջd)E�>�ϒ}x�hSs���E��!`}`���uK����98F�	��6L[�jBpۚb4�5F�1�-bv�J6D`"�жQQP��[w���(%]�ƫ#��1l[ ��;��e�!������x;xHr��C�H�L����o��;NO"K����O3f.0&I��%N�qk)���:?��7$>���yXa���(���x�A?e�3��Ȋ��,e'�T����%M�d/�{�gW���x��6��}��m<����,;E$�i���@a��P":�M��h���.�{1�'��1�6(������D�Oΐ��r�0g@��)	?cS�	����NS��UT5�K2+B�-��Ś�RcQ~�NE.0�����\r���/�z��=��|����?���#�����Ȭ�1	HO�o�t�18I� O�7�17F��7�������|KV�7�_.�m&������Fr��Qd�F5(#���F���f�{��]b�"�#&���Jf!��x^�eXݭ���Djw&]�>w֊n����}���A���=���=D��f��8&<�_�~��T��65��5����Ο����d[�
Ҿ)+���$JnO�#�v[���	����7D�.������l𝦩�i�W��L���_���u���.�c>�1��'�]`�4 PW��w
4r�L�b�=�5E����mJ�H(��������#�ks��`ˀ��*�,5J�W��UmYo7}򉗱��(�r�e��,0�?��]U�&� �c ����]�k��3��W���Oz8i�,}�ʯ�������o���b;����ڒ���{�ƹ_�������u�����dk�s�ZZ~��=���d9���|j�b-����K�d�B���LP�%��U��~(�
��,{����3W\u�+--�?<��G?�e�&sǎ-t�QG҉'|��X��.\�.�!ÈB���6BKG3eZS$k>��Fo�qQA�2^��ȼ�W��żkhkjN"+���Y�tttR�\�"p|ڴN�O�i�,��n���A*q�� ̂7��BY��߶e�ɯ�X�U|EI?������h�����'���#	��Iڷ�Ѯ����H����N���9�I��t�z�3ol���O��7�_��~�*A{�X�=lɜc���#��v=�t�,j��>��8�jbb�_M>{��)EY��e̲��+���OgΜ�Xg{{�Z�R8���=�{�b:ꨣ����ʇ�@L��X2La�5IJD�xJ�d؛��0R�#��!k�a�o�׷���AU�@�gϧ�؛^_�
͛=�|�Ɔi��t��P97F�l��{2��?D?��,ٌ���=;ojljȈxPa!޼���x(Bb,a��X�H]w�e�}珟�;��]|]��R� 胢�\�ֈEO�v9]��4�{�k�?��k_��7U/E��2R��/�����������=���Z"�T�C���+�@V�cV���d�V�S$ʶ�a��_�V9�Ы��7����6���W�}��⢽#�
}�?��/������sA5��:�-::��J�e�:B��QD�)�4����xrAh���7(��j���NC۶�THJ�4DN���*�}�Jz��J��	�a��R���9�s�$����m�����%��e)�T|$"�.pOiv���;ǜ6�����?���;��վ,��mߖHYr}�����)��M�=����m��ȇ.�E�f��i�l�RYy�5�\�Kr]c�� s��r�C@ر>�q���l$��099��!J�b�o�'��O�����N��L�_���G�Λ�/�p�ߥ+���tQ`+T֘\�U ��a�O�4N�(%(�*���zz8d17��_�B�@��<�~c�&�{�^.Ps*M�WN������ce�*��"��(�6�d��@�� ����a�##I�u��a�������^�������~��:��;���<7WѢV�i���>߫��{|�����߲�wӦM�-��^��O�ӱﻁtSDT}�e)�"��ķ��ݠ����Hi �?.��I���)Z��u*U*����|�.��/�>s�]�]�8�ύ��/�> l�(Y�Ca�[e+��DjB��"�f��0��ֻk�K`�s�&L�ܸ�W�5K;�e�u�7T�@� �>w�Y�8���C}�Ids�>/È����K�0��>�� <�HR�N�Y���Q/��ǘ\�{2'�(��������O����[�Ӛ�׈g��!ѯ\�Mz�{)$!�|��j���P�+�FT��$,HQl�0v��7��%���Cm�gv�Zե��Ҵ�nzy�5R@��ĮT�wC��
���ڹ��fΜu�y�_4����aܘ.�~}4YT"��Q�� �q
��Y^qcg�S��&ի��f��WJ5�ɻ��>t��y+����YB��H��tvL��	�8z 4��y|X��k�D`WLj#�j C*< ���Y�r�c���������$�:��|�跅��I`�d�qmo��$�p������.��x����-eW����Ul��2��o�[�,@XL�h�t�A�T"-"��_�E�L���1���vP.������H����N�y��+�m�2Ô����Sk�t`w��n��z��� S&��W�g��sf榒%�@
ʍ�5v SQ@�*kJk�fUZ6ض� 4�2���DN��!�.��y�7�	|���Sy���l�&<Ө���{�Z*�AZ�8j��$���u?)��8G��hxأ|(:�d�ò��7i�s��+�GԋI�D���ftYC�|V��̱�}&�������(��#�;�t �����!]f�~����X���b>������ag1�V|��Pr75�V�0% 3
#����8o^	�<Q�QB�HO��]�>D����S&W���^�����U��ƉV��rY����7�P`5-�b��kJ�j��Pd�ⓗ���G�~��R[��C�9#��:����	���t�C�����c��#O��h|����%�|�2�&cbb|1��㼷����E���5�W�Ej���~J��s�LJ57��X���dϮ�JJ�X��+�^/L��]�����&�5H��5Q������+-�~f~rv� �0AU���O&����1�C"~��$k�`�sY����wj��$�o����e�f�:�� )�euf�X���k���Qi֬7�@�����[�2���Q�~UC��Rϯ�Aad���ibw��f�&e���[B�Nj���	�;��1�{���ҥ���s���K���=l�1���3��U0�,XSF�^�_��oi�~K,�
6�Gn,��Xss,Dz������<������s�Q�$*��rj�����d�U���v�^�[���	(-��iښ�e=/>*ZE$�l�]#H8V_��Eꀥ�qܐ����0���<�u]�mR8.`JEf�� %�(H��w?tcv���x|����Db!�>��{����|il��a��۫T���5�T���*�_���r�Uߡ��422Z��&o]�p������7}.{LX��9���6�A���%[�i�@�L�y�Gb�a�+(\Xt��z�M����3��ik#�H�\��m��h,vP3m9�:��'bOym����[��.�\��Vz��ͥ���?M�����m���ui.s�Rc߄�QldT*�3Sa�D֗�Ϻs�W����J�lc�y+?�O�-z�ίQO&���C�xlO�7ζ�/�Y�̵U��T�uir� ]�FHМ��/?��O9����F��vǻ
�7�q5=����⋯�o��첿/����t�ݵm���@-���~�����I*�:-�?t���أ����0���$��p����q�N�:s��~�����rd��q��r+�qPj�<j�m�Qޖ}d�_z8ܬ~*>����&��pj��Wn�:T��_������1]��!����\��uR<������%��-����pbGXM�"�\��2mpijG�zZ"|UE4��<H��OiN��E��ӂ������h=oPy̥܎"�a�Cem��QE����/]���������3>���Χ�ڟ~�Û�K��m=���߾��C����i��(�R���8ψLS3��ey�KE�����j�G�%K�y����
�<��U��Ֆ��m{�zi��Wo�Nk���41��u�Գ��5�9p���s[W��h��=���z߽/�<�ƫ��'8���ᄬ���^Ir\U�EѰ@aQ�Ka�F��8`
��?մ���c6g	���X~��qwp�]1����J�Mԩ>a�	��h[}�]D����xK⸣���[�{���q�g����}�:�;�����C�~��L"?1I%1X�^Ӛk��')J���"��-��*�2���R��	����Hs�����BM�����9�3���v>R*n���͛W�i>A�a�1!s�eJBk�?y�4�d��T9�����r�6�f�rq0p�	Y�Gk5�*U%�Y�j�RdI�Q�)QE�t���RJt�6U����}��Xq'���iw*�b�uHm���I�Q�&GjT-3p�P�dc�L���	:�K�@������B�,_M���v�#q�b�=~}�ˎY���;�c��&Hk�:lٱ+֭�M��N���rEߏI{vT���X�ܸ8O~2g���a����}��Fmxށb�b&�)b����4���;�wl����9	ѫZTϖI
U�U0-	-єQ�rk/�}�%Lp�k�|���Rl~7p�H�X]H�mY<U�)NVf�P���d0�P���Iσ7����aQHj)A%����N}�FT�et��+����Y�A5x�{߃`#��4�����L�{,��ֵ��~s��H�X��c�+�|�ي�T&��y�q�����
�$E�3�˪&4���/�Ϝ1u������$qm�S�~Q�|�R+k�(���R�fВ�����]�R��ʚ�fD�HZ"�F�	�'O� /}
��=+�8 
;ê���#�����ƍ�Mw����F��g���O�*�B��A~"F� I����b�&����m
��oxp���>s��X$*5���O>��
Du�z���z�ە�B{�t��;�\s�k�V�z�&^�_���ܑG���ֿ���_��D1_�����w�m	��$��JQd����}����_�D��M�� i==�[��vY�^�Y�G�Ñ���#����}���ȏS��k�4�U>��Ƨ���)��x�v�\v\�a�ւ qH6|N��-+���۬��1m�+��c��o�-�� f�d�^�1ˠ�Y�D+���I��ݩ9��ϯZS9�ē�v4���R��w�����l����(��Q���Ln�@�/=F�O����_����/�:w����7V|�����:�k��/����ȑG�׾~5ɪJ{����}�?<}���9�۲������G|��+n���a@�M�B��^��:���}D���]'$F�wҼT�y�w��ɱ�]���3M��/��yp`�����H�<M�Ú����"�	��t:��Xi�(�4~�%��b;>�"��	����,�_�l��*� ����fOM�!�����x��O�`ك�tՏ����z��:� ��?9�ZC
�.�9U�nx޲֎A̜S�ZuY~���/�O��lU�ؾ~vl����{���d�7�eG��7W����g�fś3TC�nz�I�������w�}4	ȼ�R>_�^(�}���t�G��g�C��A�=�̻��TY���x;lߖ{�xk�>�^��h���:&�LG�\��Rv�����];'����_l�����D�U(*��4+�'D$�v�?h�	Lב��/f&_��47U��I�԰����L���ɯ���R��e��G�N_��6o�K/9���� m�����e�����]���S
���:mbA`UZ:��%:���iwP��o�8q�Pz�P�u
�=�W��>��b�T�;R(I�Y�8��g"_���59��'J�m3i{�z�sŊ?���O?������:JN�F��S����w?�������/��X4�
o G��PP���ܬ�s�R�Έ�5E�3�T���ӚF�N-o3j����yۿ�Xw������eG6� ���*vI��t����9��D�E)q<,�	�Z��s���[�<|���pX����t�.#Q��q�����	���*j�U Nl]��x�7*,q\,Mp��NLV��R4�$zv&hj���3z
�_ф�EOH�2�u�]�]$YY��6�B�6o(��.l�AA�S۲��+A#�}o��w��oѻ���֙}!(o��U�'�7��abݽ�7��Q+����h��:f��1߬X麱m�e��,�݁���n�b�v33V�.�|�y&�W��'*�hC|���J0���
��g���K�wO���ӒkDSYf%�K"��F����}�J�'.���꼘��q
Ą����	��q�@�k��Ȏ	!���VT(M��;g�U�A#A�� xe��U5�&j���u��Uc!��Gd����t�醧��z��K�g�ه��U�X~gHݯ:~�A�n��w�Y�HNx�� Z��GNă�~���ؾ�c��k �*9AM
�bu��J����$xv�Ei�-�����R*��`���1v�XյC�g��cɁ�I��6��+ϰ�� m&�m�{Wg_=����ߊ�
�*)��H�2֟�.�Al��;�:l	22;X7��Wo�7�3{Vi�[�{�2-��~�>�k���k�7�߰��/����R�꿌Opd���H6}Y���:�-ȒGb�]8_ Ae���MtTA�@u�۔b�+���6���P��$�Y�6s�^0����e��I`��e�������fp��.��nL]��J�]+����
�y��bBm�l���)`[�}��np公��HJN>��T�a�����H��Y��˗�_{�E��<�@���Ӕ	�d(�!���*ʃ����7|�W���9G]�Hg�`��EV��-���/�ī� _�]#
�]��b=Z���:u>>�`�[n\��.����(��؁	�M�G�tt���n[����L;��B��dtG�53~�m��9�p��$5c���6)���?<I���/��f}4�>�(Y�L]GK�O<fJ��lS\}��	=���ªz�e�h)�SR�a4����Q�P�1dEhv�2O�W9cY�v~� ��	$y|�\El��̂��8�W�[؀�5hf�s�[��W�,��:H&o�)Ӑ�T��oN��7�LVK��§��$�q�I��*����ϯz�Q����������W��MY���hR���aY|&,Kϴ����s���	I�XB��DR�PX-�#����|1z�x����6�V Y���@.ǰl�q��:R�R�Zv�jZ�����`6��9���+!����kW�Vֱͮ�;$J�����ۦQi�C{�v�_�������O����� ���    IEND�B`�PK
     ˡ�Z~��ٮ ٮ /   images/2cd57c9b-7217-4a6b-8577-1769ce4bee7a.png�PNG

   IHDR  �  �   V���   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���{���}��{.{�.�w � /�%�.֥����=�MF��m�D��Dr=�(M&��Ɍ�t���%�'Mc��i�ړFq'��Z��ʲ�X��\��@XX,���{���gA�@������3��9�=g��f�����Tօ�����رcxqqq�+W��v{K��n�;�d���v)ek���U��IRJ��j��ݖ$�$�$�מSJiUU5q��$�o��ճnb�[�>     XU���<w1I�&�M'Y��UU͔R:��<���;�B�u󥔹�������n����+������j����RJ��n_���Z8}���[�F  ��P� 6�{�wtӦMۖ���5���nwkUU�UUMTU����'���j<ɖR�����,Ϸ�%t      ��I�d�8)˅��R��$ӥ�K�Fc&�L)��R�L�څf�����ҫ����_|�Ź[   �
�p�=zt��h�-���ݥ�=UUmO�������mI�g���-��-7      �|�W��O�jo���Rʫ�F�|)�媪^Nr������3O=�ԥz#  �ڣ���<z��RʽUU��v��UU�/��$���N��w�Π      ���Or.�˽u.��R�骪^�v�/5������W���Z�  ��PpgC;r��Ϊ�&9��vUUu Ɂ$�z�{�4�K      l KY.��*�����dUU/$y���\��}����gk�   �B��u��Gm���N�`�C+��r0��$��      x�.�R�k4ϕR�O�\��J)O=s�ر+5�  ��B��u�]�z׶N�s���>���$�{�$#��      ��$'�<��٪��_J9������璔Z�  �mPpgMy�G�h4�f���H��'�So2      ��t1�����o���9v��L��   �F�X��j�>PU����zO�w'�?I��h       kY���L�?n4�M�V���ǎ;_w0   Ppg |�ck���G{��?��ILҨ7      ��q&��UU}����+W�|��矟�;   ��;�x��߽inn�ÍF�O�R>���$#5�      �5UU��R��7��4�ͯ;vl��P   �o
��������`UU)�|<ɿ�d��\       �eKI�SU�ד|maa�K�?����C  ��(��7G�9���I~,ɏD�      `=YJ�UU}���/?�䓏�  ��O����G�t:�f)�G��hUUԝ	      �U�L����h������?����u  `�Qp��j9r�CUU}����$��      @����-��N��������=v�ؕ�3  �6(�s'G��p�����;       �B�/v���}˖-������  �����[���,��ǥ��N���<       �9/%�'KKK��3�<s��0   w�L�ȑ#&ɧ��D�f�yx�v��$��*�V떯m4i6�     ��---�����5���)�$I:���I~mvv�7_|�Ź��   0ܹ�#G��L�W��L��5�YӚ�f��vZ��u�+��l^]�V+UU��n_-��Z�4�����f3�F���      ֖n�����$����n�>�t:)�\���:��յ��x��ʞܱ�I�Q����cǎ�Tw   ���u�=z(��%��������f�����gxx8CCC׭k���     ��k��ʕ\�r%W�_{maa!sss
�7w%�?-����O?�D�a   ���;I�x�UU��I��$ͺ��e��>::�������fdd��N�ݮ;&      ��u:����g~~�j�}~~>���������l��n�1��M�&�����o�  �ե��>|��V������$b�x�����x6m�t�v��>22Rw<      ��
�/_���Lfffr���6�ˍF��|��?�;   �C�}�:r���$=��%�9N_4��l޼9�7o�����5::Zw4      �;677w��>33����LOO���{7��ZU��xꩧN�  ��Rp�`}������ZJ��I���s�g�֭W�7o���X��_q      `�+�dvv�j�}zz:.\���B���f�|��j��ǎ�Rw   �C�w������h�Z�G���vTU����l߾=۷o��͛311Qw,      ��3??��/��W_����s���5?齔�tUU?;99�ם  ��O�}8|��v��_�R�J�f�ynW���֭[�cǎ�ܹ3[�nM���      ��---�9w�\���r�t�ݺc݉��I�󓓓��  �ݣ��9r�I��$���r;6oޜݻwgǎپ}�B;      @,..���󙚚�+���K�.��v���v�������    �
��Wu���O�R��$�ü����m۶�޽;{�����xݑ       6���ٜ={6���JΞ=�V�������������w�  �ۣ�:th����o�R�����J��Ȯ]�����޽;�����      6�N��W^y%�N�ʹs���^U��R�����Sug  ��)��3���#�F�w����,7RUUv�ؑ���g߾}J�       k@��ə3gr���LMM��Rw��y���{ꩧ�]w   �:r�ȑN�[I�ԝ�����s����w�}�;       whnn.�N�ʉ'277Ww����v?y���/�  �ۧ�N<���QUU��d�F��ܹ3�x�;�gϞ4���       p�t�ݼ���9q�DΝ;Ww��[J�s����]�A   �=
���<�ת����s���*�w��<��[��      �>�x�b�{:u*����\�oNNN�R�!   x��׸�G��t)�e �,�F8�w���;       �lvv6�<�L^x�t�ݺ�$I����SO=�w��  �[S{)�;w�ȑ�0�?NҨ3GUUٷo_�=�M�6�      �077��Ǐ��ɓ�0ѽ$������C�A   xs
�k�ѣG����I�u�عsg~��l޼��       ����<��9{�l�QJ�ONNN�Ӻ�   pk
�kБ#GL�I�ԕadd$=�P�瞺"       �F������������:c�%�ӓ��ߪ3   ����<��#�;��7��_��UU����y���j��       ��������<��s)�Ԓ���������g^�%    o�Yw nKc۶m�,���8|tt4�{��r�}���h�      �5��hd׮]ٵkWΟ?�N�SG�-�F�SSS�����=   ��྆=z�3I��:�>p�@����e||���      X'FGGs���ʕ+����#�;v��1?55��:  �֪���9r�p��&ٴ��6����@���<      ��ԩS��w������>�JUU�ꩧ���  pk&���;v��$���###��>��{���       l�7o�Ν;s���,..����$ڻw��|���Uo�  ps
�k��#G~6�Ϯ�����Ї>�����<      �ftt4����ٳgs�ʕ�<zo)efjj��y(   �V��[;z��D)��${V��͛7�~�244�ZG      ��u:�|��̅V��I���<���  ps��pk����U,�o۶-�Ї��      XU�v;���m۶�<vkUU{5  ��Lp`����j=�dt5Λ��ȇ?�����8       ޠ�����F���W��+KKK�<��3�W�@   n���j����R�}ll,����      �U���>��������I2�l6?�Z�  pk&��w��]�N&��Y�f3��G311��       �-����׿��,--��q�v��c�^Z��   �9������d��I�w�K�      ���y�����^��;��_^��   �9����}��䯬�Y̽�޻G      �m��{r����:�g<8�Z�  pc
��ԩS�v������������       �c=�P6mڴG�~l5  ��Zu��>�����{��޴Z�
���ŔR���v�YZZ��v����7��F:�N��      �E�ݾ����h4�l6SUUZ���ە�F��+�ԫ�l�=�yO��o���׳J)�L���   n��; �ۿ������I��y΁�����GlKKKYXX�������t��tn�x�����M��      ��X)��Z��Z��������q�����p��f��ƚ���~7'O���1W�\�����_��A   ܘ_50��R�Zno6�9z�h?�X�VJ�����t:������B:��u�W�      ַn��n���>9��l^-�gdd�����ѫE������̫{��G�����7�d�d��n�;I�I?  ���L)�~�q��ጌ�������t277��5??���i      l<KKKYZZ���|.]�t��VU�������^�}�j�۫�|p���Ù����9�F�(�  �F�}���~n�j�r���~Q�RJfgg333�˗/����������       o[)��{�7�j��+�oڴ)�6m���x������C���g���{���N�L�ԷC   �����u���?�h4���3���w桇����������W��+�����,-��      ����hddd$ccc����Zz���X�����?�>�l��������}   od�� i6�/��m���r��������\�|9/^̥K�2??����TU�f���_~��       ���fvv6���9w�\�d����v�I�������dbb"[�lɦM�����C���K?�_O�#I�  j��>@J)����v����h?�x[J)������tfff277�����Z����4�ʹZ�LLL$�I�       o���p����ǋ�����ʙ3g��t�j�2::�M�6e˖-ٲe�u�$���ٹsgΞ=��c>���  �9���h?7���{���m�t:y��Ws������d~~>�v;CCCi4i�Z�;&      ���h4�Ns_q�ҥLMM���ddd$���ٲeK�mۖv�]c��8p�����  ��)���nMr�_�7���ٳ�_ۿ%�N'�ϟ�Zh�r�J����n��.       �������BN�:�g�}6CCCW�۷o��=޽{���jeqq�_G�~衇�=��g�u    7��> ����T)�����w�^���+���W_͹s�2==���Ō����jehh(CCC��      ��w���+W�䥗^ʉ'�j�211�;vd۶m�������F#�v�ʙ3��/..�`����   ܐ���xw?7_���KKK9w�\.^�����4�]��v       �]�f3cccI�'�?���9~�x6mڔ�[�f��ݫ2�}Ϟ=}-�WU��(�  �:�QJyg?�߱cG���r�JΜ9�.daa!###W?�      ��m��K)���ʩS�2<<��[�f߾}}�t�;w�e�k��}|   nL�}p��ƣ����{�Rr�ܹ���+�������u��      ���h4��o<==��g�fhh(�v�ʞ={�h4��Y###����]��u��>>   7��>8����m���^�.]�K/�������4�lڴ��      ��PU��O�>{�lN�>�͛7g�޽����+gl۶M�  `�Qp����[�n}[__Jə3g��K/���fdd$���w)       �]�����p���O��hd���ٻw�ۚ�u�֜:u�.&�΁G}����w�u    o��> >�%�x����������/djj*CCC���       �hV�{���ʙ3g�cǎ8p �f������ߢ֥K�v'�[�  �7Rp �VkG?��ݏv[ZZʩS�r�����      �]WUU���s�ҥ|�;�ɮ]�r�=��V��v��]�Fc{�  V���`�[���lftt�-���ٳ9y�b;       �b��~���LMMe�޽ٷo�[�ڑ��4��,--�+^_�  �F
���hl�v�}�����gff��sϥ���      ����*�v;�Ν˹s�r�С�����׍������}ɴ����/  pS���t��m���ͦ��Rr�ĉ<��ө�*���       ԧ��TU��Ǐ�ĉ)�������w�E�  `�i3����������M�[XXȓO>������~E       ���j�2==������������~w)�o��  pc
����޼��6�l"����Odii)UU��x       �cUU������\�x�i�Z�<ߴ8  �U��>���~�����/����      �ni49y�dΝ;w����o�   �1�����n6��=>�|N�:ej;       kJUU9s�LΟ?��>wSp  Xe
�`�
����9}�t�{       �����>}:���W��~��]��  ��4�@)�o+?�/--��_��1       �j^x�,..&��w�  ���׹�i�N�J�ۭ9       �}���:u*��Tw   ��`ff溏g      ���ҥK�t�R�1   ���7�����#       �]w����#   p�)��s���~c      �uiff&�n��   �E
�����\�       �/J)����;   w���:���Pw       ���   ��unii��       �7�n��   �E
��\)��       �7�  X_�          
�           w           ��;           A�          ��Ъ;        � �:?��g�������d1I��\ZLJ�Hf6�������������  X��       n�������O���޷���RR�N�{��,]II�JJI��d��,5�n#�k$3�d��t������\�Z�\���ݿЋp9ɕ�<7�d�f�U��  �;       @͚I�)z��Z¼�^A1ɥ��Y.����-$��k%��Y.�_�k���k3�u���T�i�  �Ƣ�       ��j%�ֻ�����I^�ke�W�Y�s�Bu���  ��Qp       `P�$�w���	��|{)ח�_�.\��Z.�  �@�       �����I�w4m��q*�J�u>ɹ�z�J.���  ��(�       ���L���i�e���$gr}������*��K� `MRp       ����[oII.�7>�M�?��޵ӽ�3��y  XW�       `pL�֡7{aI����Sᯝ�r��*�د�  p7)�       ��4�d_o=|��d:�M�w���:��d���d��� ��(�       ������Ջ�����I������rY  �B�        X���n:�$Sym���$'z���:S%K�
 ����        ܎��7y�S�sym����L��dv5� ��(�        wS;ɾ�z��w�r����6�}e�3INTIgU� 0p�       ���HrOo}�F/���������U�	 @�       �A�2�J�j�X|_Y�UIY��  �}
�        �Z�-ɣ��z�%y&��I�J�d�v�J.�^D  ;        �^lN�z�:�L~�~�c���J�V3$  7��        l7���)�����l�?���W7"  
�        �F�Nr�������������W���	 �Q(�        �ض$魫�)�?����\%�V=! �:��        p{nT|/%9�������U2�� �&w        ���Jr��~���K������Ǔ��gW;  �Z��        �?�$�{뱕�%���	��n����U2_GH �A��        ���&�Ho����\_z�f��RC> �Z(�        �v��{몒��r�}e)� 떂;        �`ۗ��Jr���T��z� �=
�         k�[)��J�� ��(�        ��/���O�$�L�I��J:53K��    IDAT� xS
�         �S�����{�:%�n���7�J�Ք ��        6�v�G{+IR���|;��{��VɅz� ��;        �ƶ7�c��$�%�^�o$�f���J��+ ��(�        p�V�����&II^N�$_K��$X%WjK �[
�         ��=�~���|'�޿Z%�
 �
�         ܮMI>�[I�T���Z��+Ur��p �ڥ�        ���L�po}*IJ�t��&�J�߫�kK �
�         �����IR�3Y����$�[%'j� (w         Vþ$�譔��$_�r��_V��� B�        �:L�޿�����U�5f j��        � 8��S�um���I~�J�k� ��F�         �V
�_H2U�o��s%�xI�5g �D�        �A�J�h��&�R��%�RI>S�C�F �&w         ֚�$O��$ϖ�xI�aI~�$[k� ���         �������I�J�$�"����*)u� �:�        XO�IM�I��䥒|�$?e�; >�        X�v'�Do�� �w         6��Ow?Y�_+�O�d��h @��        ��uo���䷒�/��J��Ws. ذ�         i%�H��'9Q�c%�\I>Z���l �a(�        �=��I�����FI>Q��s����         ��+�O&�B��J��%�%�]s. XwZu         �5dS����%�F�/&��*y��d ���         w���#I>�d�$�J�%y��\ �f)�        ���p�_�r�����rI>Z���` �V(�        ��w8ɧ�|5�s����KҪ9 4w         �wd����$'J�+���:| �:�q        �ճ?�_��d�����-IUs. 
�         P�{�<���Y�������         �;�����+��Q)�        �`�/���'K�wJ�p͙ `U(�        ��?��Jr�,�_,ɡ�C@�(�        ���p�_Hr�$_+�gJ���P p7)�        ���H�$�O�bI�X��*ɦ�s�ۦ�         k�p�ǒ�z�S%��%����0         X�$�I���dI~�$�9 �w         X�I��$�)ɱ�|�$�� oF�         ַ��|.ɋ%�bI>Q���C��(�        ��0��$_H�RI~�$�9 \G�         6�mI>��%�^I~�$�� 
�         ��=���%9S�/��%i�
��I�         H�f��'�B��%�\I�9 ��;         �z��|6��%�vI>U�Mu�`�Sp         n��$���TI�ǒ���@ �_
�         �[�%��$��k����
��E�         �]+S�O��WK�޺�>(�         wj"ɧ���5S����ڥ�         �����u`�Qp         �-Y���'���?U�vݡ X�        �~y4ɯ'y�$�+ɡ�0��        �~ۓ�I���K%�DIZu�`�(�         �����I���Do��}5g`�(�         u؟��ϔ�J�#%��@��        �:���D��d�$�-�֚3Pw         `Pܟ�sIN��WK�`݁ X]
�         ��ٜ�SI���K%���Tu����        �A�H��$�<ɓ%�LI6՜	�>Rp         ւ#I>��tI~�$k�@(�         k��$�N�LI�T�+IUw( �w         `-j$�x��䉒|�$c5g�mRp         ֺ�I>��tI~�$�; wF�         X/�$�t�gK�Ų<��5D�         XoIK��QI~�$�C���        ���I~=ɉ��bI����Sp         6�}I~!�E�_.�}u���        ��d"ɧ�<W�/����kZu        D�?4��������KI�r2��x<I2�I�I����$C�׶�$�I������$�[���d��4���dx(iu���dh,i]s�xz��L�����$�koMRe�����o� X�IK�XI~/��O�;UR���)�       �������'����ㇳ�k��[�5�d[�����d��J9�F��[=�R�I2��R�p�k�z��f��?�dS��M� �`�3��DI�A�߬���3lH
�        �g������Iv&�ջݳr����$���M�?�}��Y)�Od���%��z���Z�<����kO\sM��>y(ɯ%�;%����*9[s&���       �?KI^b<�=Y.�����w$9л߾�0+m�W��ob$��߷��b��,O���r��F���� ��؝�L�7J�I�A�<Us&�A�       ��,��nU�k$ٗ����Y.�ߗ�`��I�ϓ�5�[og��hn^~����Y�?�6�`MM�3I�RI�E��_%�_s&�uM�       �����To���,ݯ]�L�@�K�U�3ޖ��:}_�9����k֎޵]��+�we� ���H��I~�$�J�w��v���# w���޽��u�w�}�&Y�]�d�ۉ���\`�P(�R
��K��B�mͶ;���v��@��r\�PR��dw�
˖�z�mZHi	�v�e[������Q�m��s��H���q�����<l���{���׀�$I�$I�$I�$I������wg��2`3����y�lT��r|��F����� � O�ᇁU3���:�+I������G"�:�� �)�$I��wI�$I�$I�$I�$5�8���q�>�J��9�^K�ϥ�9���J�}����ߟ���@���J���	�xo�;I�&Ijy�%I�$I�$I�$I���#�3�\�xf��J�Y@GC�K�8���q>*�߇�5TB�kf�UT�t��$%fx�X	���7�$�ep�$I�$I�$I�$IR��;s|n�ǲ����T�W�� �����ӝ���<�k�r6��n�[�a"I�@��ہ���� ��rM��r�'�$I�$I�$I�$IR+)��}�ǻ�k���Qir��M��j�/��5Y`%����q�̱a����+��E� �x]��	���R�I�Z�wI�$I�$I�$I�$-c�3ǬN�Y�M�s�C%���(O�s��,���s��N�X�m�%��2���WG�"p'� 1ݲ$��p�$I�$I�$I�$I�bu���1k%���l����_Zk�9Φ�J���3��g�W(IM�f�O���~��S�I���wI�$I�$I�$I�$-%��O� Y�2*����R�"p���q6}|w����$-� ~%�]�o8�rM��T�K�$I�$I�$I�$i)+�t&��3�<�J��%��tJ[|� _�9���ww|�����F(I�s��/�v8�rM���K�$I�$I�$I�$I����q�̟W�t����!���#��f�3� ��t��+�+��ߗ7�@IJ�
`�����H�%IR��K�$I�$I�$I�$I��� �|��S�k�8ƹ;���v�|�H��$��6����"|xw8��IZ��K�$I�$I�$I�$I������x)�
*��ޔ�Z���gꦲ��
*�����z�Kjj*�O~(�g���|�5IRCp�$I�$I�$I�$I�.�~�ޙ#\�x��~���8���g�?. �x:�>��eTR���$�r����� @)ݲ$)y.Fl�7o~'�I�;�����g.�i� I�$I�$I�$IMo1?;�1R*%�����~��:�����T��?�M��K7���Ug��:͢$��� � �i#IIqu�"���$I�$I�$I���c)U���g�k� ^<�;M�8�3�\�T��7�t�����V'I \
�6�+>�p4�$��A�$I�$I�$I�$I��f� }T:����+źtG�f�Y9*)ӹ�����W'i���5�G��x"�$�n�K�$I�$I�$I�$I�8����ہ� � ^�L�.ͣ|m���� ����.B���Tt[�[#|�� ��\�$]0�$I�$I�$I�$IR�&�O�?|�����R�K5�3s�ٜ�u�P��>{\��wIu��,�3>�J��M�&IZ0�$I�$I�$I�$IRs)�� �^C%�~C�ui���?�,C�������	|*@L�,I��wI�$I�$I�$I�$��}m��F���k�� .K�&]����x:�~#�l`M�K��x��)��> ���rM�T�L�H�$I�$I�$I�$I��#�{�4��
x7�X��.��5�ǀ��j�UT��?�J�:I-�:��G"l�БvA�4�$I�$I�$I�$IRk���~	�}�(�T����������ʪ��><Ĵ���j�;��#l���#$�)p�$I�$I�$I�$I�Z[x �
�P�B�>p"͢TE*��n���|8�Zu�Z�
�]T��;#\�vA�t&�$I�$I�$I�$I��Q>�X5��g�d��>M%��2��J��[��rx,��$5�������pc�I�,�$I�$I�$I�$I��4F%��r`p;��T+R�JT����ꆍ�j�`�2����4#���Dxe�IRH� ��M��Bxs�uHI���\�|��F����֨�$��Q(�.cQ���fzz:�2Ԅ:::�.�|>�v	M�T*Q.�7uV,���Jm�jLLLL��c|||�'�5b,I���
��Mռ6�@�OY��1&>N�Bd��T�%%�ٯQ������(��5�\�|u/	�]�c����c�%)Y����ߝvRn ~x��Zb������7͝���`�����I)0�.�!FGGo!|�A�ŋ.����o��ì]�6�2��{��w�޴�P������k&�app0�2�ʱcǘ��Hm���z��<����O|�X,6�F�]o~��ӈ�$I�Ҳcǎ����mmm%�EJ�RCƫ�5k�p����ː������\�R(�b�ER�����䩧�J�����d�ن�W,)�վ��e˖\�yW/IZ꺁�R	�ߐr-JQ;��3�s0�.	�o w��T��HZ:���$I�$I���Ӯ�lB�r����ehh�p���5�)�`�]Z�f�5��g��p;P�N������I�"Iup�0��Ww�R�H�� >l�tR�O��s3���$]��F�aU�IZ���$I�$I�����{ xV�u�K�|>�R��|>���t�eHJX3ܛ�&I�5>>���p�e�$�p;P�C�|�;�R$�޾F%ϼ��J��(��"�e*+^���Ӂ���J���`�X�{#\�vA���yr#I�$I�$����R�d�A�z)
-rf||<�2$5@�ʛ�I�xꩧ���O����n_�޴��M �S�5_���Z�R7<�Ӂ��e��� ��&��
����?#</�$-N���F�$I�$IR�	!����&Yʼ��|��W����Ç�]��i��7�L&�봤ƈ1����k>�ͦn_@��j�/I��u�6`5p+�P��Y�>�\Si��a�[�%�q2����G�J�7Dȥ]��ţyfG%I�$I�$-6U��B�P(4u�k�����C���f�KZ:�;���H�e�S&�i�ŉs���i� Iu0F%�|5�ޟb�������V`p������X���x�Q��wD�I� I��II�$I�$Iuw�]w�6V��f�g2r��l2400��#G�.CR��&X�,uHj������/j�p��]�KZL���W��;1���x�ʊ�[�A������)�%)Q���E��ͻrVR�sFR�$I�$IR�e��H����f�M�l� ����f�i� p���S�N�re�e���|S,����c��eJR}|x�@�[�o�Z��V�"����{���U%)A}�;��'�Ui$��8#)I�$I�$)	/����T��la���A����5C��YB����ɓMu�f�MSO���!��c�]T:���J�w霎 ����6'WQY)�9`:ź$�]����@��Dh��zIM/��QI�$I�$I�ʶm�21��]�B���ri�qZ3�"��B�/ j����t���7U�f�'���<�T��d����� ��O�y�t^_��g%p�a`o�EI�����m��w�J�wI:'g%%I�$I�$��������Zޓv��L�\�)j����ȑ#i�!)Ei̛�Z()=SSSi� 4Ͻ�\5��<+$�q�@���(0�n9j����[�����m����^Y���b�}��"�+���b�]�$I�$IR]�����=�X�����ٙv	�R���1퀽�t���144�jͶ���M� IJ�c�V`=�n�UܪZ�{*�qn��b짨�O�X����n���^��&�%��YII�$I�$I���Zߐv��l��l�u
�=�����C�s�� �Ei�.5�'�l߾�?�Z$�E�҈�"*�ƽ�V��t ��^|ؗfQ�.Tx1���#l�БrM���3��$I�$I��&����}�p�tU+V��T*�6���fȼY�͒��ѣ,[�,��u�M���|>�1�R$�Ռ;�T�q�k��U��n�P���n��i%�Bmv {#쌰.�$��9g$I�$I�$��;v\F��֢��dRx��Tƕ�Y�*��X�r�+V�2v�;�O�u�J�	�"I�j�J3�+��9�r���T��ۨ�7� ��+K��� [�oD���&�$5�3��$I�$I��&�������Ki<{zz8~�x�ǕԜҺF6�YR㍏��2n���̧�kd&����$�]	�8p-�*��-G��#���s����_*��$��<�Z�o"�]���ЖvQ�À�$I�$I���	!ܼ��$QJ�d�ن������1%5��:���]Ҭ'N�����1��I���V.���.I��O7 � ��n9Z,� ��C�O�&�,J�B<�`��.N� I�rfR�$I�$IR=-��{3K#\u�ԩ��'��5�uR��������}�M�����%�:e�~�J*Y�o�[������+����o��0RK饲1���W����%�׼{�I��T*Q.��.�l6����R�)��LOO���SSS����j�J%J��7�;y�$SSS�.��s�\4��H�$�c���+��b͝sZ��-��,�w!z{{9y�dCƒ�����t�����
��!b�վ|s��H�"T��E��c����Z�����ˀ�^t�X���e��9�����x<ݲ$ՋwI�B���e�T"�p�����������=���'N��Ocdjj�c�-hz���Xm�0���d2UmB�P(P,�4!T�Pn�ׄ�:�^�	�ٮ�������d�Yr�\S>�,�J������_'s�n.�W������YM|����}�T*�R�п��j��$�ϟ��!055E&�!�����ٯ��׎�];g_7���L���u(I��TLOO�B�Zឩ����.&&&2���`�]R3�����G�&>V���Rc�}��ݻ;���7�H�&IZ�f;��	���j^\/��8�əcn��G��)�%�j#���#��a���b)I-ʀ��Ei6�=7(;�ϳ!�ُ�����F�ccc��w1��7�ƙ�tn�l�B�@[[����7�a���4���LNN299I�XL<��כ�^O.�[�B�������f��xM�\n����*I���B7/�}�.������l�X�t.�pm��x���	��B�j�V�r�|�ʑ��n�Jwޏ?��:Պ�(���G�E��Wm)�%�**kT^|3�o��t˒��%5�ٰ�l���@_aذgϞ�
�ZX�Tb||��V��L��˗���I{{{"c�EN�8��'RKi�e�����}4J    IDAT��X���%IR<��7�ʮ7�u&�H�P(�PW�wi�뤤���eV�U�{���S.�/ǀ�$]�)�7��n�	��Y��S<v�~�x	��p1�>���� �\����̀���}��e�|�ozz�/�������r_���ʸW�NH&�0XR���������.�+�;v���1��c|4������H��H&�9c<R*�����#���O�r�-n�&I����ݻ;���j|���d(
	UU_�����|�r�ʆtE��z&&&:^6�%��7tLI�/��199�x3�|>O6�Mt�z�1ֺ�ίmݺ���G��������`[���Jg�a Oj!�
|�� ��.F����U�Y�s�==������j�&��c�;���@�����"�������m{��q>l�]Z��T~�?<<B���b��ŷ����V'I�R3::���gk}_+(���k�йk֬������!��, @y�Z%\*�񺻻9p�@�c
���n�Z ��d˖-�N�IZ�.��$��@���9.O�IU;	���� �[�&��$~�7��X,� ��"�F*��+R.KR���,CCC������r�́7�*-Q�!��*�˟�1~�-oy˾��$I��s��m��j}_.�#�k�M���"�b1�1KtI�����K:���A���$:F[[��7�Zv�	!|c˖-�.I����� �O�-=W���W@w��H����	�o��Dk�
H���P��c��n |R!�B�|��^_,y��'���J�2I-b:��'1�nٲ�/CKv���������c�/�X��ںu�S.S���cǎ�Bxa��k��I�s��|�ݰ$��wI͢����{�&:F��W�T�.?1�лe˖�I�$I���v���ғ�-|�c�X^��]��y��E�����N�i�3�%m����@6���d2=1�@�\@��k3�L.��5��Gc������ozӛ�7��0::����ǀ֙���CCCttt��u�r��{�2=�������r������eڅ$af�`�T�d2C!���r���f���|8�x_�X������`�%K�Tw۶m�����[!;G+u�L:�b�
N�8���%��Z:�C+�!��
�ccc�^�Z)�^*�j��d2Ͻ�۾�`I���借��関%�����QeG�7 /��R+8 �>�{��v1�R�O��ھ}{&��)�p=�	���g�z}|�4�[�>R�s����ۯ��r�c�a�ڗT�L&����Bᬟ�1�w�^;�K�Ɵe2���v�m_O����뮻.�d2?<x���C~i�֭��|^I�u�]w]��d�\��B���%QR"j/�j͚5<�Z7Ig�耻�%�O{{;G�M����\.�:?��[��N�I�Yu�ފ� �x_^<a��)�Y�V%�Z��2Mp���������+���~����?/�?��d~q˖-���q�鮻���f��1�\*i�
��V�:kW�Çs�ر��Ԣ&�_��[n�z��4�s�==o^�Рa?<22���w$I����1����L&s�Ŵ�Ȁ��4p��Lx�';+�&&&jy�ooݺ��K�I�y�~��|��H�����D����À�
J�������8�r=Ңg�]�Ǝ;��+�����]~wzz��o{��R{*�cǎW�>�N�UovK��y'n��<�L漟?��|�c"��w���i���Y?W,���#���u�O�������g|lbb�}���T�f��s[[�9�绞��Z2_-g[Q�r�L�X<�k��������1R.�O_C�#�61�/f����v�m��]˹�ڵkU�T�=�p+НB	��u����¸�$�l�Ν��t����r�r�*JF�X��~�B266���%�6���0�?�xb�}f�*������L1�/�~��7%\�$��^��J�-)'�� �k�#��t�?KjnG���tv�� ������֙��att�;��A��i����Boܲe��n䠣��m����j��f��󴵵��f)
d���۳�,!��,�L����l(}�1FB�'4�>|*�J�?6�{-���!��.�fr����r���i���x��'N�*���ի�|~�'j�z5q����v7��p����|�\>����r�H4�L&s��0�a��k��f��P�w��������_���)��J%&'')�M���$�n�֭�'�B�ھ}{.����Hw��2��f���$�lv���������P(���f3==����!:::�'�tN�%5�+V�gϞ���j���܁�����[o��n���<�������k��1�{����}TB�?���$��;�'��<�v1�b�la`�&w�}�E�R�S4���|`dd�n��ğPn߾}u6����s�+mmmm�������g��p�� �l8q�����f��dhkk��ɓ|�[�j�������ĉ<��S)WT144����R������R�
��>+�J��eJ������4���LLL,��-�!��oٲeGڅl۶����w;�N�7�z��^���p�=�tLLLjnž�;s֪���)~�Լ�Kj&���<��&ƭv�u����[�l��K�$Uo ��������V�� ��y������/KR<��A�G�.Fju���H:�L����H��*}jbb�'�����}V����ʤƨ�\.G{{;���
����	�\.��f���b�@���|>O��~8� ��ի)
�ٳ���t̬[����^&&&R�CJ��F2����f��OOO��OOO3>>����L1�lݺ��B*��w����r���,���'����o���i�!Iҹ�ܹ��j}_����*JN��ҡ�!�?�ȹ%-���������f��d���Jl����\.�4�B��[�l�'��$I���7�B�d�o����9��nï~x���V�p/po�}i#�"��e���~<���Ү�F�c|����d�O<�0����m4�@oo/���ttt��>��ٮ�R�tWZI�)
�����o~3�f����ߟZ}}}�[������j�Z�l'�ـ��Ω���LLLp���9�Ȳ~gdd��F�z3k�����lvx]��\��oݺ���.B��sٱc�[B�k}_6�%��'QRb�\\�j�*>���%��F�;::�Õt^�B!�z�v�c�u���ٺu��$U�$i��z�NZ���Z�'�<����w��� �'W��:*I���'H��ud���|���1ޒvpM�󣣣k�yҝ;w��,)����<7n��k��+�`pp���6J�SSS���3>>ΩS�gbb���i�H455E6���k�M���'8z�h*clڴ���a������>99�����������Er����\}��\}�լZ��e��޽{;�ؐ��;w�|Y6��g�;������mQ%I�즅���]ۚ]ҡ�V������6/��sIr��V{�4��b��T-���t۽��<���:x5�i���x8�;�u�-�����Լ�Tv_��/��Fh�x����D-)�;��݁���_�+�>::�l�O��z��Z�B��/��͛7���gzz��%HK���8�\r	����\.'ڵ�\��,W_}5!��{�!����I&''����k�aӦM���^o!�7����Jl `��ݝ;v���	�V�8�߷o�s�.B��s	!ܰ��ջ�D%�sH�԰Ml$�*.��4�\.�ع�cE��xݼ����j�$]�c����/�\��� �V�� S���R*�L�<Iu�nv ߙv_�r]RSrvR-�{��1�@�u\�1�?��?8t!'ٵk�e1�?:�T׼r�W^y%_|1�R�P�����i�U9U�|������-^%����!�Ftt�Ν;)��ܹ��b��­�ւ�g�]�$Igs�wv����t�L]�����D�/I������$Bo�F'5.�̶��]�T-�����{��'S�E�ە��+j}c�Gf���~
��:�&)s��ߎ���).`�]Z�Z�)�LLL�hK��:�lzz�3�ΰ}����'�u��V�^��_����]Ť&Q.����f�ڪs����6���
����.EҌ��	������kikK�l�Ν;�^'����;w��e�/���:omJ� I�Φ�����c�.��l�K�O�ϊZ��{�8���*E�T_E�שt��)ע�m-�N�7/��&��{�˩tu?\��$%'C�k�ׁG"|3��ύKd�]:��ռZ�Y��/
��m۶����l&��X��!+�f;�vvv�=YjB�r��˗/�N�\��.�̠�Ԅb�����y�f��.hS�s� ۵k��z�����}��}�E�U�ԗ$5�R�t�B�׊��$;��r���P*i�k��6$5^�όZ��(�PS�L&sS��H���	�ǀW�I�-^}��~�BN��3]�WS����:�&�q6[�/ �#��5�HWjU�N�]Z������룫��e˖Q(j��^�����Zްo߾w�.�f�Z˖-��crr��:eHKI�\��������K��+���p���&''���gӦD�w���Ol߾}�������^RǺ.X���v:;;���aŊ�]�/oTm�$�"����{�ϜW�s"��_��ծՒorr2�kE�ܡ��A1F;�KRk�$p50
$������O�7^��tu�x���=���^�G%�~�7FX�r]R✝T�ٹs�_ /�浽����Q4����$���LLL0>>���T��"?�u��?��w�u��g2��р���Y���~$U�����~xQ�p��'�ŭ�����|�k_K��~�ȑ�m۶�꧚1ưk׮�c�e �DQ�(
ttt���N[[mmm�����i{�s�"�����z��-T���ܹ��9mmm-�,�ˉΏ�X��'N$v~I�C����\���G�6l<I�)�������Ν�b�H�X����Ba��~��$X�$)Y�� 7�]�����:��x-�&��z�[R�=De�����N�����VT��\L��2{zzf����_����A�-[V�Bk��ٵk�y�ٽ{wg&��(�����z�j��R������K���i����dwi����檫�J��/����Z���ή���O��G���e˖188x�~shh�������������)T�����������R���z�9,IJ[�]�%�#� z��.\Kw���)���ھ|��@�w S�	����I��p�k�����Vup�����uV�\�T�Պ.(�~6�B���>֮]�ƍ�/`���r�������s��X,�X�t!+V�`dd��iuI�hbb��7�]Ƃ��yV�X�r.$ULMMq��W���!�_۾}���ntttͲe����Q�L&COO�ׯg�ڵ���Q(�~�<A�U�"%I���{�^Be�䚤0�r�����j4:pn�]R5�^��j�Pj�7%Q�$�����R����R�E��/!��N�*�뀋�w��=��� ~��d����ϋ�O�6iA��������վ~!Ls�lܸ���a���^�/�1���>�cǎk�ے.�����+Wn�Z\{{;���i�� �_~9��.�Z���$W\qE�Oۖ����{�ys�k׮�c�_�1^_����f<}Ym��L�<6�.Ij6�]d��E�X,�]�����wI�H�Z�jw��zmwIZ<nnN�\��7��l���P�p�$Ƒ�0�9T�|8��#��X�!Bjz>MRK�1S��B��!���7����]����7����m�2!��"��Tmmmlܸ����$��� �b�%��n��R�Ć�z���o;��v�����r�/��:�}}}lذ�������3�h�]��T2��5y_+&�V�s��j4z�V�^Kj����K�ZL�	\�Uʵh����@wR�p��P�O�00��x��x1�>�K���E����-M:7�j)3���c[ĹA��ު��_�㮻����?����xv�c����˙��TZ,&&&I����\��c�eH��#mmm�=o������v�8aǎ�!�6�������Ɇ�['�yh^���|$���$-D��ꅼ���������Q�M�Zq����ݕs�$I��7� �'S�E���� ��(��C���z��I�)�a��� � �G�f�{g���-Mz���j5U'5Cu���f��z�����Y,7���<����+9u�]���fŊi�P�60>>�v��\.344D[[[=O�<���:��m�r�v�'��_�9�|B�jժ���ӑ1w�ĉ��:�$I �py���d2-p���L���g�ԢB���s�5��򗿼��Ix��φ.h�TI�[�TJ��nٲe����j}>�����.I�S�J����I�-.7P�!�!]�<�N`#p�׍WRCm^O%��X��s:�_�rmZ�|z�VSuФ&ܗ/_�E]ēO>ɉ' ������7�ځ�X�j���I!)%���lܸ�G}4�R�+�Ͳ|��Ļ�Hj���I.��2|��z����;w~xK���<�|���X�jUb���T*=�ʶq�$�jtt�-Ƹ����b��B!�Mb�����.�l6��� k֬aݺu�C�G�mx�S�N�f�֬YC�����㏳g�N��	�����Fuvv�Ts�BM'!��O$[�$)E_���X�n9Z$.�x)��F`
��?��[�\-->#T:�� ·��SY\�7����B.)Q��R2��p��A�t�� �l�U�Vq��A>��8���$hoo����P���utt�]¼6l��uHZ����ټy3?�p=O�g4xG���NFFF�J6_�³\���6�k�[l���@�?�
���|�rV�^���+W�<��G�mx]Ǐ?�����r�7r��!����޽{9t�P�����K>�grr2���"�L&C�T��1ƛ.G����n�	|�7�V��b�?�ˀh�������#��#���`#k��P�tx�̟�"�� �E��Qji2஖c���Iw�X�b�|�$5��?s$��K/m���j755źu������v)������m�%5V6��������z���O6���L~^�����%IM�\._����b8���/g5�7I�O�+V�����?<7l�(���t``������j&''y��'ٿ?{��q�YZ�����.ĵ܁c�!��j!IZ���O�{��-Z솀���Jд���E�5�U�[q��t7� Dx�J�}6��P ����ZJ�qe����p����\.�޽{[�K͚5k|� -���Mp_�v��vi	(�Jlܸ�|0�Rj6�h�*���w�}�[n���'��$%dA�V����f�y���$-LWW+W�ddd���������<y�b�8o�mmm�[��u��q�M7q��A�������9t��;VK�]��*�:u*��'���޾]�vm��P9���R����9�r�� ��-�4
0	���y�[��[�ۅ���8s�vy?�K������ ��U�Z�w���j_؈/_������k����\���~C��111���H���200В($�n||�����o}+�R����۰p;T�{e���u��x��'7_oXQ�$�E��Z�@Z�{{GG'O�Lt�:{Jj!�����wvv^����C��{oooկ!088��� �\s�b����~�������V--FI/d9~�8}}}�ߗ�S���1ƛ0�.IK����nZ�+��M�'T����YH���*V��[����Y��T�/�9 �p�*�����/�Z:�pWK	!����Ut�����N���ٿC�]��.��p���4c����ӝ$�%����\.G�XL��y���044��q���y�n�R�Z�K�Rc���{ҝ=�Ј���CR����dxxƁ�d    IDAT��+W���S�󏍍��|��[K��L�\��+W�r�J���:&&&ؿ?O>�$H-�/�����)��tvv�T�*�~�]B��x�I���8� 𧁏 #閣W ��JG��J�<
l����7SCcSI�Rp��@�}�W���g�� v��w����tww3==͡C�>v-:::�&-A�ry����nݺ��J����I6m�Ŀ�˿�]�y-[����t�����y"f2�k�?n\E�$=Ӷm�2��Z�B�5"k�N}�L$��e˖188���������'6V�\Nm��z�I���Y�~=�ׯ*�8p��q��і�%U��b�5����-��V}�c�1�r$I����TB�?�r-jmY���@ʵ �����x;pU�UIj"#����#<B���׀������S�Zo&@K��ݻ;��bU[�d2�Ժ�011��]$.����KKP�Xd�ڵ|�[�J���Z�����
!P(��[i.�cժU��?�B��5*E������Y,��}/��O�|���9u�ccc?~�Ç399Y�b/P��'��������200��������ɓ��再7׉'={{;�֭cݺu@eW�p��A�z�)>�ܑ�"�����eٲe������N{{����~<��B8=�3��}���/|��a�c!W�H����#���@�~��b����w�\�i��{#�>�2�?/J�*IM*\1s��;T:��ʎ�_p���!��eLNN��6��F����������ݔｽ�M&������K8mpp��6�U,ټy3_��W�.廄X�jUj�%a�{�µ*E���
!\\�{���8�kN�:šC�ؿ��.�iK��A����-�ϟ����1<<��s�!�f�P(�f�֬YT�Ǐ�СC<x�p�ر��$�:I/�k��î�.�����룻����.:;;�=>������ݻw�_�`����^�TB�7�\�Z�@7�f �U�g �>+;�<���&���9^>���P	�xt�����EpW��f�+�}m�PH��y�r9V�\ɞ={R��l.��"����.CRJ����f��J��Kapp�)Ij�r�ܔ]����ioOw�l�{��ڻ�{��o~��$I�3d2���v�\�bż���蠣���k��Ӟ={x�'ؿ*??LOO'z�B��ZWfI�B���~������������z������N3\��iOO===lܸ���I:��ÇOͼ���T$p?u�T]ϗ��X�bCCC100�� ��,_��e˖U�\�\._�wIR�c���R�iՔ4��]�����|��[#���Y�7ݪ$��>*���\v$V:�c��M�|����e�VV��4��Py(��Օ�Ç3-_��)����8�R�����X�����KKX�X�K.ᡇJ�����<���i�Qսl�\�
�|��H������ZL�uo?���v.��.����"{����Ge�����_�B��x��|>�\��@mmm����������ٙvY�J3�݌��6V�ZŪU�N�����#GR�KKM���k666FWW�ݟ-[��5kְz�jV�\ِ�tV�X�w��^[.��>�lE��R~��1`$�r��~�^4�DT�=�~�i`+�>բ$-}�����(s�<3����E����e���j����%\Mu���8y�d�t�ڰaC�uI��x}}}������Hj~�L�iv��ʽ[��ƪ����d2��C^�wIRJ���~>�\���׳~�zN�:�c�=�#�<�h�;&���L&CWW===������GOOO�uf�V�MTf緛�zu�����4G���ѣ9r���6\���tX�T*-h^9����0�6mb͚5��Tp!\�p9����T�	|���kQ�z%�	�ǀ궗IA�1`G�Q���w ߛnU��^�ƙ�"LQYx��<:��|+@�u�X���e�V����F<��F6�e``���z*�R���M����Ft:���ի��I隚�⢋.��GM�:;;Y�|y�e����v��c��4�I��!Ƹ����s�������J���
�x�	z�D�^�aᛤ��d2tvv���s�������ٵH3�c�ԩS-���L�|���A���1�=ʱc�8v�Ǐ����ߥԈ�n-;8�r9.��R.��2������j��Ȁ�$�<����| ������>C%���UP����'#<��J�N�Ij��q�8�+A�ǁo�� ���5��Ժ�pW+i��;@oo/�N�3�ƍ���T�˖-;op2i˗/���$���X��]=
�����%Ii�Pˋ���	�X�fk֬a���<���<x�n�oD� �J�)
tuu���>{tvv.� ���8q"��O�<ْ�s����v��g|�ĉ���=#�>66���ZO>�����|>���޽��U����<�2�芤��@�����c�&��ip��N����/c;u�NO+���q���y��49�q.M�6'�݉�$M�؉Ǹ,0`$hFs�{����#if�Z���z�����گ�F���1��g��}~������l.v8������S� Z��N���y:��V�v�M��bvv����ŏ�*��Z�ƕW^�UW]ŉ�YN2J����Ç����$i9	p7�g�a�Н���G7�~�lɵ��3�g8�8�F��!�\�n��B���%��D�G�ߏ����^�8�>2�U!��<�k6�Qu�
!�e��~��R�q!^Ң�;w��#��]�$1==͖-[8q�Di5������k9):�]�}�~�w���$�P��G6���d���k�Z�ڵ�]�v��c�����}�[������Օ�A������㌏��q�F�����8�:�SS�x<99���D�5a῿ݻw���V��ɓ'����IN�:�f�0::��^������Ǒ��/u:N�:u��Ǐ�ĉ��ߋ����i�֭|˷|KT����fvv6��m۶�ʹ,IR����#t��RV�
�!�J���J�7�?I���~ ��xfI:�F��_�J��ݗ�����o � ǁ���m]3��H�$U�,�e�֭?~���_+]�;zH:W����f!AIձgϞR�1=�\����ѣG P�$I�fgg3w۲eK�,k�޽�ٳ�|������ϯ��R��΋��i�,�/�C7nܸh�q]7������� _�F��֭[ٺu�9�n����frr���)N�:uƯ���J{.��j�###lذa����ht'E�j�7dLOO���O��SOq�رBO.���֕:ġC��j��`˖-=z4��$I`�]��۳�w��G`C�娂^��r��%גI�G�������~�?6G�ⴝ����NН��q鯏������	`8<s�xݽ��q�g��jl޼��Ǐ�r��{��PVRu��Pf���>ؓt�Z�F����B�ؤ����t�	�u:�˲��6oޜS5�!p������g?�Y}��5�O����?R�5����^6l�. Zewo���X���Š�r�$azz�S�N1==���4333LMM133��y�����h,vW;'��p�[�a��1::�޽{ٻw/�݄q��1�x�	�x�	�{�\����f�fN�Z�뮻��v��u���w� �;9�#IZ_>
�%��5%ע�
�ݐ�c%גY����%�����\RjQ�T�M�_�%�y`8I7�~���g��瀅�I��;t����/�����?[xϥf��W2s��pW%|�CN�$�y�E��ƍK�K�����i�&C��0;;˅^��?^��7m:��r�l6�<�&�c�$I !�}Y�N�ܗ��o�k_��g���{�?���@]��`hh���!���⯇��h4�K�]�Cg�zhh�N��꿗V�E�ӡ�j�$	���$I����;���������Y��444���0��Ì��,~\���F��������ɓ'�.���y!,��W�n����eff���fgg����ǹ����ܠ	!,ރ�Cgo�Y���Bt��uv����ݻ���k9y�$G��G��g����9u���nC�t�M\t�E%V�[��p�`��H�֧/7 ?���ZT=W L7�^�SdB7,�3	|��?�o.�*I��&���+*�<�����Z���_�������V=>1v�t�V����(��ӽ�����v$�m۶�p߸qc��Lc!���<.�pu�%I��`OֿPV�}�E]Ķm۸���yꩧJ�e��7�6�M����ymذa��m:r��m���b~nn��u:����K��V�v�}Ɵ/���l!`_�Z��0Z���u��f�F�A�^_�x����&���B#49yv����a���멂�K�Z-fgg���gnnn�5??�x?[z[���Z-���!,�̹p_,��}ka����h���=��M5���ٸq#��СC�8q�|��~�o������n���^���0�p;d>�(�V����M��!�3@������ܿ�J���]�v��/���� �QnU���a�]�P��.L;6ր;t;�� uǎ���%U�֭[K	���.�����{���X��&{��QIR9ve<>>��۱�1n��v������~�����Y@4!����lݺu�m�6FGG�.�/���b�;o���K-����t��,P�ը��g|n!ľ�ϥ�/�py5�\��~Zz���)����]���ξw-�~�+.[�l���E/z�>�(_��y�g�.+�={�p������e�g�$��X�$i���<�q �)|h���~;�7%�r��ܟ���w��È$UL�O��B�y������x��F�a�]Ҳ���K�nQݠ$U���\pO?�ta�+�Zkѫ{f�$�}�{���=UPI�$A��ewo_�V�q�70>>�����c�V�I��ܹ���	�m��֭[�؄�,�:Ʋ�A�w�ԩ�KX�
n����V�-n�������hp�e�q�e��o|�/~񋥜��V�^���𒗼��RR��l�픟��$I����_^Qr-��	���o���Z�"t7|�)���]�룫�$��ϐ��Rup�}�uhh�� ��͛K��,�ʸg���R�n�����B�����2��O�FFF^PD-�$-�;��͛7�Uǚ:t�뮻n�1E�.S��d!v����_�b����;��[n��+���;vn�"C���.�;vp뭷�W�bM�4El�����߿�M�6�~�~�0/�p�=�lͳI�@x
x5�>`�cx��m~���B�)�áp�����˭H���O/T	I��zx{�`tt�����-����Hx���q�K�VT�\�^�G?wLS_�$� �ͿI��jB� ���W\A������������7ϟ�j��w�f߾}�ٳ'�y����pߺռ�4(v����_�r�|�I>���q�x���������֖$	��yظqc�S����^]I��_�n����"�ಔ�����Pr-}�p8���x7��#IѲ��*!��.:�C��Bc�J*�\Et$<�訧}IZ���\a��*̓Rܯ.�I� ���?<�g�;ccc9Us����*���e���n�~�<N�۾};�_=ox����[���K+�^&iy�V+��hZSSSe� ��v��U�z�_}�9E��*��f|<�4�����$��o/���BT)c�o �,��<8�n�2�{�/�\�$i�U	I�������Ha�*�ۘ��*�Q�=PR��Z-v��Qȵ�p?��ji�����Z$I���3Kmܸ1�R���k�墋.:��U���h4����yի^�+_�J8���p_�[R�����.aQ,��%/���x��^ǁV�b�U���,��$I�K���Q��Ce�J�@7�����K�� ������,�$I��U�&�^T�ccc�t���":�͐��^�m�V�u�x��)��%I��t:������!n��RNw9ߓk�����o�&^����җ���y����*�)l/�CCC\��|۷}ۊ����}ff&�k�!K��'[K���,p���\ɵ�:��_�Xv!y
�	p_����O ��Y)I�wUEυ��.KW��
Y�����lI�(#�^��OR��Y�
�FHU�ޟ��6�&I*J�����p%��6�M����¯�ր���0�^{-���9t���uljj�����T�]�vq�w,�ͽ�h�~�V�E����:��%�\�W�$�	��zم�2��/�_v!Ep�� /~���S��	��G>���^�н}Aw��<&�Z�$9Y}=I�S���������U�"I��,�c�޾Ԟ={���K_Ĝ$��G�F�����׽�u\y啅�$�+�PyL�H*����o���5�"�$IR�S%2�{>�$�<�)p�?�.D�Q~x{م%��	8 |�cI*�wEojj*Uw������Z}�))����%�277����F�Q��Q���!�C�"II�l�2�j��:D�V�ri����^�k_�Z^��U�+����)�i�]�r.��b^��Ws�݆�Eͥb�?��l6S?!d�wK��FO �?_r�� ����.�H����x��$i`pW��ƞ4��p���N���5$U_u�*2,"����6[��ۤ�J��4ܓ$���R$I؜ep��7n��/���i�&^��s�72::�{M��S�szz���$U�����~;�_~yaU���&�|.��RI���,��t�rϗ\��! ��?�.�h�
p�n�����V$I�_u�XI��
��	��"�PU��`nn.�kH��z�N��,��{�V��hT*\*�x�7g��eV�{P�^OS�5E�"I�i���H^u��꫋�7�Z�=���W_�w����Da5I����L�%,J�$�������u^�җr�Er���3̏�K���3�ˀ�e�����O�]DL��x-�ْK��u��T��6{��R�4��ǖ-[��.UT�^'��<_�/}-����¯������<�@��|7�p���[�I��j��t:t:���⯗�y�$��;��&I�������Ť�ɻ�k��Н���ή6�PQ�H�[�$���iT1�e�����7-[�k966ƍ7��Ν;s�AR�b
�C7PZ��9$k||���Tu�M�y�=�P����\���%עjx��?^v!e���K�&�_��(�*IZ_�+zI��I��J��CUE- J���0��=�V�BX6<���r�K?���"�:u�v�]�5�Z��}_��	����a��������/}�����O��ê܇��zܷ}�����w���E�$IL!�LǬd�D����r�]_|17�pC�mI�S�wIZ���P!׉���V����<�$i�� ���rKQE��n����]H�Bw���	�x�=@�IZ�|R��.�5f�+qU���}dd��������/ї�݅?[._x-�yv�|=;y�d��,��NQA��-������v�_�2������1g��3���&U�z��f���B�0�.I�[�N�U�1�>;�B��/|!W_}u�זT�u(6�.����_�p�p�Qu�zI�֣����?I7�,����f�	���>�)��o~��1��	�z�R�v ���z�@�yZ)ܼ~��>Yd�Ж���BW��B@|�Ґ�r�����K����y�8�orr��kNMM~�2ݕ%K������������9�����ˍ=�}Ζ����ￚ����]��j�[/l,X��i��ԕ�׫j'-��_	�~��H�\�����p^u���)}1<<�8��[nabb"��J��v�}���1�j�TRq���^�|-6��$iu ������kQ��F�>��!��o�_��ȸ�*I2�j��k@��y�ϛ��Ƭ�$/�>I�U��g���p�jA����ϝ,\.|�����9���'�2:�Z�=K�Y6�(_��$Y����V�\�{�I�����q�F��k[�:g�s����'+����Wm�Aʇ�/ȻI������S?u:���s�"�a�    IDAT�=44D�$���s�m��i�ω%�)���gM���&ﵗ���\�?/�g6�$	!�j-bI�֣�n~���RT?�O��;@����~
�~�ݤ��I��L8)j����_���w�W��y/�mٲ�������ATF�|zz�$I�T"���ުm�맥�������mS`�N�I��݀�$��R�U��,���^�b˖-�x�lذ!�kI�����X���4����U����Yܽ��� ���J���������Rr-�������@\ǒ�(�I���#���O W�[�$�/�VD�y:z��)6bT�iޡ���q�l�¦M�_|���.����h4�/I����I���KҊ�����$��+u���r'М-I�$I�:|���i���E܇������KZQ�a�k��"�RU5���y�s�=W��^����)��G�.D��=�/a��s�����^�ϒK���pWԒ$ٛf\�v:B�۷/�c�GFFr}I����d)�-�s�����ah��榛nbbb�N��{��R�ww�s�=[��E�4�v�ޝi�^��q�\UެZ�Iŋ1�i�]RE�s���+wBd��lڴ)�����A3K�+�;��}#V���
f� � ��x��@�,%�`�`��%I�'͸X�I���tرcXj}�s������ù���������S�J���j�s>��th�Z<x����s�������F;�l6��ϯ~*������S�$i����f�&Y� w����CR<�K���69���U��S�9���T�v�J����c����\���]�(��n��2|
�T��?D��&I��Z��{!����v�f�ɡC����[�����B�w����%U���,�V��kOOO�r]IՒ�����M�6񒗼��n���h4h�۹^?�4��z���J�$�V�5��~N��\��������K8�wIi5�)jcb?e�#��mC`����w�[�G�.D���׀j�L,A����x�t�IR��JKg	!����uBE���V�E����/��/^q\�$�>h6�>$��SY������t�ް�ҽh׮]�ڵ�N�Ñ#G��׾�BK� ���\Y@)��5::���,�{�Z�*�����*�1�j:�sss6X�����9�5'H#�yӦM��t�$�L� �:��%ע�����9�C�c��> �#�]��V%I�0����5����I��$	�v����/O�h7==M�$��T��%�À�����}9�Z��.���.��S�N����ϖ6�L3�!��]����ܫp/*Pj�]R/1vp�nw�VS�<���34���-o��?�$i=��g��喢Ƚ�m�5�dɵTB�)��~��	��J$i`pW�zvp/z1=IZ�۶m�/xA��U�0���;&i}��,�gƼև��4Y6�lذ����% <��<��Ü8q�а{�#��K�r��t2}�ᴽ�(*�^� ��s�}ӦMe�!)bE���x�E/�q~�$iy3�? �eɵ(n��I7�m�=� �>�n������uπ�bE��P�֭[9x� ccck~/�bPf���҈)���͛y�_�3�<�C=���d�sҔ��/��/����o�xGIR�u:�F�PvU�vp��X;۸@R/E��pϰ	t6�:$I�A��<�Vv�N�N�\K���?��t��?l(�*Iʏ
���^�| 8??ϦM�8x�`ߺ���4�.)����Үm�]Ry�i��ضm۶m�رc9r����\��)缵������� I��k6��v��z��Wg�]R/�vp��.I�(j�Sŀ��%I�?�<�I+�	��U�s%�RI�J�_o=��^nU����{�g���|�V��^(���g||����s�������09Yމ_�%�144�����^�s�Nv��	�ѣGy�ᇙ����l�����y;��0�.I����|���c�]R/�vp7�.��}awIR��.p3��ޒkQ�n�x�LɵTV�o ������ �,�*I�������4���!3�P�Rvp��2;��Z-�������>������yn:���`bb�$I8r��?�8����5o!P��I�9�k��$I�H�$S�2I��J�U�.�磪 $'� y��{I�(j�SԼ�$�u��$�?� |�	�E%עx]|�x��Z*-t7H~4�_^���ܪ$��pW�R��\k'���y6l�����ٱcǚ�c-�K�AާI��Ϯƒ֧�up_N�K/��K/��$Ix�'x�ǘ��^�6e�ݮ��\4��S�N'��,c��%�k�|v֦VW�<��*3̑�˳I�
�8p+�߀��[�"�b��?Ur-���:��	\�(����R��52�h%I�'��s\���v����8�^zi��W�w�Ԁ��^fggK?�uzz�M�6�Z����=������j��4�4B�ٳ�={��;v�#G�099�z�O�y��%I�h�Z��t�j�����K�%ր{���%ţ�yN�j~6�:$I*г�����iɵ(^/>|���kY7|�+�	|/�c�E�V%I�pW�B�:���p5I:�[�l���/g||�o��U��B��v*������.����WĜfzz��7�~���ܹ��;wp��Qy����Vܧ|@|��>����w޹���$�^�Og�Y��Ww���S�ӛJk�^R<���Tq����n�]������лӥ��vr�6�ɒkYW� �N����]���[�$�c�]�
!����4�p�BY��&��\����h�w�sdd$���T}1����#����z=�PǩS�J�/511��� ���9r���z�Z����R�G��}�ù+IXo��g���)��8;�K�C��v�(I�)j��e�e,��.Ip�x�y �Ѷ4W��r��R֟ ��ǁ�'p-ݠ�w����"f�]�J���^c:\�Z-���ٵk�\rI�]�fggs8[�_R|&''�.����T���s��h||�k�����9�9±c�h�Z��j�+1�.I��4�jwXGP\��%�&�MBvp��KQ��+�0�|.�:$I*�/O �l*���
�S���v�W�%�~���[���V%I�2஘]�k���(W^y%;v�(���w�v0�.��"�E��*����333��w?q��A<H��泟�,�<�L��z ��$I�)�U@p��9��8ļI��z)j�Sŀ{�9��%I�� 7��)��� p?p�ՒkY�<	N��o~��r�����$E1�9�ݸqce��PL�thh(�kH������K0�.)���51l�I�^�s��B�<�r$I�+�7�V��g�gwI��9�Y�L���<gei��I���]���}�n���e�h�>�/���`6�G�����\��T:��/��/� �z�)����;D�l6]8��S�*�J%�'�^�6ۤ�z$Ib�]���B��{���fwI�i��e�������K�9�9+K�I�V���]�4�
��Iم(Z�|�U� ���� p��$0W��'O�B�q���T�?y������T��U�J*��ϔa�w �:$I-S'I������������D��T���9!�|���`��]�4(�^|��B���?�*��A�� �v����$ ���4���6�.)1:���tH�)�M�6�d�z\r���|wH�R�$Oe�!����R�<$i5��#b�K*���e��%S�4HN�>Rv!��.����.d��� ����%�%i@pW��$ٓf���hޥ�UޡҼ��J��V�EȤ��x������T-��a�[߾}�%9�"I\��U��^Š���'���%�ƀ��2̏��.I4m���-�Ek�n����d>�-�����$�s����Z�r;�K*[LaΙ���K��f�����tOL��lR��S��t:r.G�4��vp����b{�<� ��rp_Y��q��y6�R$I����f��C��	���K� �xpݮ��z�*��+V��###y��Wy����I���O�Ȣ�aI�ʻ�{�ݎ�T�,�~M�$�<�R$I(��)�>;;�W)��ՊY.5�.i5��#�K��z�7�MAv/��jy;���U+��tW��~���K���pW�Bvp_�z�)�^��ɒ��w��w/J��3�`�]��wY�U��ZŠ�$-� ���P�y[���F㹜K�$)v��
pӗ���}�������*��ہ���4&):��$I�]�N����\�רZ�_R�b
rV1�"�XElދ龘F��ށ<�$�od\���z��������EkewI�)j���r9)סZoy�[��T#IRy��	x��B�-��/-��)@'�'�	��<RrY�*ʀ�b��:�OOO羨gwI������aI�2�~����$I��.I�v����{���F���T�㨤��jq?�1�.i5Eܫ�L,���N��$=�o��,�Ei!�~Cمhy����e<���EI�ŽJ�A�3��l6{��E�����'�X19��.�����ܯ�}1���ѴC/9|�p�_@I�@��j��U����dwI�1�.�ʊ��T�႔��y�!IR�|����Q�6��ZrZ�Y]�/������V%�
�^%�@��{�=�;U���<�-"&����.�J��~�s�����/ɱI� �t:��2ހ���KZM�<x���+K�&�t�uH�TAO�\v!���	�ee��<v����t���"O�ERT�+:333=������]J_�2�.����U�H*��ϕe�g��9�c)����w�����g7�p�;�KRoU���ϧ�f:5I��r�n���.DQ�^^v!JgIW�7{�� �+�,I��{�T�V��
�W���wI1�)�i�]R/�f3�΅U�e��$��9�"I\O�Xŀ{�^/�I�>�{}��e��eX����$I+��~��B��o���
	p"�������ݍ���+>�ZmO�qvp?W������+I��&U�J*G�+c���F�M�vp�$�]�$O�[�9Qk+vp����7�p����K��$�wI�V�~���Q�F�ܿ��B�6���^��ǁ�r��TW!�N�c�52�.i5ssst:���XT�P��r�=�;u�T���oY6y���.I���ӎ�i�mZ��J%��O�:_�+%�ƀ���΍k��wI�zK�F7+�m���/��]�� ����[�?)�,I3���j��iƍ���]J_��Z�_R�b��j�h��e�!)ryo��f�,�$I��.I�C�{�ݦ�j�YK���]Rb�{}��e�}y���K��������X������.D�/�� ��	�
xp�ܪ$�UHE'm��܋�Vm1OR�b�cM��244����Z-��s�݆��w���|����A�:���LVTWb�V{���bP�gbi��I�p�$)���	P��=*J�����\��(��.^	�P�#�%��*�R���=����n�ٌ��ZI�*�$������.AR���	�i4Y�&��۷_�c9����D��1�����R����$�.�y�|I�*b�B�\�=ü؀�$I��
��Z�T�:�� �_v!� � ��\���۵�����
��$I�*�^��N'�.�yw7�T}1vK7�.��"�U�,�e�j���X�$i ��u�"� �v���H����Gka�]�jZ�V�רZ���;��wI��������.Dѩ?���B�� ��p'0A�k�'��8��+W!�]iU�����L�GOp��K��c�IR\���T-x�eB0�.I�$I�u��:&��Tm1�c�./�|El��}Ȁ�$I��#�e�Se���? �,��+�� �`��O�|�{�ra�]Q��G>��5.���H�a�("�i�]R/1vp��&Iq�����tpO�Ā�$���������z��;q����S�<'�M@+I;/9�s)�$�w	�<^v!�N ~�e�bx"��n��w�Œ˒��wEe~~~"͸���J�ZD����y��c������K��"�8U�lcwIR�����=L�o��p��K��UZ��T�"N��y�JR΋g��ַ��kK��}�n����Q���d�E�X�\�����"�*����tRܳ�zbPDh*���`�]RqJM��EY:��=zO��~�ZځU��*"�%��b]�!��]Ҫ���W�S��������λI���f�%ס8�x�E�^���R��'�V&�l��up/"TZ��<Iŋ�Cq��{Iq)"`��q5�%Ix$�����<�����p�װ���^b�W�k��b��odd$�k�S�9�wI���I�V��K�Cq�q��@(��'���R��+*I��
�g����Д]s$�c��j]�%���D�6�d������&P$I�v$���up�b�vp��K�A�"���yN��Ei��!�gr.E��Atx%�e�(�(𳘡��%a�ˀ>حD*�7g�f]vp/"��I�1LcM��R��j����=[�n�0�Z$I�Ѵgff�t:y��wvp��X�{c�,/)E�s�k�=I�c9�"IҠzx�ɲQ�~�(`gQ-:�����=`'p'����r+��w���k�I񘟟/��sT�k���qJM��EY��!�}9�"I\���$I��p������KXV�uI���ϕ�T��y�!IҀ�����Q���K��+�#�3>�Mt���(�2i�3��p_�"�_����jE�5�j]�%���%��z|��1�.I�Z��:��=Q��E�$U[�M�K�ŀ���K��Yເ�^v!��w�xt�V`&�'�\��;���V&�O��T�6�]G_ѩ,���kx3ֺ$ţV��G��u�!d
���]��oI�d
�OOO�UJ.�op��K���t�z)⤚"6$�S���wI��7��hم(J��@�&�*E�N�?	� W��� &˭NZ�+6벃{�"�_��k~~���k]��Q�&�v�]��Y���wIR�=��3O�}�J�:�������j3�.����~�����wI�������Q��r�V8M��p�{�	�n�<PneRu��Ulv�d�s��]�jfgg�.aYU�J*^Qs�X�+�2N�Ā�$��>�O;�j��K�A�A�X����Q�<�jw;�K��6�C�(�E�ہ���.D�`:�'�7�x���'�j=��Jd�]����?<���l6+��^D��}M$+�N�I�D[��8���B�S�|��2�hd�]��w!�GҎ5�~.�z�5�k�^R�$1ྌ��k��wI��� ��Uم(J�n�}Sم���tw������/�[�7�F�ݞH3.c��t���t:�ܯST�KR5�"�����5�Y�܁��$	y�"ILI������bdd$�k�s��^b��Z��8���J�v��z�inn�X��H�����p�E(J7�l-��N�� op%����'�J������n�w�W�����L!�1�.i517vHZM��(�:1�'��1�>z��w��kK��V�������A�z�5�i�]�j������֋�!�\��w��]՚8K����x7ݮ��R��1paمh}
�d��xK���~�-�ǁ�ʭN*�wE#�pA�q�<�+*,e�]�jb��>77Wv	�"V���M����M��Q�$ip�j5�硨�+ր{�uI�C���8m��2�ft4�:$IR*��Q�Sv!���tC]�ֿ �7t���^��O 6(���J�*$/���%��V�Q���c�:��N�VۗS)��e���&dIqh6���.�U�J*Vk�U;I"�\؀�$Iq�Y�M��u�ˀO�.D�#�l�O��n� 7�>	Tk�]�Ȁ�b�*྆n��2�.)1��vHꥈ�{����uN��t�K��*�p$������&9[�^�}��J_I�!�l6�.-�$^    IDAT��%���gbU���]��J�e�>���.>���B4�L�?���l��x��l�J}f�]1ٖfP�:�����\GR5���KX��I����j�m�ΉC�%I}��3�|��5g�D!�.�N�r�Iŋ1�cM��Q����$� �x0Sv!���i�ƒ��
��v �
����S�(�'�F�$�ӌ˻��**�iwI�I���VT��ɒ�W�<'�@�i4Y�.�U�$i0>|xx2����(�4�.���B�k�9DҀ)b~S����΃C�%I��'��TkaKE����R4��� ?�5�x��	|�K24���f�]�!\�f\����.)17��.��Z-�[�0���=�`�]��w!�GҎ�Z�"֟�8��T���vo�����l�ר�s´�$I��\�$IZ���8Yv!��p�N�R�<���
p��x/ݍ<O�Z��
�I��{� O��.)�N�0uH������@7I��9�"IPI���W��{�)O������p�%�����^��~��=�$y"�R$I��}x�Lم(:��ǀ�+�)� ���� �v� ?�,�Y��kE�D�b�3�^�ף[�賂�<��K�%��f̵I�Cs�*�&�q���$IB!ɫI�@z(���܋q��WR/���p�ԋ�s����u�$�������K�Eq�?��K��|�����n��
��%���n�
c�]1�p�ڢ��B����-��1�&)E�u�0�87��?���H��(��`���;��se,�X����CR��K��"N��ڳ�=�K����  xr���� ��Wr-�y�����Gh93����PIej pWL��P�tVJ�A�]��K�A��ɕd����1�.I�$IL;�j܋N �Tm��c�GR|��inn.�S{bb�h��H����p����%ע���t�o�-����sn�}8@7�~p5p=���2��pW>���=W����n�]Rb�W1T*i���-��$Iv�O5��A�$�WҞ�2;;�s5�ewI1���Kl�H�O�6�~�~���I;��w��B�$I��e�!�? ��\��������Ԑ� �χ�%�@���n�W ��kT���.@� ͸*.��L�0Y���9Ds�^R����|�\�6z\�$����w�K3��粃��^b[��I��{_�٤ѨN���s�$I�ȹI�����jم(J?�"6ր
�D�O�;��B7��f����~8$�U��yUB$I�{U�nJ�A�{lYb�MR��W��jր{��2%Iyxxq�A�WF��b�zx�FIՖ���݇�΁k��wI����wr�_n)������	TkqT�A�i೧_����~�0�B����T8�B�$�Ҍ[C��ҵZ�ܯQ�y����|҃�$Š���vٕG����R����i�����8�tdd�B�r�K�%���6�]���p?���l�qvp�$���r�C��kQ|^��:�dɵHQ
0|��kQM��ի�+���������pW�$ٞ&|Y��+0�))1o��b�TR��ؤ�n��t:Q�/϶��ˎ<�$�iC�sss�Y�	!0<<�k���`��/�{fl�H�O���vJp!|=�R$IR���L���U%ע��|x�LɵH�`�����ng��<��}���:��*�B�Vے�ahlk�("�sgfIq��K��$�R�\��np�$)���833S�P���wI�j6����h�T�.�y�o�p�]���%��.IҺ�$�2�A�kJ�E���+���̰L�w���vy߿��>�b��w�*Ā���$��4㪶p�j�r��wI��pO��Q���j�h6�e��Z�٤�hd�op�$�]�$��gX<y�Cp�����SSSe����p��K����tr&V��6i;��%IZ�/ǐ���b���ہ�J�EZ�L}�u���9�����.���0�XlJ3���3�.���;��]R/E�u���+��txx8����y�"ILI�|%����(�=/������%����Q�7l�Pv	�"W�ܦj�6i翝Nǀ�$I��Q�����J�E��s������Z���8��9���n�����{�����;��N*��Ag�]�Hp�bw;K��wIU�f��e���]��w�x�;��}��'����NOOPQ�p��X�ī*�T�"N��ڽ(��wddĀ�$I��q�]����Z��O����R$�-�4���׊�n�}!�����tЍ�Y�zg�]Q!lN�b�"$�����$�R�}��3Ώ�����o|�{�s2�z$I�A�G���g*"&��b	���]R/E�m�v/���I3l��ѣO�]�$I*�	��� �Rr-��6�]����F$UL�ct_��Ɛ����.y��e��m��^1�����F��2��K�ܽ�K�E�Y�.CCC; ~�
�3����4b	�W�k���1��垘V����>�1��$�O���pcɵ(>c�� ��/�")/f�'N�zJ ��o9�9�ǭ��'(�wE!I�ͽ�T�{;@�����wI��p�&�;����̶y�^�oΧIҠ
!<���h����;@��th�Z4.�JZY,��uM�T�"�z���J������$I�z�n'����J�E�~�n��*�I� O�~�I�����z�M�0�?��M��l�������_ͫ7���������b�����g8TR/1wI��6Iqp���5̑w�Q�$i�%I�`�qU�朙�a||<��H��X��!)^)��k�l63o�/���l�&X!��(G�$�k
��ݺ_^r-�O �=�gx?A7�*Ik����-�ZIw����ߎM�F7,���!���et7��v��@?N7ho�]q!l���J�V�����6*�X1o�����8��}ek�#��X*I�|%͠��ټ��"y�$U_,�򱱱ރ$���z���J���t:�%I������^r-��{�	���VɵHR*�� ����M�)
I���ccQ�UIIZ�����.aEvp��KQs�*��ְ��ZO�%I��h4�e�����7�U-�/�x�:�8�BR�p?���t�qvp�$i�L�~��B���>ϓ$����ѳ�d�Eum�ۅ\GRu�|-�^)����,�����J�$��[���'�������TjCY�Vcxx����`�]R/�:��.��g���L;��<�$Iљ��+�E�u�o�̒D�vR�}�CN�����5t�,]�V�C_�z�;�q>��WJ����:U�e=#�`�]�����6`~~�O����u�o�������Y����<_�����C�stt��$��w��
'I;v�G}������$I�ȹ,I��Y�;�_�Pr-�ӭ�� ��Vn)�T��%���4���sss=�Uu=��{w�N����K������KXQ���U�\��'J�a�\~:F��^}��!�~�i�z�)��6[�la���l�_S����i��$�z����p�'>ؽ]R�po�Z<��<�����,��W��S7l����$IL��w�|Wɵ(N� �����Z$��U�����i�U5 Y��r�:j�]R/�1��&Iű��ʲ��$1�.I�E�Ki6�����S�B4&''����+��67nd߾}�ر#�S�;He�]R6l(5�>>>^ڵ%UG���N� 8u�>� �<�!�������S�g%���_���$�"�� ���Z����_|��Z$�p��T�8�b�E��$U���p�%����wI�)j�S��Y�!��ڝI�օN��4�KW���v�����o��o梋.⢋.�w����*3�*�:FGG9~�xi׏�k������<���g��{5nI���ԛ��晾)I����� �[r-��V����~��R$�X�U�Z��9M�*���n��,iE1wp��6Iq0ྲ5l2�"I�E�Kiƥ���h4h��9r��z�f��޽{ٷo�yՙU�A���L�z+�k���X�חT�-�~��	��կr��	��:!�L��R�{_s��$i=i�O7���kQ���_����ߕ\�$ƀ�J�j�6�	�T��oQuw:�V444Tv	+2�.��4�!�����5���8�[���?~�oݺ�E��Ƶl\���t:}�Q~�a���سg����}�Zޡҹ��\�_��`�]R�:����^��{��O?�C=����FwZ��1��������$i=� ? L?Zr-�S ���I��IZ���t�Zmc�qy�����n�ۆD%��^�S��난E��{Iqh�Z�\���ͬ5'I2�S)�����;����|������]��!1q�t�;�И&�@B.���^fܫI��T��!@�E�D���4!a��	d��NHl�x��NM.�&� �4�������GQ��9:{����j����ߟe��ֻ���nq}}}��G�^��ޱ�q����庮�^����~%�IO;�{�)��N� 6� ���{�q�N{3�1==�.(��m8ԾT=s��Z:� ����Z��~�� �z�r�yIl	`S#��0H�s����:<�H$���='��U �H$By� �`=~]�Z���o�v�7���Z  �%Yk�HZ3��ʟ뵰{��{*��-�ܢ�o��ecx*%�������4�L��;��������P,�1���B�,�4�p  �YI�Z���p-�wJ�)��r� ��^��Ѧ��b1_�	ch@��R)
�[��� ��h��YQ�7��; �Kg$�}�������V�����ٳg��ޮW��Uڵk׆�Kw a���(��??�U(t��yMLL��I���Z[�s�O
   Qg%�B��P�� ��$�%�����Im�B����_��V�+�կ ���iMMM]�����z��ω�b:� ��sf� O=�,7*�H�T*�̙3*������wܡ;v4u�x<�Y��rY���qO�`s��{&�����J�mJ��.^����I��8��w��庎��;  X���9I�p-�����|3�Z ���#���tp�����^MTC� �Ắ/��Ql4����p x�u�3Ƙ5��#�T"�P�X��ӧU�T��եW���joo��mmm������R��t:���D_���^غJ����odn�R�������ַP���<��;  X�ok����t!�}�����>p- �R��:��Wp��;���50Aw k�k���.�i��C� ��q�؅	�US�JE�Z���B<��쬾��o�Z�j��ݺ��;׽H�Ӟ܋�bh_�TJ����gGG��c��b�����Y�3<<���~
��qc�������x\
  �~GҼ��]B�]ҧ����h�� @˰�- ��{�������$�_ �	c`���u@4���/��	� ¤��gZҵ��z�~���l6�'�xB_�����߿��^wN.
��@�c��	�{<���:�Z���i=�����'�;wN�J%���r�������?�u-  `����_��ZL�IM�l\�u���{�V��;��hdW��:� �j��ǉj�&i x�Z��1�Ƶ�)�ˡI��,��ХK���d���ڹs��1^�.U*�<=?��!��h~~��q���}@��p/��:w�FGG�8N(���9_C�v  ШHr%���A��G�-��4p- �!��mXC��B'��+��aQ]  �?a���Jյ��-̯��_�l��D .�7� ��0Ɯ��济)�ˡ]�[.�u��i���={��կ~��݋������411�����������6���˪T*r'Ի���L��;  h��k���]B������\ 4��;g�-�ӽ���ڢ����0��X�p�#�e��l���E��� x��z�}:c�b��&&&���{~?Bw ��z��j:::@�x}�t�ĉ�f)�x¬��c̠�  ���$�K��$�K�j^'�)-�ܟ� hJ�g ��c�z���~�7y
`=a���& �122�[�¨�(��"Gkm��R  �$9��n�=J��c����B�� �T'u:�XK�RQ�R�<��G�g[=�4��� �F|XүJr�.�v�������fDk6 ��1�b�]�������v� ��0ykW�\�O<�׾����e��2w�q�� �$�R��Y��f���½�������oH�����j��Z�J$׽�Ů��q���_���X�N����~�s�sgՏG��*v�L��1�!�4�u]���#k튁���V�ܥ���<���α����U�TT{���V:�v�����x�/J��Jeů�
� ���S-tp������iI=Z�^�� ���Yk��������RQ]  �?a���& �;y�N�8!ɟ{@c�o�[���S� �$�СC׎9��Ե�1Q���:PU,�Am*˃�5��K����}|5������F�7�/6X�z�j׫y����.}m�"��u��*�����{���Y+�,�e��Ղ�˭�^~L=��Xk����.��C��Y�5��5�u_��j��bp��^�����9O��kQ��^�  ���H*K�3I�Y��%}H��%��� �3����\��TT;�p��(�L��zA��R�JEO>���\�r�Ǽ��B��O�yQ  ˼ 鍫�X.�e��LP��{>�_5Խ������[����2�\��@�mma�1fŏ��U;_�����������x+�f��p����}̰Y`��k����ޯ��k׳��,�/���k��_����������Խ]����v��R  ����I�K�����#�;%�S�X�� ������9�S^�s�R��X,F.|�W7�0V�W[[[���������������x���"w�Y���:�q:� �pZkܥ���Q	u{ğ��Ӷm�<h�J]���4<_�/�׎Y��>�_w\-��4�_{��y�C�Ajkk�}�0�k�r�,c�*������p���k�õ�i�cK_��sk�����o�/@Z����D"q��R  ���w�b��ꥷ�j~P��%�]ҋ� k"�����;W��B���Q&��e��v�௶�6�r�i�K��$]�xQǎ[1,So׫���T�ܭ�Y�J `����zs=�R)2�z3l����bGl ����wؾ��]�j��b��旾�4$���������
���i�b1_C��u�_0_)t^������n�0������K��KY �F�P�\Vy���t�  ���$%���hL�!(�!阤�����k�UpG����� �P(h���W�Z�DB�D��pV�TR�Z�S�5���Z�[[�P��O?����U��#�b���ؘ��N��j��G�0Ƅg� `3;��~-bk�ä�Z%���.�������RX��O�Ӛ���t��N�<y]h�<C7 ��u =j� �Ͻv��w�M  ��'$�K��$�c-��>-�?I�@�� ���#pƘ\��S�|��j���d|	���_�]wݥ��O�]~�*Q����?�ϟ�s�=���~�߮^��|>��R���%�\.OyP
  ױ֞Z��g��~����| ѰV�����fgg}@�43?�(�u#s�T�}�1fЇR  ���I��)I�y�� �$�_ҫ$����[ �Y4f��Yk����$���P\,�����C��ի�� ���ڂ.�:tp��\.�/}�Kz����K�tp����⋾��*M,��7�|3w ��:tM��Z��s^w%����&���G�k2�`LMy?����X+T*��j���P  �ھ(��%�j��I�H�t! �w����X��_m?����rY_���t����L��O���x\�d2�2 �d~~^�<�~�a����w���ᷳg�FjA���|��2���  �^��b��W�G��(݃ ��8�/�!�`=�e�u��jZTv�i�w"��T    IDAT��:   ^򘤟�4t!���$=!黂. j�#p�J��n��G��Z�����Z�:uJ?��r��� ���ۃ.aQ&�nh�VP,��o}K����t�ܹ��yݡ�v�$-<,}��=����7��  Vqj���n~����c��s� ֓J�|�W�J���FƘk�  P�7K��D«$=%�]A w����Դ��Z���DsQa&������-���K_��Ξ=��� �)L��0u��z�|^'O��g>��>}�頺��%i``@�.]�u�f5p��{T
  /c�Y������J111�X,��8 �+�k���D���^�{~�Y��i��  ���!�G%տ�2��I��~ILXw���ϕ4RϱQ����|�v��Db�Rѱc����kr���V�Py���h���1=�����?�'Nl8���cǎinn��q�轱�8<< �i����N/Q�G�Z�d2��8 �+��{T"����/�D�z��<s4  �o�J�!I�$�zI��yI��`#��������Hv�)�˾u�X��䤾��/��k��*���bJ�RA�!)\a{ S,u��Y}�_�?��?���_��n��A�#-<���W���]�w�u�� �&��p�BP�\.�6�|����Q�P�}L �266��8Q��pw]��;  ���,ۡ~o�tL�w]����;B�Z[W��Z�[7�V����e��r����^���gu�ܹ�� DOX��a�@s��.]��G}T��ԧt��1�r����G���!�����Gu�lff���1� ����{���:&��$)���6��Ԕoc�?v].�s� ��H$Z>��r��9I�V�u/�lkk#T  ��V��HI���w]����;¢��F�<A+
���{�c��y=��3z衇40�=+��ttt]�$�@����^�#�<�O~���׿���A��p����q}��_��J��p��Z��S ���1kvq���e��w��������Y��ܜ�c��D"��xa_t��������Y�  �tV�]�.]"�C��$�_��p�%� $��fG�����t�7zYNK�:uJ�jU�d�׮_�����c�=���.}�w~�n��6�[@{{{�%H"����V333��ȈFFF|��G�}=z�G��7�I�T*�r5�C� ~;%�߮�b�\��֗� ��s.�\.+�J�n�@8�(�T*)�H�\.�>6���!U>�׶m�|�\��~&
  ��Z���UIw\��Hz���C�ݒƂ-�V@�aQw�l6�e-533�s��IR(�5�\NO>��N�<�׾�������sy��r��{�DGX:��%h��V�����G�JESSS���T6�U.�S6��s�a�z������_�����7�fqN3[�c� |e�=���*��J&�~�ԐR��{��P(�:�蘝�d�x<N���c48�oN;�J4pg�=  W%���G$�&�Zo����'�D�� ��H!,.�{`3a� T*=���[��ҳ�n��ggg��3���g���߮;�C;v�hQuX�u]�����J%U*���ŷ�b�Ղ����&K]�m(���}Ƙ�0A<�1F�XL�XL�%	9��D"�D"����dR�x\�x|���dr���WX�a	�be�JE�Ri1Գ�ZT�V�Y���Ţ�o?ȩT*r]W��.֗^�ja�fԮMK%�Ic�8�b���6�q�����k��1F�Tj��k�}N�;���Z�|>�����?��󚛛��̌fff6|�?��Db�~m-SSSz衇������馛<�k=���b1�  _YkO���T*�6���)288���'*�� ��t:��¼J�������+��G�c�%�  �dH!�/Kz]�� :^%�iI=��,�Z lb�
Ƙs������<��5�|�IMNN.��Gط�pV=*��Ν;�s�Ω��K��r�n��6uvv����U�ZU�P����uo�����uo��Rx��a�z'^Q�'	%�I�R)%	�R)��i��i�R���3�ݚ}��{:������.��]�jפb��r��R���ئT*��g����%�j���k��ڢ�Z���J�R���_��痆�	ϗ��� z���..��-HX��|>�����#t�����)�z��Gu�w�{��{]��D��t�}�M8p��r  XQ&�9](\I���sW� �%���*�Jy�{:��J$�up�u@p��W���	m�����8� @،j�+��$�!�R!iI*�%����`���,C(���9r$+�{�c���C�ݫZ�ꩧ�ҕ+W���H��]�\.�\.�'N���[7�x�n��&�ܹsKu�.����_�S�[���y>/���|�b��R��2��2����ڔN�߶��+��,�Gќ����K`�LXk����,�6��Q6��뺋 �?��ܣ�����}����M��Ƙ�� lj���?z��Ek���ߥ��|`�}^�� �� ����1�:�]�z5��gff�gϞ����n���a��  hFVҏIzX������[һ%�� �w��yչ0��j�޽�Ӹb���{Lccc/{͏pa�RQ,����lV�lV�O�V"��޽{�k�.�ٳG��ݑ��\����)�Ͽ,�^�{�Z��-�Z�.�?XK,S[[������ޮ�������d<��ummmr'��s�ȇ]�R��ܜfgg5??���������_ HawMLL�_����}��|�bG~?Xk5==���{Q  ����j�=���XL�2�/_�+^�
��,
�z022�[o��k�E�tZsss�������}��@�_M#��ƘAK  ؈����YI?p-���KzV����k��D/�������r���t�رU��~��|�P.�500���I��8ڶm������ե�۷���S����]�U�PP>�W�P����� {�P��qU�U���hfff�c2��:::��ٹ���'�;@��q������D��&��/~/���jzzz1��N�����|��G���ܹs��^�:�~���p333��⻋^� �z�1'���\��0���r��/���+�N+��V�p	�T(�L&�� ���E�-599�m۶���{���C^�  ���~R�g$�%�Z-��>&�G$�/)|� "��;��\�NNNzYGCfgg��Ϯ�c�PP<�4�d�u���V�p��d��ޮT*�L&��];��q%�ŷ�%���&����[�ZU�RQ�TR�\V�TZ�S.�U,U*�x���y���wTH�R���m۶i���ڶm�:;;�L�������r����)MOO/�������L��Sa�G�������멧�ҩS���׾Vw�q��Y'&&��4:� Q�VO�� �u]U��P�.699x�♙�H��+�o�)L!R �J$�x1�5��ňa�cn䙔���;  �y-��?!��ׂ�y���t��K�� �xJ�0y����ǽ��.���:y�.]�Tw���O�����jjAc ,�Ţ���ˮ%�������K۶m[�wuum�`AGG�FGG�)
�A�\.�f_mg �kE�|-�i����g�ы/��׼�5����=	�5p7��� �x<~|�y�b����6�*Z[�R	�+�$]�|Y�y�k|Y� �R�Ԛ���P(:>��0Ƅ�i���D��ܳ���k�  �*EI�!w4�����s��p- "ls��i/mY]ױ���r]Wku �V###:w���״��yp�1�Z��ή�ټ��C������RWW��������VA̃#\���̌���455���	MNN����׋�R��'睚���O?�o}�[z��_�W��Ujooo���Y�Y�V	� q���KG����m�cJ�Rh��h ��B? ��.�]��}��]��ct�ʕ�ː�p���f���t)���>s�}���*  @c���)�%�L�� zvK������&<4��;Bcrr�lwwwQҺI�J����)_&��ժFFF400������d+{�0<�6�Z���ի����ھ}�v�ء���ŷ~/�iF��0u�YK�\���&''511�\.�����8h���6�L���)�bQ'O�ԩS��w�^���+^��
�LwI� �0��Ç�4���jǄ�K���܊��r��y�~����lqSSSA�����~��tr��t:��njj]�ð�j���^�  ����p�K�?�Z=��ߑ�o%����`�5��������r�ȑ3�^_����]�������4::����m��u蕀;�J�����낆�㨳�S;v��Ν;C�a�d_�����N�C����f���0��䤦�����K�_�"k����5<<�x<��{�ꦛn�+^�
����5;;�L�d�СCl# �1渤U�R��jVf����X�e\�X,*�H4��&��t�ҥ�ː$� еkׂ.�:��j||\7�pC�u�J�F�	� �(��z%$�7�ZMo������>p- "$|�2lu'Ug�}||\w�qǆ+
���Q.�S.����r�\������t,ck @��jjjJSSS��_X|Z��ٳG�v��Ν;�}��@���{��[k5==���	���ktt�0;2�dRsssA��r�JE���ԱcǴk�.�ٳg��z��f��[k�� �1��Z��a��������\��}��,��t:�kS�S2��)����ٳA��2���joo����nD��   ���_�4!��ׂh�.��%�MүJ�� Q@��b�9Yo�py��\.�Z+�uU.�U�V���U,U(T,ߟ����̌�[`����1��1 4fi��ܹs��ڵK�w�֮]��c�_��pb�b����q���kllL�-f�^�|#)��@�S��ؘN�>-c�:;;��ݭ��nuvv���M���J&���bM��a�? @Ў��bmN'�9�Z�0����-��Bw`���ϳ�k׮i׮]\��-�������X��ȈR����d �7��qī:   |�I3�>(���y،~Aҿ��3�N\��#���y��GFF�я~4R�vggg�����	:zѐ��u��U]�zU���;w��޽{�{�n�޽{�.��L&�H$|_�#���=��/vg�v횲�l�~^ �gў�Q�]bzzZ�/_^�fv�־���  ؈b�x2�L�Z�W�\$�T*�42�����u�m��c��8��K�.]�u�[��t:�Ԃ{������!�z뭁,�lp��p�x  ��C��$����9�����_�t$�Z �?d*�T�X�P��֝��uk�R��j����nO��j5R_ �ժFGG5::*i�!�;�{�n�ٳG{��U"�h��f�-=g�����FGG522���Q��ζ| ��z�^,�d8���IƘ3� @������=z�����Վ�T*�ܫժ���B�, ���q���N�C�(wppP�w�� >rg�E�aR*�t��5�۷��gd��h���   ?��:�LR:�ZMiI�%���� i2�r �w�������=za��KU�UO;{!�Jyz��:�h-�u5>>���q�9sF�uwwk߾}���{�n�b�����ـ{�X����b���I~�6�F6�����[�k6|W�V	� g�=.i���w�r]W��8{�������`゘�YO6��-�ܢ|>t) |�Ǖ��.�.����7��븍ܟp  ��g%�M�g$�����wH���~^���@�D+�-�u�cƘ��Q�Iwu Ͱ�jrrR���:}������٣n�A7�p����>ggg���o���N����𰆇���f#�3 @���T�J�"k�綵��mu-  4Ḥw����?���T�X�m̍*�˚��V:MC,`+H��:w�\�e�hff&rMg 4'�J�̙h�������8ڳg�oc6Ҥ�q�QK  �W%����Kj< ,�E�K�M���m'4 ��,$B��I?Sϱa�Bz%^w$#�	l�JECCC����s߾}��曵o�>%�u�D��q��;�����ڵk��А�ݜ���!����&�}/�߿�յ  �(k�sk-���~�Z�jhh(�݇�\��׽�u�/�b��y���~}�w}W�h\.���l.���ڻw��M�*�JC�5�r����   �qIo��EI�����;�~B�/Jz!�r �w�����N8Yke��TW���Yc<{@a�U"��}ko �*
���W����ݻu�7ꦛnZ�cz���9���k�jUccc��ࠦ��}�@X��0��JMܣ�j �i����Z��J��eF:�y��E�z뭑��P�d2�^�3\k-� `H��:{���%��ŉ���U.�u�M7�:�
^m"���;  ج���o$}Y��ׂh{���$�I�}I��~�e�#t�ĳ�J�*������F�g�PP{{�fgg=#����\���ȈFFF��sϩ��C7�t�n��f�ٳgqB۶m�׶<l_�T4<<�+W�h``�k I��E��i3$�1� ���>|x��g�׽�:??�k׮�Z�z:�2��'�nk�w�ℳ�����U*�j�� ���6��/\��;３y`�J��z���f<��@�Ryf��Í���z�������\S���\OOOѓB   ��IwI���;�і��~I?*�IW�-@P�[�4���5��ݢ��N���d2��?J�xovvV/���y�}�S��O<�+W�x~-Zɶm�T,u��E=����'>��{L���<������n۰f�y]�%� �q�[�j���nw�Z���i``���eI�����gk��ė/_&�lR�dҏ��V�TB���q488�ǿ�8pತ/)��|���٬'�opN{ē"   �岤�t"�B�)������t! �A��d��F�zY�'��H��Z`��Ţ������}M�����N�}nnN���'��Ojpp0��� D_6{���;  L���ܥ�wq�:д�Y�q~�����%����!I�o� �?�����^�X�L��g�r6�J����	����N�?$I����r�ڂ�����_c������  �kXқ$=p��K���OH�p- |F�au�����:TU*�<=?��!�N[QyH X^/`�Bw뺮�{� � _�JE###�|���s$Ƙ�Ƙ������}���B�ƩV��p႒�d�N	 `mmm:�|�e��Z�" J$�\��1��������x�^k�������ҥKkٳE:�  �*+�G%=t!�4�%锤�] �pG(5��]�^���PU�X��� 6�w|�� ��um�/:t(��Z  � O��jbbB�������й�a�y2�}_OO������\���V+Ǜ����А��x+O  ����Dn���ի�d2A��2��N�>��P�|�������w�}�Ƙ_���E��8���_�lv�����oh0  ���B������W�g$}XRg�� �w����ۏK���A�&���z��H� l~Q�^F>����^ߋ����/� �����W{�ـ{�T��ؘ.^�����@~���]�R����o��R.�{P�c�wrrR��ӑ��p�d2�k׮]FS^|�Ev� "��p{�u�_5Ƽ�f�����Ƙ?�i��K��qdd���Q�ܿc��  ����wH�xЅ`�0��KzA�O\ ����t�=��1'�=>j�%�U�T������~pP��wnX�n�Z��V� �F�fZuV#;LU*�r9]�rE�.]jI�&U%�?��x`�Uz}}}���^ݫZf``@333��b�<- ���i�9s&�2�V(4=���% !W�ot'�:�ޡC�V��MNN���g�(��u]MMM����P.�k�k��׍�;  تJ�~Vҟ]6�%}Z�'v\ �pGhYk�Ċb���`U"���� 6���Q�^�W*��t1L���҆��tp ������^[k�[�Z��ܜ&&&t��e]�xQ���*
��Yk��8?��"    IDAT���[w��C�]�t�յ*��*���� <��588�W��3W�\��
A�LF�N���d�y6���������+U��'i��V0??���Q]�xQ�/_����fggW�Gu]��9,�qV��  `�Jz��?�l:�tꥷ 6�-c̱z���F�+����� ���`k�:��=�����K� :ƘUw)����󚙙Q6���ؘ�����߯.hppP*�~����c������_m�{{{�\ҟ�����a���2"���pg38u�2�L�e �S*�҉'����u�g���J���ZkZҚ;�x�X,jrr�{с����hbbBSSS���j���@��   !b%�GI�t!�t�j���'^�;�M"z�l�ܥ�u�:\������;��x�u4��&rN<x��յ  �Q���W{�P(��ի�v���Ɣ�f��k���l6�����!�l6{���[X�$i||\gϞ%d
D��8�|�r�e���VgΜQ:�� k��b*�J:y�_���1�=8[�'<x��-�B�Z�j~~^SSS�����Ȉ���9�[�T��   lr�Y�=������]�^��n 6��;�eLLL��4S��Q��n�����Һ�0 �wQ�r����G������E�Ǎ1ѺA l	�x�|�5l���w����Ǿ���r���W�־Kҕ֔�m�bQǏW,���>`+H&�:s�L�e�\�T҅�!��d4<<�K�.�9������]��t����i!��Y�?���v�  ����nI������%�#��tK�� � �p ����\I��{|�{���'>Q�V��׉�����c���  Z����&���Q�گJz]oo�?��q]��<��9s����L"�ЩS��.�3sss:�<!w D��\����Ǖ�f��s�����f?����w%}����Z���k   �OKz������VI'%�+2�@d��f�9V�Q��.y�*���b�� �A��z�܅&j�ۥ���Z� �0;t�7�������������:����nI�V�[�ffft��q���6V�>}:J��������ٳ,��L&�8�Ξ=���}�D�j���}��MOcl6��O�߶��@8��ɠk   ��J�K�PЅ`S�&�%��}��	�j���p��r���h{{����F5��u���{v�uo����md�(  ~3��c�5��ik�����5�x6�t����[kA�g+�u��	MMM)�N+�Hx5��R)�r9�={6��ɤ�c
?~\�d2�������b�d2�T*:s�^x��˞��[����t��x���R�����۷1ӊ�r|rr�A  b'�r?t!ش�Wғ�>"i{�� h@��Rb��3�����A<�   hV"�P�P���QUXk��R��� �V�V�]�:��~+���u���������������㌌��ĉ:}������8���2��R���D$ae�Q&�ѹs�4<<H�DB{��	dlI:u�fff�Eh�x<�d2���;��(�N����Y�;wNǏ�ŋ��M�k�L�-���j�	�������=���U������}}}�z�	  �~I�Fҷ�.��#�=�^�􋒢��آ����;|���1���X,�T^��n���� ��b�����x\�xܷ� D����522�����b��g�o5�uU*����'z{{���  �*�Zs���3����|�Z{��`�rG�}���c�2A�_�ŔJ��N��L&�L&�H$�����8��Y\@X[�g�U�R�\
�mmm���h�u�ܹS۶mӵk�<��^�1Fw�y�b���ݤ�0����b2����3�u]U�UU�UU*��e�E��e���@���Z�p&�y����=۞��ѣ���wE�������}_�E   DH�����������{%�	� k a�(������(><�M^z!�_  �uy��L�:�o��ڱV� @�c�#G~O�_]�W���v����YDOO��>�Vc����+�:�ժ���5?�\>my@>�H(�L��_:7�4(_���(ب�����!�={6�r�����)I���
���V/���b��n��6utt�P(�o�P��U�K���ҟ_��z�\^�S(T*����7����r��<x���hzzz>�����8��H��r�����U.�����   ��YI?)�IzW��`s{���Z�)�7%�Z�pGS���b��K^����  `)���t�(��{Dk�7Z\
  -�N�?Z(~]�k.eR��m۶��s�=��H9x��??���op�$�>�z��р�R��p*�R<���|�1f18o��㼼�����:k*O�x�P-x�Q���T�^�֪\.+��jxx8T������߃2����t�s��jU.\�$��i�p����T,�.$\�ڂ�V���wX[�_�{��<|��u_�-��1}i��ڟb���P��K����ޏ�5�C�>�����q����F��m@�Z�[�à  �����[҇$�'�Z��%$�haQ���
� �E+�-������%�L�䁆_���F�s�)�Y�͚�y �)��^#j� X�Ν;588�����g��B���X,v��o	 �:>�:c�S�2~�m�u��x����ެ����#�H[�P���_
���$�)�HH�b����ڜc��X,��P���+���W�Z@5��5/�Z��^��>�u�U?O�������=�$�I�x��}��EXU4c�J�V}=�L��@���ne��9����F��ֻ�l�Zג�,��T���kZ-X^�VU*�$y�<���~=����� ���������B�Ŏ jX�*�\�}ߡC�.]  �&`$�����l���^I���K�#�|���������'+����v�ܩ�9vQ�2� ¤��M�����{�@Bظ��� �AS�lvG__��[ ��Ç�����A}���J�ox���Ӵ!�R�K�t- ���}����;P6�U.��* �Ȝ1�&''��a��������WI?���~;!�3�X�/8p9��  6�{$��$��CI҇���b:�Z�-��;B�Zk�=:!�����Y�#J�x�q��o����g�m��E,S�X�l�_���ju��kx����-��  /9r�.I'�fN��tL�?9��������?��?����󋒢�u!�@�رC۷o_�������� Ѐ�1�Oc�������.f�������^��EI��.H:m�9&驞���  ��~Lݵ;�.[�5I}��B�5 wD�ѣG��Z��z��Zx�����ު���� �����.{�l4�N{z�V��.?������V� ��>򑏴
�I���I����tJҀ�v�3�nVRnjj�B___Sۢ���Ç_g�����]�pڶm�v�ܹ�1��jhh��E� ��YIu]��:t)�b�q�ȑ[�1?(�fkm����v�g��1�T$�.L�/�ڢ��듕Je�q��B��}���7��   �y���K�t!�R��tH�?]�pG$>|�Ac��z�O�R2&��^�o�����*� �bϞ=�r�g��"�R�$�m|�oc�O���|���  ��ѣG������ZI����l�Z{�q��j�z�����������6G�����ƘwJ��V� <��ѡݻw�ul�\���!w ky�Z���b��	w   $^)�aI��l9��ԣ�]� �$	`lyG��ek�_�{|2���Dc�f���tZ�_� ���;��رc����<#Jܛ�>��Db׽�ޛ��&  >���8�/���vc�%ł�	@0��������縮���a�E��1����Jz�Z�ȡC��]   ����>+�_]����K�m-4d�1Ç���L��G)@�lw�F�ݻWSS[���u
_ǋ������fgg=#*��Xk���������  DÃ>����b��~-t��I������ǵ{���Zk���455E�`󱒲���ڬ1f��'��c��~�q�W��<�@>�z  �z�K�����lIC�������m���H�!�ęJ�bU碌(M��Qk:�&�  B���C��㞏c��D�}�oe   Z:���ɗ�H�>��ǆ��w����Z�#����0�t[kwH�!i�c/��J1o���8ڶm��o߾��L�1���V[[�r�����[X%�VY�S�1���AI�z)��8N�Z�u]7�ǳ�J%�ҽ   ��I�?%����ׂ��FI)齒�$}"�j�M,���%G��,�z�5�(�Jy\Qk��=y߾}�f��� z�� v�ޭ�W�z>N"�P,�|���T*�T*�|�����~���  �����s�^/}{���@���WZ<��@T%	uvv���sC����EMOOk~~��G����3t������:�q�[��>�'R   �hx���]���$���ǂ.�lH�!J�W���<L����q%�IU�U_�A\+�r}�/��Q�r�@�tp  -U�-ح���-�4(�4$�J�.�R�W��+k�������Z����'*�r@�9��t:�T*�L&�yc�T*�ݻw�Z�|>�|>�b��b���@cd���8rg��X,��k����^�f����g�pz#��Ea:    $> iBҟ�,$��FI�J���ߔt*�j�M��:�䌤��{p=�0��W�r��={�hbb� Dw a�8�o�(Q�>���roo�V�  �
�C�����۶m{媟��J���ǖ���]��=`�㒮�/m�9�6:�Ys��D"ђn�Xl�<�JE�R��s��,��v���b��Be�Q[[����$-�;��6U�TT�VU�T�����b�V�>Wo�Q��q�X�o�&�L.�ˋ���3�ڿI+�]�ok�ז�,��}i���juj�.�a6   lB.钤OJ�l)���.�m����ߐt!�r��#��Ȱ֞idR�����خ E8 �r����e����Vҽ  lz������׿�����/�˒B�K�/]�]ug�Zx��V�O-��J�ӊ�מ�wG�Db���z��!��^M<_u��d2����ߚJ�T.�599��1~����ŋ�.�7�%��~�E�j�v_��(��H��b�z��3nл���}��ǖ_V
����ɓ�"    `=_�t���K�5�Z�u9��-�%���ߑ4hE@�pGdc�4r|B�~NBONN�q��� x�� �����j5���j�Zi����   @�.t�V��۷oW:��uL �Y-��t!     �W�$}���J�Wׂ�-!�=�~N����{���� Z:#2��j#Ǉ=��w}sssھ�]x |[PasB� j�1�w_ܬ���گ��          j�Iz���\ I��'邤>I]�VDwDơC��$�=>��ն%�Rػ��WP!ϰ_�����K���Y�VC}j��l6�}�յ          4'��~7�B����;��Hz���`����;"�c%]���0��`��ccc��.��g �1�2n�Zd�z4y��z___�[�         ��Z��I�w!V֩���W$��7�r�p#��H���7p���lH��%�X,jǎ�� |�� H�DB���������\#�1�{P
         u&�m���.X�CR���Z��� ��#R�1��a����v-�ˁ� <��p I]]]�-�s]7�!w�         @K������5�Z�����7[.�)�tp�x�Ji�뺁�522������A;�*����@�*\��&�����         `�8)�$�`��vG�Òn
� �#Rǹ���a�[kSYk�N��@���[kCw}�;vhbb"�\�tW�V1�<y�=���         �I?(��A�"#�W�EI-�u����;"�Z;���^�Ҕj���FFF�J��.@����� ��k@�R	Ž�R��c���G�       �?{�'�Y����O��]�ժ˶��C5-�1�)R@��L�b��C�'���PlH�`LOO�KH(!زqlzq�-W���Ҷٙ9�~����JVٕv��y�^�5��Υ�ݣ���|  @����BI�t8�����vāoHz�$�4� w�c���ܾ�
K�0��.�c�������f���z� ������������3�Ķ��        �E��F$�TGJF�{��/H�K����q�ơ������[��Ǳ��طo�r��� h���i��� ��\.�T���i��E�~w_�n�ˑ         hs��t�����Y�> �~�v�X�2���R����� �R�J��i�Su�JE�c p��G�0E@����j��E���2����_{�K^�C         �����'J��� ����Պ��t��4�2���V�|��cȲ�iJS�۳g����� �Y��7C�@c��ߔ;�dY�tG�Y��]          Z�Ò~Eҿ�,B��m�~"��W�h�i"`�� �k��j�{�1g-䎞������a�UEMY�j�JW�X�R��:
�i��n�,S.�s@���v��G��}�Y�4M���6��e�}��F�         �ܴ��Pm2��EQ�×�����>&�zIc.CK��;ZA�j{I�&&&,�i�q:�3�㦟P|�=�hhhH����� h�f�.�r9��B��y��4M533�:�q�a�l�$I�{�c�z{{e�y��+���A�         �vg%�H�K��%���LI��NI_�t���N'��hk�eY6��ۺ���l%ң��*MS
�@�h��R���<V�X���	�1$Ig�C.f��Z��         K�s�.���u��%m�t��;$m���4p(���Xk\p���rE9�V)��8p@+W�t�2k����&h}�bQ{��uc������鎒t��          @����%}�u�$=A�G$=,���qX8
�h9I�,���h�Vn�۳g�zzz\� ����Ln�m�)�d����J��u�E��*��f�>� nq         hcJz��Ϻ,�I�'駪S{����D�qPpG˱�N.����Q�i�r�T+��i*��]G��,k��S�_,������\�8aQ5��G���9$"         ��fT+_!)v�X
F�Œ�A�I��t���@S������	��,������u���p�2h���uY�5�d '���_{��~;��f܆nw          � שVuXB}�.�t��$�G�N�PpGˉ㸩&�gY�(�ڦ��k�.�\��u K�Z���(���X,jbb��w��K��!۩El��}9s          x��$=Q�w\��FI,��M�<�w��(��]g�KӴ-K�{��a�;�F�4m��{��`Ha�Z�j��:ʒJӴY��S2�|�u         �=,�%}�q`9=A�GT;b�?Iz���i"t$
�h9�J�y��>�=I��/���,�t������ꬵJ��u����u ')��yMLL���,�,S�N��I��z�UW���         @�Hz��?��~�Q�G$m��I�I�V�S%���9(���$I��$��8n�b�|qk||�I�@�k��LdY���V���a�B����1�Q�]�����澐m�����%])         ��~I�6�hwT۩�vIJ���g�2��\h9Y�9ik�i�(�Zf�R��XcccZ�b��( N@�eK^�\n�T���|>�0;��^W�����]w���F�         �1}]�%��� @m�t�j��J���H
\�B������eYC'��i�8��$IGNN�D����1]h%��CN�e-��d���J�Ttŉ,�EQCv�ɲ��_�җv/��   �4:�����'    @zXүH��� ��%m��I�%}Z�ݱD(���T��E��N�C k����$IZn�R��ꡇRoo�����8  ���vu�S�nd    IDATE@��<OCCC:x�J���8Υi�j��������ey`   4�V}o�\<��4     @S�Hz��+%Ug\�t�je�%����%�.C�u��`��J��lܳ,S�s�v
��ڷo��岆����4�4M[��FLBp����T,�s�N��p��D�8����~�<��W�����l>   ��V����$     hr+�i�v�8�V�>n�tP�U����e(����,a��Z�,��_�ڹs������ӣ��q�m@�ֶE9<�2%I� �W��H����ˎ��1��K��d���yǜ8y���Z��s�����<(   �w;�1F���     �f�]I���qI��8��%=v����Vx����%Q���C�)�J���n�=�399���I�r9��R��j��� .�����4����A���GA�T*itt�u��T/��K8Ƙ��^~?�$�J���r��{  �Ǳ��L.�'�˩\.��     p,�^,�*IWK
����y��K�'�V������� ��;Z���ĢF�i�D�eE����3�u>�W>�W'5y�X�M�w��;.,�ÿ#��p�D��o�e��e�i�Y����(j�w�$�+�.y�7��E.���Y�}_Ƙ���������?���v�������?wT��������S���G��G��?Vi�xGzH�DQ�\.�T*�X����Bw����y93  �9Տp�|ZG�     �+郒~ 鳒ָ�4�U���.���K�wI_Um�{{��(��r*�J�:��Z�v�wc�\�?ù�b�����Z���%��e����� Mӹb���=:K��o�r{]�$
���;��1
��Q����TU/��/�K�b��ys������e󯋢h�v��B똚��s�[  `�5�{�(�(���st�f�   �I�U���A�%n� M-'�Y�˵�Mw�/Iߐ�]�wEὣPpG��U�Pq\^4%k��8����F�@���!_ק^
�g6��M��֏��e����^n?����3U�aͭ�3��#yԷ?�����y�����ow�
�4U��:[�T�v�  �5��홙uuu-�H����}
U*�Q 4GN   ��Jz����.���[%����$�J�M���7%��Q.4w����k���19�Y�fT�>���za5��?75y~a~~q^��t�zi��0m���˿�2�(�c��Ȥn����s}��3��;��K�A"�2U�U�iJ	X&���%�   :Q�sC\���*
Ns4���.
�@���M
    �@*iD�w$}ZҠ�4@�Y-i��"I���t�%��&�1�$k�1f�u��$I����0����J�Ƙ����C�u>]����
��էZw����N��\9}���#���v����Sсֱk�.
�   T*������R��|>�����0T>��=-�*�JG��   @[���'H�A�gZ�ZZx�G�	�ߞ]~�ڎ%hQ�5��W�!�"��������'��Y*��R���TJ��$yY$c3y6��L�}d:��U�<z��+�d\�?q��~~�e�C?m�)@|�s�V�`��呾G��z׋��@g�߳�Zcd�[�ô   �Js����]�X�o�d�+�5b]'*���<ϓ���c4��8��B%IB�G���Ւ�jVq+�"�1�ɦI)J��F�ϋ��gl�-��تoTͬ�j�UB��Tb�?���jdHl����=_��7�\g  X&yIWK�R�8��0%�Iߒ�_�˨�DX6�h�*������ �a�X^R�I�
l"/��X�J�3�r^��oU�B`U�BϨ��          ͪev��F�U;Q���r�=0S��J���n��go��  Zݥ�>%i�� @�-�NIߐ�M�
���pT4|�tFF�;��Z���Y�f�s��T��B�t���B���<���:          tk���$�_JǦ*鎩�~w������̗o��[e��   a���Hz�� @��J��j����CI?��Q՛ �`4��֋z�bvfw1�9�<��s
9�Ԯ�,��w������          �SM2�Lf���(�}�T�����-7I���  ��t���%��� �,�t����Vv�s����:w,�������%��>������y��
�p��՛�|�w          ���t�D�s)�u�l�S���:  �Q<Y�g%mv�!���{�<G�Z&ԌqR������S/*�q�9��ނ�nE���+x�G�          �d�M'ɮ��ޱ��Ɖr�7#���nי   ���QI/v�1Œ��cI?��?��ݢ�~�h cAF�^�S���W�ד�.�-���{���          ���Vzh<��5}{�d�w����v�	  `�6I���:�E�$=�Z��g����.HJ�Ek��(���'��C]�_���������          �v6:�D�G��;�|�-�o�^�r
  �+�I���Ǻ`IĪ���t������t�]��Bc������Z�7zQO>���˻`Mo�q��]�          ����4}�@��F|�'��u  б
����:�A ,�i�����Vx@�Ò��{�|�U�F���AFF��zw��Zw�a����`Ӫ��`v           �n�D\}�`�����]o��M��:  �H/��QIî� pꠤ]�v�VzHҾ�e����$YGO��662�5Wx��s
�����6�s>�9           ' �V��E�;ƪ��wg����7��  :ʰ��$���  �^�Z�}���Ic�ˁ#,���T+�;Gٹ����E��|�������n�I�V�닡�k          ���3{�Xt�C*�x��n��u  �Q^!���\Ж�[�U+�W$MK��T�4!)�=��^���G����k��u������K�4 �_����⮾�/���ˇ{���W��u$           :�}c��}��>6��n�V�u  �N��	I�t ��3r٥����wWv�/=e0������           ��J�ݽ������F>}�ݮ�  ��g$�Z��%u9� K��{x��[~k����5}�7��           M�g����O���Om���<  ��'�3��: ,��Mh䢋��3�m+{r��2�{��.?t�	           ,Nf�v���8��䫟p�  ��@ҟ�.��, pR(�7�������.��oۼ2��ނ��           �Ǝ�h�;g�|�S�\�:  hkJ����\�E�ݡw��WWt��oY�lݼ2wJ!�x=           hc;Ƣ��V�⏯�~��,  �m�H�F�6�Ђ�p5��E=g�ۆ{���X�;�;G�          �Ns����Ov����>y�G]g  m�%]/�L�A `1(W7ȵ����W�6�凮�            ���~��:�?{+������:  hK]��.鍒|�Y `A(�/�����v�r�����           ��Y�G����|��?����r�  ����6��\�A �x(�/��[�?m�?Zߟ{�C���S           �/J�~��r�h9{���]�  m� �͒�")�8 ��%2��g�5����5���l�          �	���������񶑑[�y  @�9_��%=�u 8
�'��+��l�7|����3C��           ,��ǣ�wV��-�~��,  ����H�;%�g�C��>oy��Vn����U�1�           ,k������}�ϻ�3���:  h;gH���_v �(�/�{_�����_���xq_��\�           �a��ew>T���}��WI���  ���I�\ҵ�zg 
���Wmy�����sW�/�<e           �����������-���  ���>,i��  :m�c�zۥW��"�?���{��
           �WI��x`��������7D��  ���I+i��  :��#x߶K^{�`�O�X�r�           �H<�|g��{�'n���,  ��tKz��?�8���Pp��b;           h%Qb���_������nP�:  h;H������sPp�tͫ��洕�?���y��K�H���v�_���O���x�9��          :��dmv���뭕��ٻ���!�q�����<����o��  ڎ�t��k%ѳ��:����˟���W�9m07�:�x�����#�`�|�2_��Ne��e^0{ޛ=��_          �1[t�Y&�t�|Z+ϧ��Mk�Y"�&�N��i�2��a&���;J���n��u  Ж%�[ҫE�2��̻^~�O.��c����LG>��y~N&��s�\���2~ �e���y�         ��d��4�Mc�4R������X6��%��i,ɺN�����ʎ;w�?���ܾ�u  Ж~I҇$=�u �������?uE��>nC���Q�tw���充Zy=,��e��ly=t�          Pg�,�-���٥�,�*K"�R�of�Sqt����z�����u  ЖI���g�zg�f:���[�Z<{u�u�Y[xio��\�i7^���+����aA&��
�A�u<          �R�R�D��㊲��,*+�˲I�:!$U�L߸o����#7^�:  h[�H���_w@�h���_^q�<v]�m�=4�O��C��.y���\�2��g           0�Ͳ��{YYTQ����ьl����q~����';�'���7���  ��3%�_��� h}m[p��Wo���+�>oua��,���"{�K~n�О����           m�&�#����hFi����e�k".���g���7�u  ж<I/��>I�g��ڮ�>�uknh��g�|Jqk>���߷d���+�/���u��w)(����d          �dӤVx���VKʪ3J+Ӳ6s�mLWS��{Koz�Ƕ_�:  hk=��(�͒� hAmU ��[~�1k]?v���T���B��|��b�d���          ��ڄ�JIieJie���Iʬt�}�_|����B�Y  @�;C�_H��:�������ykV�M�+>�ζ���_�UP��s]m�J          :���)�i%�)��I�Q�u���]����G;��Xr�  ���%�_���� h-_{��K�=~C�߬��C�Y\0�_����'�ا��'��c          �06K���j��ʔ��l�������_�����]���s�  �=O��$]-i�q M�e�oz�{�썾�]O朗���k�ٻ�{�Nz           8+��ڄ�dfB��8����3�T���ɋF���o��  :�7K�}Iy�Y 4��lF���K~��u������:�r3���{�Vh�ꗟ�j�W           G�j��g&�̌+������TMc���߾o�7]�g]g  �lI��k�� h>-U�~���?��/?~c�Y��R���/t+�WjgB;           Khv�{<}P����J�va��3{�=����o��u  �Q.��nI�t@�h���{_��瞵�|c�`n�u��f�Pa����
�d��u$           :�Mbťq%��Ke��u$'���k�L�����]g  ��&�?�u �D���m�^u�)]��-x��,K�
{�*�h�W          �6g��<Y+�O�)�ʮ5Tf���-]�{��]g  �Hz��?�t��, j�Z�Ȉ��}��ק�Z|��5u�	�}
{����\�           ǑVgO����i�q�Z��{J������K]g  )��
I#�ֺ����m���e����u��ίv��d��.�����[E�          ���U��O�SR�tgYY+}sG�+���W��:  �X]�� �͒g�@MYp�[~�]�(���,'��w+�?��w��0�:           XbYTQ4�O��^eQ�u�ea�t������o(�  �%�I�U���� h��+�ൗ���N���|�5]�c���!����z\�           �V�M�U4�O6�]�YR�J_�Q��7|諿�:  �x�%�]�+%�� e �T%��9��S�~�4U�c0F��!��W+�h�g           4����(�U<}P�u�hIX+}c��?\��_�:  ���$�U�o��;Ж�����7<7��P߹`}񱮳,��X�|�j� t           4�,�jS��V�T]�9i�J��3��?�����  0�TI �
Iy�Q ,%�u��o{�����[S8�u�c3
{�Եz���7+���?}           �	�W�է����ݲY�,���u�NY>��S������nt�  @Ҹ����i������@[p��~�+�}��r?ڴ"��2Ǳ�W���ם�����rב           @�0���R�X��aIRV-I�ns� ���2��3N�4yӝ�~�u  �Y�ݯ��Jz���i" '�Y����_�'��u�pOД���¼
C�Ե�l�z�d|�u           ��?PسB��52^�4����u�E�Ѻ���S7���׾�]��   �S��]�G%e�/��@KrRp��ly�SO�e�;h��T>U]k�V��'c<ב           @1����_���y���l����`�o�Po�u���_���q�  �0��3�'��4�E1�^��W\��7?�_�M�?/,��r�r�k<+           �cY�hr�*�PW\�Y��I�ֻ�g��s7�r�  �VJz��ߓ4�8�hh����_�_:��c�9�i*�^XPa�)�����           ܱV�Ĩ*�T�D��,���������铟��u��  �SJz��+%�v��14l���^}ɋ~������MQ#7~���&u�;[~��r;           p�����J���2%Y�:�1�����������:�Y   ��,�6I%�IgJv��5��~���}��N��BO����c1�Sa�u�?Ga��dh�          �&b���>���H6SZ)�NtL���ugn޸��;����,   �J���K�Y����bT2�4�����Wny�SO-~���7lZ�ф=���p�¾!�k           pT���*�RV-)K��#�1Һ��I�m��[���'��   ,�>+�_%uK:O������^�̳/��}�PO.�z���*�>C��Se��e           �E�P����¢�ʤ�e�#=J���	~}���x��;�:  �"�J����J*I�@R�i"��-��F^~ɦ'�R�k�@���(?�NšS$���           ���4Qy�}�&F]G9�����q��nd���u  ���+镒�@�)�� gYZ�##[s�]���e������O��           ڂ�u�=S=A^�s�Q�\�_5�?��9   NҔ�J�,酒��6�Y�e�����y�������"�b�
�N���ޖl�I6��R�ZY;���R��n�&��M%Y�,����l*k��uGP���Kee��_         ����|��:��x���d|���~ndf��A�ƞ/c�d��c�o;w��&��s�����"N�n������ћ>�:  �z���Jz����,@[[��߾���qzϫ��q�x��֞��w����X�U�Ʋi"�ƵBz��fI�|���M��I�D>[`����L֦s�u          ��?�1~������=_������ْ�_���e|_2��z~X+ӛe��������轵�oMbt*�n�S�8�w7�u�  `�H�IW�6��[�w���v�k/>��C���7�~�[��ϕ�+4|��JY��keu�%R�)�RY�Ji:7a�f��L�RR�<��t          @S3A(?�]+̖��ys��y�kㇵ�h��    IDAT��s��p��1���2��Ο)����������~�/��<�9   ��'�bI�$����m�},��ǿxՖ����ݷ��\�\�*u�9�l�����Y)Kf�Y*��2;{����2޼C�y��M�Mo          �/,(�\�m�ͤ,���L6�������'��</�	ByAN&��n�b�D�]w))���"�6P~�ݓW���or�  `���t��+%mp�hyKRp���{������R<�bVnPaթ�^mKɒHY\������c�$�����Z[;���ݓ����Sp         �ֵ�����G�n��g؞/S�;e�P^����y� \�m�Z��G�Ĩ�$���j��Ǐ����箳   4@Nү�6��Y�8F�	Y��!�wzכֿ/�WoV~��Ʈ��X�,�֦�'���:7�ݦ��M$+/8tں12~�pp           �cd�@G;xx�3�DiT��r�y�'y���B� '/���u�w�@ƨk��rEU���:�z�w���H:�u  ��$�0��%镒^-i9���I��/_��>��F�cb��ן�\�pWꐵJ����Ҹ��1�S���Q4�WIyBY4#�F�i*�L�? x�?�A�|C_�GK�3��           �����\�������Mt�y~(���k��L6��VKJf�M�U<5��<��2�,*+K"�nH�??o���O�������p��S7&7�y��]g  h�1I�%����%����e �U��;�k�x�yOٔ�Qo���=u�;[a�P�V�V��Ҩ�,�Ȧ��$�M)�d|�����vYo��>�4v          p�����uOZ�զ�gi�(�������Eya�$�ͧz`��{w�����4��������u   �6I�-I�$mv�hZ���qdD�i�k�.�w�=����6M�Vgf��ʦ�Ҩ*���V�o�'��          ���3x�&���+S�Y*���P^��	r�r��y-��}~p�$9/�����_\��EIOq  ��%�W�Ւ�&�2�
�.C��?�;���>�.X_x�R�9���iʯX��U��e�*�JJ㊧�O�W4�G�����,�%��$y~P+������I�3��^          @�1~ ?WtcY��xAm���K��Y�4�Q<5�xj�ҙq�Ւ��*���ɴƸ���;W�wiuo�a�ƍ?��{;�r  �=�Z��K��/釒��N�ԾER`�Nh���e=�q
/Z�0ǒ�V~p}#W�8�*�L+�N�FU�qE�2?��g�f��g           ���S�m+M"%���ҤV��2aAA�W~��iK����J�%�qg|����G%}�Y  ��S�t��^��$�R�Y.C.���+��X�6�p~�W=��m�7�YTQ<}P��~E㣪N�*��HY&��x~���#M�         �u����12���4V23���^��Ie�eIT+��'4{p�)�T<=&�&�b����8mcz����,  @��MI��t��jSݻ\�mэ���ҫ/:����H�������9�|n���ҙ)�IE6�%c��N�)�X��>�4v          p����g�u�b�%�d3ya^&�+��WP�uZ5H�S�z���������ǒ����T��   hI/��I�ewt�EMp�k.^����[7��8�YaϊF���JiuZ��AES�ܭ�R��d�����r��0�          Z����]2R�*��T49�dfBYT�1F��kh���͔�'������`z,>�+߹���B   ��D�O%� ����k��͒�s�fQ����s�q����
s���_]�Oo���:�xz��}��G�V�e�T�v^�'��;          �.
�'�x^��`�l�(��P4�WieZ6�d�`�����~�S�e�d��u4�]�cN�|�Gn������   h=���%}^�����;�Ђ��oۖK��x�r�9\q���+�[))O(�>�4�����$yan�V
           Pc�@F�d�����IF~�[A�_A�oyzƨ0|�J�t|az���X����;  ��*��8�$m��UүI�s�8iK��-����a��a����A�L�̤����ܭl��^��>{H0,&�         @�b��r3�	�/e��ʤ�ɽ�*%Y���Y�^��+*)�+K�K���5P���\�����3�B   �����?�G&��&&��-h���W<��g��/w��
C���ql�*�>��<�,.�y���%y|           ��V+��6S<}@��^����b������:
C�4�Џ� ���{�9���6i   K����ϑ�bՎ���0�`����g��]A�v���UX��#�L+ߣ��n�4�1F�e�pof,�         �u1�ݝZ�V�H�3�&F�VJ2���N�q�\A��>�4Y����[��>u�����{܍�  h_���$����%}A�nI���9��qw����>����̯hD��\��	�Ϧ��v���OU=�S6M�s�{-           �f<_^�(ɪ:�G��?Su|�l����hGc��(��Ѐ��!   :C*�NI#��(�4IWH�AҴ�X����}�P�-�Rg���ohQ�I�3*�@�]w+�ʵR�.SB            �� '/�+��4��nU�?�,�,�1r}��)�3��_[��w�  ���/�:I/�4,i�������L���ܯݶ��F��$��+�-�=KZ�Qe����HJS�9��          ��b�'/�˦��{��̞{�E����䅅eNxl�z���[��4  @g+K�.��$�"�tI�?{Y�0:�1����omTI��L&�>}U4����@�f���           xa^���ޯ��eqt��ذ[��Hwt�sW9   ��vH��jS��J�mI����e(t�����K�̡ܺF�90]�_�=��6KU������1�� ��t            ��k���轪�)e�Qok�ݚ(����Z�_��˞y��   8�1I�(饒�U��~��f���Q�����2�qA��j|:��x}R�Ry�=�i$�?�m            �/�+��*�[��ԑo�56]��!6���.   h���$�D���c�H����\h#G,���5�9��5���@���Z/8�
+U�?���n?����=           @�3Ɠ�T=��6����@Q�i�;H������[�Zt   ��I��)����DI��Z�}�]4��#��;�7n~��ҁ�$��#�g��{�M#?8��           p^*��*��'e�!�K��Ɋ�h�����o\��NC   �d����A�
�C���,i����hh%G,�o�~��!&f"%i�8W��"�,Uyt�jۙ�           p�j��L�;j	%i��Q�S����p�V����4    �R�Z�����H�t���J�7I�Β��=����W\���+r��16u��V��P��           �������k��h��C�3��§7��  ���H�OI����HZ/酪��)��CRp�k�rj80}���d�\M�yd/a            ,1#kSE��$�8w�t%Q5N��%�
=�zM�%��I    4ڮ�勳_�Ζ�tIϐ�I�Jj`��=j��)��g42���C���⪒�T##            tc<%���ir��cSUG�j���_�4    \J$�D�u�^.�$���E�� �$頳th�C
�׼����	�Zy%J5��\��L�7{           t�Jf��lb&R�f�I�����x٥��   ��LH�.iD�$��t���$]-�FI{\����џ�^�ȕ�MWuY��ػw�J���)w��ݷ��fw�#�XĠE+$.�M�6\�HHD|���H��Hdh�D 	��l{�>>������m�o��^�<�T��v���Sү��\�<V       �N4��F{��x�hg�}�o���şG�?�   ���߫븧qt��oGį���^D��u;��������}.�&^N�?o�:���       �fk�?z1Y���F1��x|��a� ���������8"����W���{ߎ�*p�������d�a_�_Lў��m"b��5        6�)Gݴ�����w��'"��no��  �6UD�lu���G�o�Q����z��9�������������i��ɲ�Y        \ދ�b���kOƏ���<�����,  �m��븧qt��w��I�ߎ�߈�a��x}���`����~9]Fݞv~;        ,�&&�2vw�{�=.F��n���w� `��E����#���:x?~}z����*p����w�ضGo�       ��/��O�w  r(#�g��mED|-"�ߊ�oD�7W_u��;�lyK�#"��������o��4r0/cY5}�       �U̗u����}���ů�>  .����������""�Ǜ��'q�?����?��S�U�~'�����`��(        ���d������~�;~��P  X�&"�gu��3�����8��?Y}�<���g���w;�wp㈈ݝ���6[V1]�}�       `���x�x'���^�>�S���G�;?����G�� �mD�����s��^��W_�E����z�����ŏ#"팿�ǰ_,�       ����7Yć���>{��֟F��  ^�E��W�E݉���qD<��'�h�������_}�;���^������GD|�;���!U�����z        k�w���D1�:����w{  ��2"~���e7�����j��(���OO"b�������(�?a�ŏ��ç���5.{���e�]       `�ꦍ��2�<�����w�O{  \�d�uo�7.��۵m�w��t        �y1�����z��P  `P�(�󮇼�-����       pS��:f˪יw���:  \qw�u=do�7x       X��ɲ�y�wF[_��v{
  ���5�f���:�˺�        �`���i{�W�Fq����  W��>�r�ޡ��       n�6�oA�n�o�:  Tq�x��͛���i�M       @w�&�h�;�=O��  ���*�tu��e���T        t��������m�'�  Wl�qW7��#�        �^�MH1��  W�ǣ�.n<�����.n       ��&�*e�ˬq�
� `���$p1qz;       �m�w��e�h4���    �b���jb2��}[        ��?\FӶ���Ž·   i�"F�����7t       Fݶ�rZv>g�(�  �A�b���=���#�        NO� �?n  �*�}��yeݬ��        $s��bY�D  ��Y{���v       ����)�  ��Xk�^7mL��:o	       @b{��hۡ�   n�����e4X        6FU�q�p "  �kܿ<��S        �F3  �������yY��v        ��2�z  �X[�w�X׭        �A�p�;  �k	ܛ����r�       �ڟ:  �����2���L       l�y��lY�  pí%p�S        hH  ��v�^�M.�}       ��^N�h�v�5  ��ځ��ԛ�        D�m��� ���v��R�       ��� ��V�(똗ͺv       ����ʨ�v�5  ��Z��7n       8����Y9�  �u����        orh"  pUWܧ�*ʺY�.        ���**]	  pWܽi       �Y����+   7Е����        Nw0sx"  pyW
ܧ�*��]�.        ��eU��  p�\)p9sz;        �v�1  .�J���        ��E  �.�ϖU�>>
       �sLU�M;�  �r�����        \DZ  �r�        t��l9�
  �r��}Qձ���v       ���.�h�v�5  ��R��dVu�        �P�E�   q��}^v�        ���Ls  \̅��m�M       ��M�  �b.�Ϋh��       �[���X���k   7�����GE       p5�  �.�{�        �&3�	  p���n��       �[j���i�'  ��](p?\T]�       �-�F�L�  �C�       @/4(  �y.�O=\        pMw  �<���eu���        ��|YG�C  ����ݛ�        �CZ  ��.��}�       ��  �rn�>[�}�       ��
� �wxgྨꨛ��]        ��eM�G  N���}�pz;        ��F�|�I  N���}�#�        X���  8�9���	        �ˡ�  �Y�ܛ��E)p       `��  �g���M        �˪��Q�   '��ϗޔ       ��e5�
  @Bg��^5}�       �Ѧ   �9;p/��       @7�)  �i�q���        �!p  Nsj��4mTu��.        l�E��  �Щ����        t�nۨj�;  �S�e��       �n-4*  �[�ܝ�       @�J�;  �S���?       �1�
  �S��n��       �S	� ��8�       �AhT  ���q���        ��Q  �v"p��6�v�U        �$e%R  �t"p�f,        }��6�V�  �v"p��        @_�*  �q��C�       �&r#  p܉����        @O�  �qNp       `0m3�  @&'w�;        =q�;  p܉����        @O�*  �q'�!�        `#5b  ���;           A�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           ��&`    IDAT p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
�Ϯ    �Ǝ�Hp          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap     �ع�'�0 �5IFc@�K�y��W\:[G�n�t�qt%���@�?�eUC�P��(     A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�  v�.�    IDAT        � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          ��y�vW����8���q��n�}��z������<�K�      �#l�/ƫ�����i|�����/w���z�����p  `a����ß�<����<���4V+���>���       x��n5^?,�`�3M�q�_�n�۫�^����r�=  ���           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �         �/v�/4��������]��eM7�l梭�FlQ�MYP���:0�FE;�i'�HdA��$7������J=�A�t`�a%�������߿�e����.���^7\'�' � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�    c�.�    IDAT      HA�          @
w           R�          ���          ��           � p           �;           )�          HᲢ   �����D]]]���E}}�������={vDD����e����W�V�?�O������GDę3g�̙3q���8u�T�<y2N�8q�:y�dLLLL�       f�;  @2�j5,X����`���?~466FSS�������5k֤o���8�?~<����������_~�%�=��㓾       ���   ihh��������c������T*=��T*����!b�������~3>>G��#G��������q�������ٳ�       �
�;  �$X�hQ���E{{{���Œ%Kb�ܹEϺ$*�J477Gssstvv�>>>?��S:t(<�}�]�߿?N�:U�Z        �;  �Ev�WƲeˢ����U___���U*�hii�������{#"�ܹsq���ػwo�߿?������k�K      ���  ��������������n�!J�Rѳ��r��������<�HDD����޽{�o��ݻwǱc�
^	       L�;  ��T*�lٲ�����θ�[�R�=k�hnn����X�zuLLLāb׮]�{��8p�@�;w��       �%"p  ���j�q��bŊ��鉹s�=iF(�J���mmm100Ǐ�ݻwǞ={bϞ=q���'       ��  �O���Dggg���Eooo\q�EO���͛������gϞ������O⫯��?����y       �?$p  �/*�J�u�]�v�ڸ��;�Z�=�?Q�V���;�����~�/��">��طo_LLL=       ��   �dɒX�fM�Z�*��ꪢ�p�bݺu�nݺ�O?�4v��cccEO       .��  ���̙��w_�����7�\�.����x�'����]�v�|���q�ܹ��       ��;  0�,\�0~��x衇�����9\"�r9zzz���'�9;w>�(N�8Q�4       �O� ���n�G}4z{{�\.=�It�����`<�����������,z       �?� �i�R�D___<��c���^�
VSSk׮�5k�ė_~[�n�����Y       ��  �R�\��+W�3�<�]w]�sH�\.G___������hlٲ%���ۢg      ��'p  ��R�������OGkkk�s�������+���۶m������I       0c	� �i�T*EOOO<��S�t�Ң�0-_�<^z��W^y%:T�$       �q�  ��w뭷���P���=�i���+FFF��?��_=�;V�$       �1�  ������>�l�Z�*J�R�s�F��r<���q������Hl۶-Μ9S�,       ���E   �P�f͊���ǎ;b����v.��/�<��?��      �$�  Sʊ+bǎ144���E�a��?~lܸ1^{�X�hQ�s       `��  S¼y��^�͛7����u��ǻ�6l�rّ       .6_� �������ދ�+W=b���188���q�M7=       ��;  ���W_/��b<���1w�ܢ�����[�n�����V�E�      �iA�  �S*�����?z{{���R�Ćbxx8n��Ƣ�       ��'p  R�3gNlڴ)�{3gN�s�/iii���~;֯_�R��9       0e	� �4���cxx8�瞢���V�144�7o������       ��$p  
W*�b�����o�5�\S��Gz{{cdd$�/_^�       �r�  @���_�����5kV�s�hjj�-[����@�ˎ�       �W��  ���=�o�w�}w�SࢫT*100�7o���ڢ�       �� p  
���[�l���Ƣ��%���o��V477=       ��  ��T*ņbӦMQSSS��K�.�w�y':::��       �	� �IS�Vc�ƍ188��3KCCC��꫱z�ꢧ       @Z�  `R466�o��V�*z
���;��0�}�C�B�*A��0`�D�ƙD�n6'j93�K6���L��L���d���$_�I�RS��dh64eQQpąTmi�>�y߼�D���9�uU�K��*i�s����imm��~��q�5�D�R��      ��c�  ��1c��7���x��^���*�J\y��O��O��ښ�       u��  �U'�xb�~��1jԨ��+��Ϗ[o�5��ڲS       �n�  ��u�{]�~��1|����Kg�uV|�k_�A�e�       @]0p  z�Yg�_���cȐ!�)P�N;���׾C��N      �t�  �7gΜ���[���-;	��        ��  8�f̘_�����5;�	'���ַb�ر�)       ���  8b�M�_����U9rd�v�m1jԨ�       Ha�  �'O��o�ٸ������n�#Fd�       @�� ����׾6n��hkk�N��0bĈ��W��sLv
       ��  8,�Ǐ��}�k1p���h*�ƍ��|�+�l      P*�  ��6|���[b����)ДN9�oG       �T� �W���-n��8��c�S��M�<9���/Ekkkv
       �:w  ��V��/|!N9��(��ӧ��>���T*�)       Ы� �W�n�Y�feg@�\p�q��Wgg       @�2p  ^�����q饗fg@)]y�q�Eeg       @�1p  ٬Y���`v�V�R�O}�S1u���       ��  �!1bD|�s��jկ����5n���;vlv
       q-�  @�kmm������g��tuuŎ;�^��������>���===�w��8p�@DD���EKKK���D���#"bРA1lذ:th6,�����6x����W]uU����9       p��  �G>�8��S�3�����غuk<��c����O<�<�Ll߾=�~��^;����СCcԨQ1nܸ8�����Q�FEK�_-3�x���/~1>��Gwwwv       V  ����׿>����gg������G�|0|��ظqc<��q����;�o�۷o����������8qbL�4)&M�S�L�#F�Wf�sN����}|���N      �#��  xY'�xb|���(�_|1֭[k֬�_��W�q��������cÆ�aÆ��wÇ�3�8#�;�8��sc���������/���?����       8l�  �Kjmm�/~���֖��Զm�w�uW,_�<֭[����N:l�<�L,\�0.\�j5&O��f͊��??N:�켦S�V���|\v�e���Og�       �a1p  ^�5�\c��K��X�pa�u�]��#�d������X�vm�]�6�����ĉ�o|c�����!C�d�5�!C��M7��\sMtwwg�       ��f�  ���S��{��쌦���q�wƆ�s�lܸ16n������f͊�/�8f͚�j5;��M�:5������W���       ���;  �G���ⳟ�����q�������/����g�ԍĲe�bٲe1nܸx���o|����5;��]v�e���&V�\��       ���
  �G>����ѣ�3ZOOO�u�]q��W��������n��g<����/~1.�䒸�;����NjX�J%>����q���       ���;  �{�sN��-o��hX�Z-V�X�]vY|�����/;���ܹ3��o��__��W���+;�!<8>���F�R�N      �W��  �����>:n��F��W����.�,n��ؼysvNCۻwo|�{ߋK/�4~���EOOOvR�9���mo{[v       �b�  @DD\}��1|��쌆�y����c���iӦ윦���O��?��x��������s�>��5jTv       �"�  @�?>���wfg4�^x!��կ��_��w_vNS{�G�k��O~�{��윆�������Z��?       �÷�  Pr�J%>�OD�>}�S��ŋ��xG|�{ߋd���ŋ���~wtttd�4��O?=��wdg       �!3p �����cʔ)����3n�����'?;w���)��;wƧ?�����g���i�]w]�3&;       ��;  ����������h�V�����=�_�";��X�bE��}�+Vd�Խ���Ǎ7�ժ�        ��� ����kcȐ!�u���'n����?O?�tv`׮]�`�������_�ΩkS�N����m�       �� @I�|����7�9;���޽;>���w���j�9��Z�?�я�+���{,;��]s�51t���       ��� �������V�J�rz������X�jUv
���G�+��2�-[��R��]w]v       �Y�,  PBg�qF̚5+;�n�Z�*���ؾ}{v
�@WWW|����~����ӓ�S����7ŤI��3       �e� @�T*�����3��O~����?]]]�)�
�Z-����ł���3;��T�����>��       �-�h @ɴ����ɓ�3��m��7�tStwwg�p�V�\W_}u<��3�)ug�ĉ��7�9;       ^��;  �HKKK\{��u���F|�;����ڼys����m<����)u�뮋!C�dg       ��0p ���Kb�ر�u�V�ſ�ۿ�wܑ�B/ضm[����]<���)ueРA����       �'� �$ZZZ���/�Ψ+�Z-��_�5����g�Ћv���^{m�Z�*;����-o��O>9;       ���;  �����9rdvF]����?�avػwo,X� V�\��R7��j\s�5�       �G� ���j\v�e�u��?�q�q��h����O|"~��_e�ԍ��??�L���       �g�  %0o޼8餓�3��]w�_�җ�3H��/Ƃb͚5�)u����N       ��3p �&W�T�+��Ψ6l�O����ӓ�B�}��łb����)ua�ԩ1s���       �w  hz3gΌ	&dgԅ;v��?��ؿv
����7�pC<����)u��믏j�G       ���5  4��/�<;�.�߿?>�я�3�<��B�x�����p�ܹ3;%�����.��        w  hf&L��S�fgԅ���6dgPg�n���G���+;%��W_---�       ���;  4�K/�4;�.��g?�;�3;�:��C�g>�����NI5v�ظ�⋳3       (9w  hRC��׿����n�_��3�sw�}w|�����H����?��铝      @�� @�z������������o�={�d�� ���o�ҥK�3R�=:�ϟ��      @�� @�V�񶷽-;#�7���X�~}v�V��M7�O>�dvJ��/�<*�Jv       %e�  Mh���1r���T�<�H|����Π�tvv��>��طo_vJ�SN9%fΜ��      @I� @���K�R�����������N�=��q뭷fg����˳       ()w  h2#G����>;;#�~��x衇�3h`?�������H3u�Ԙ:ujv       %d�  M�MozST*��4۶m��o�=;�W��⦛n�]�ve��q�      ��  �D*�J\x���n���ػwovM`׮]��}.j�ZvJ��3gƄ	�3       (w  h"��~z�3&;#�ڵkc�ҥ�4�{�7~�dg��T*��w�;;      ��1p �&�7�);!M�V��|�+���M��[�w��]vF�������C�fg       P"�  �$�:�hoo��H�p��X�n]vMhϞ=q�M7������R?8      @�� �I̝;7����������=;�&�z����O�����o{T�>>       ��� �&q�Ee'����~۶m�Π��z���3�dgnԨQ1s���       J��  ��������Hq�����;�3(���θ��[�3R����N       �$� �	�w�yѷo��?���ⷿ�mv%�p��X�fMvF�f̘�ƍ��       �� �	̙3';!Ewww���Gv%s��7����3
U�T�mo{[v       %`�  ���5�=����-��[�fgP2�=�X|�����(��_�����       ��� @��>}z���eg�������J����v�ر#;�P�.� ;      �&g�  n�ܹ�	)֭[6l�Π�����[��VvF����7f'       ��� ��U�՘={vvF����	����Ŗ-[�3
u�gƨQ��3       hb�  ��&O�C���(��O?K�.�Π亻����o��(T�R�7���       41w  h`ӧO�NH��$����3 /^�ׯ��(���ƨT*�       4)w  h`ӦM�N(\OOO�y���{e��>v�ؘ4iRv       M��  T�����N��(ܯ����o����z��X�vmvF�.���       ���;  4�3�<3��훝Q����'�	�'����f'�������5;      �&d�  jڴi�	����e˖eg��X�re<�����8p`̞=;;      �&d�  j����	�[�lY�����'j�Z�q�������       hB�  Ѐ�'�|rvF�,Y�� /kٲe��Odgf�̙1p���       ���;  4���:+*�JvF�:;;c�����zzz�?�avFaZZZb����       4w  h@�'O�N(ܲe������g�y���/dg���=;      �&c�  hҤI�	�[�xqv�E]]]�ӟ�4;�03f̈��>:;      �&b�  �o߾1a�B�ݻ7֬Y����G?�Q���dg���5fΜ��      @1p �s�)�DkkkvF�~��_�����3��<��Sq��fg���=;      �&b�  f����	���/�� �ȝwޙ�P�Y�fE�~��3       h�  �`&M���P�2]æ9,_�<v�ڕ�Q�~���9眓�      @�0p �S����m���'��΀W����_�";�0����	       4	w  h C��Q�Fegꗿ�ev�*?��O�
3{���۷ov       M��  ����R�dgj�ڵ�	�l޼96nܘ�Q�ęg���      @0p �r��'g'���F��ё�P�3fd'       �� ���m�s��غukv�j.�Z���Q�s�=7;      �&`�  �l���?;��������(�I'�#F���       ��� @��T*q�'fgjݺu�	p�/^��P�s�9';      �g�  �㎋dg�,��in�/�Z���Q�s�=7;      �g�  ��O�N(T�V�M�6eg�a۶m[<������6mZ���';      �f�  �l��[�ƞ={�3��X�revB!�&M��       ���d   �����N(���4��+W�UW]��Q�s�=7֮]���hkk�׿���ix��x�G�3�!T*���K�Z-�]��{,����     (=w  h�G�Θ2�.    IDATN(�1"����]�v�СC�Sz݌3��n����ݻ7���9rdvJ�+V�7ܐ�a�����O:;#͍7ޘ�      DD9O�  @5jTvB�\p�����Ľ�ޛ�Q��'Ɛ!C�3��Z-:::�3�L�>=�����=;!���������      ��  B߾}��c���(�����d'�u�=�d'�Z��駟����Q�{kkk̚5+;9s�ҬX�"��ٓ�     ��;  4�#FD�Z���8p �mۖ�G��ի���';������-[�dg�)�Uj8T��zj�=:;#M�    �zS��  4����~���FwwwvQ�w�M�6egb�ԩ�	��ŋg'��9sf���?;�Z�ٻwoi޴     ���  ��Q��
��Of'@�X�zuvB!&N��������������4GuT̜93;��ܹs��,_�<��ݛ�     ��� ����O<�� ��,����8��S�3�?�l��>�hvF�2_���d���q���gg�Y�hQv     �� ����SO=�� ����_|1;�S�N�N�%tttd'��5kVu�Q�P��� Ȟ={��{���      ���;  4�c�=6;�PO>�dv��������3
1eʔ�^��Ҵ��Ō3�3�.�y�t��ؿv     �� �6,;�P۷o�N�^s���g'���O�j���橧���7fg��7o^vԝq���I'������o�     �z�f  h �sLvB��~����5k׮�N(ĀJ=��gesΞ=;��훝ue����	i���X�fMv     �� @�kkk�~��eg�^������5�ׯ�����B�~���	���F�V��H1p���6mZvԕ����4�/�dg      ���;  ԹaÆe'�g��N�^����6m��(Ĕ)S�x	۷o�6dg�)���Q�Fń	�3Ҕ��     P�� ��s�1�	�z�駳�׭]�6;�eMֻ2�:�̙}���΀�0���4;v����7�     �K0p �:W�����۳��=����	�8���㨣����%,Z�(zzz�3R<8�<����e~���ŋK�s     ꝁ;  ԹaÆe'j�Ν�	��6nܘ�P�>}�����3x	�>�l����i�<��ϱ��{��3�,Z�(;     x�  P��v�����N�^�e˖ػwovF!^���f'�2:::��̛7/�U�Qn��ϏJ�����駟�u��eg      /�7y  P���P(wʠ��'6mڔ�Q���dɒ�����Hq�1�Ĕ)S�3 ռy��tttDOOOv     �2� ��}���	�2p�,6nܘ�P�	&d'�2v��k֬��H��ޞ� i���G��`     ���  �\[[[vB�����(�#�<��P��O>9�U?ԫ2�<�ϟ�J%;R�����g�֭[㡇��      ��r~�  �l�w�ޝ� �x�ǲ
ѿ�7n\v/c�ҥq����Ç��N;-;R��Q�ղ3     �?��  �\��.�S[�l�N(�k_���^Fggg�^�:;#ͼy��pC��3�8#;#M��\     ���  �\��]]]�	P����x��g�3
1a���2�=/����T*�P�9s�D�>}�3R<���iӦ�     �/0p �:W��{OOO�߿?;
��c�e'����lٲx���3R�9��N{{{vB��f'      ���  �\�����Z����)����N�N�����{�';#ͼy��0���>;;#͢E��     �C`�  u�R�D�~��3
�o߾�(ԓO>��P�c�=6������ё��f����	P�ٳgG߾}�3Rl޼�4�    @�3p �:֯_��V�����{�f'@��mۖ�P�J�cǎ����X�bEtuueg�7n\�|���P�����4e~�     My�2  ЀZZZ�
e�Nٔe��#b�׾}�bŊ�i�<��<���bƌ�i-Z��      "w  �ce���K(w�I��ϛ7/;z�y�����)|��x��'�3     �CT��  4��]p?x�`v�^�����B�׿{�7^x���Ǐ�N8!;zU��(�<     Ј� �����';�P===�	P��\q7p�����˗gg��;wnv��~���̙3�3R�j�X�dIv     �
� @+�����;;
���f'����N����q{{{v��s�=7���bݺu�y�     ���;  Ա����B�SF;w��N(���cȐ!���V���{.;#�ĉc�����+�� G��    �Fe�  u�wh~e�GD�7.;�������t���4s���N�#���5�;��===���     ���  �����4p?���8e�v\�+�4�s�9'�>�����w_<��3�     �+d�  u�Z-�_�{zz��p;v��N(�رc�8������g���H1iҤ8��3��*�e~`     Y��2  �`j�ZvB�*�Jvn����	�9rdv����'�.]����R��ܹs�3��iii�ٳggg����.��2     ht�  PǺ���
էO��(ܞ={�
s��f'p��|���׮i>g�}v4(;#��իc׮]�     ��`�  u�����	��V��B�tuue'���N��]�6~���eg�8����5�yMve~`���     @�� �:�;4�2]p>|�YD�V�%K�dg��V�q���gg�a�V�1gΜ���˗gg      ��o� ����{KKKv�L��}��СC�38D�-�NHS��4�3�8��?s���x���3     �W��  ��������V�eg��c��N�mذ!�z��g�uV2$;K������N      ��;  Ա����뗝 ����dg���N�X�xqvB�>}���矟��Z�Z��s�fg�ؿ�X�";     8�  P�<��P(wʪL����X�|y޼y�	�M�<9�������={�dg      ���  �X��mmm�	��L�]po,�<�Hlٲ%;#�9��΀W��h,Z�(;     8L�  P����===��q���*�����SֱhKKK�w�y���U*��������sOv     p�� ���j�ػwovFa�� )�4pw���,\�0;!M{{{v�b��zj�92;#����K�wg     hV�  P���ٓ�P��}�Fkkkv���;;�0�g˖-�y����{n���eg�+R�3:::�     �#��  �\WWWvB��� �kii�N(̰aòx�:mmm��3gfg�+2w��������_�2;     8� �ν���	�2p���:��´��F����3x�:::�V�eg�(�5l�)���ƍ��H�lٲؿv     p� @�s��_߾}�
��y�yꩧ����Hq�y�E�~��3��������i     ���;  Թ={�d'jȐ!�	P�J��������1�u<گ_�8�s�3��̟??;!��ݻc͚5�     �b�  u�lw��)�D�Z�_��9oL.�Z������W�i�|�p�	�)�,Y��      ��r}�  ���3;�PÆ�N�B:4;�p�i���~���s��)ݛh<\pAvB���a     ���;  Թ�;wf'���N�Bs�1�	�2dHv�RYG�mmm1mڴ�������;v�}�ݗ�     A�  P�v�ؑ�P(wʦ�w�עE����';#EY��4�ѣG�)�����b��ť��     ���  �\�.�{��	P�Q�Fe'���U�K��~���';^����Ҕ��     ��� �Εm��;e3v���¹����:&<xp�}���������۷Ǻu�3     �#��  �܎;�
����΀q��{c[�dItwwgg��7o^v���;.N=���Q�ղ3     �#��  �ܮ]�J7�)����7n\vB�\pol�w�5k�dg��;wnT�>N��̟??*�JvF���Q     ��o�  ��<x0�{��B�S���Çgg���W�Q�1�S�N�΀?R�7lݺ56nܘ�     �w  h ;v��N(T/ZSN��zj)��e'p��.]�����H��ޞ� �7lذ�<yrvF����-G     P�  � �mۖ�P�1c�d'@!&N��������	����X�jUvF�y��E��#5�C{{{i�y,�$     ����  4��[�f'�wʢ�����hmm���0�u\:|��8�Ӳ3 "��F�-[���͛�3     �^b�  ෿�mvB�N:��^#�\�L����樣��N�0-_�<^|���eS_�S�N��HQ�l     �,,F  ���{���c̘1�ЫN<��>|xvF�����SWWW�\�2;#E{{{T*��Jn�ܹѧO���-�N      z��;  4���#"N9���UӦM�NHտ�����^Q9rdL�0!;��+�6m��=�Xv     Ћ� �lݺ5j�ZvF��ivg�uVvB*��r�������HQ�q1�a������HY�    �21p ��o߾عsgvF��if���1}���T��a߾}q��wgg��?~v%6gΜ�۷ovF�ŋg'      ���  �SO=��P��N;-;z�Yg�G}tvF*��hѢ�cǎ����ggPRe}��<O>�dv     ��� �Alٲ%;�P�sL�=:;z�ܹs���7�{�':;;�3R̛7/;�jkk+�[@:::�     �� @�ؼysvB�&O��� G\�Z�ٳggg�3po��˗gg��?~v%4{��hmm��(\�V��K�fg      0p �QƁ��I����;��3�5�yMvF:��R֫�'�tR�p�	��L{{{vB��k�ƶm۲3     �� @�x��G�
7eʔ�8����7e'���jժصkWvF�y��e'P"����3fdg�X�hQv     Pw  h�w�;vdg굯}m4(;������ܹs�3�BkkkvGPwww,[�,;#EY�i�c֬Y�|@���'�.]��     ��  ��͛�
U�V㬳��΀#�.����쌺P��H��tttd'��0aB�3&;��(�~���3�<��     ķ�  �@}����M�6-;�������	u�����y�Z��1�jmm�Y�feg�(�4     PV�M ��iӦ��M�>=;��SO=5&M���Q7ZZZ�8�zzzb�ҥ�)�)3�裏��(\www,[�,;     (��;  4�x ;�p�ƍ��#Gfg�a{׻ޕ�PW��铝@/X�hQvB��N;-F���A�koo�NH�jժصkWv     P w  h �?�x<������?~v��C��\��QWܛ�ڵkc۶m���T*1w����XKKK�w�y�):::�     ��� @��j���n�N�{�;�����u���9�j�X�tivF��^צӦM�A�eg����|���     �`�  �`֯_��P��N;-F����J�����xGvFݩV}$Ѭ�zmyʔ)1|����TY���{���3;     (�o� ���q�1o޼�xU��ַƐ!C�3�NKKKv���'�|2;�p�j5�?����P���*�3     Pv�  �`6l�===���袋��kii�w����u�O�>�	��ŋg'�(�mzיg�C���(ܾ}�bŊ�     @w  h0{��-[�dgn���1q���xE.��1bDvF]2pone��|�Yg�r�L�*�+W������      ��;  4���?;!�%�\�� �쨣�����*;�n�7�M�6�c�=��Q�j��g��Π�T�՘;wnvF��>(     � @CZ�zuvB�7��q�QGeg�!y׻�Ç�Ψ[ժ�$�ݢE��R���6�cʔ)�׼&;�p]]]�r���      �o� ���W�������0 �ϟ��������vF]s����������c����4�y��e'��뮻��_��      �� @��쌇z(;#Ż���������4hPvF]+�C:e�e˖ؼysvF�ZZZb����4�J�Rځ{Y�     ���;  4�իWg'��8qbL�:5;^։'��^zivF�����N� e����g'�N;�1bDvF�:;;K��\     �� @�Z�jUvB������	�>�DKKKvF�s��.\�Z-;�p3f̈��>:;�W���K�.����gg      �� �A�_�>����3R���1f̘��\pA̘1#;�!��^[�n��7fg���5f͚��A�+����o~      ��  Р8���o�3RT�ո�+�3��4(,X���0\p/���U�:N�Ș0aB)�۽{w�Y�&;     Hf�  lٲe�	i.��=ztv�ނbذa�������Z���Q�Y�fE����3hP����	)�,Y��     ��;  4���#�������+�3 "�w�z�fg4����*��۷Ǻu�3
ׯ_��1cFv��o (�     �?f�  �瞋��?;#�E]cƌ�Π���ԧ�3NOOOv*�h��W�9<'�tR�p�	��۱cG�w�}�     @0p ��dɒ�4---q�u�egPb�J%>�����óS���x��R>�0{��hmm�Π�����E����     �� ��-Y���c�����ԩS�3(�K/�4�̙��ѐ�˥������b����4������     �O� @�۱cG<����,Xժ_o(������@vF�2p/���W�:V��;vl�?>;�p۷o����gg      u�  ���%K�RM�0!.����JdРA�/})Z[[�SV��<QVK�,��fgnΜ9ѷo��DY�X�pa�j��     �N� @���^������?C��Π��j��?�c�3&;����^>�w�5k�dgn���q�gfg� �:p/�     ��f�  M`�Ν�r���T��}�C����>���9sfvF�3p/���X�:Z�9rdL�81;�pO=�T<����   ���޽GY]���f������xC�
3d�.��g%m�ilOln���$ͥ���+�9']��JN�6M�jM�����&���T@@E�@DPQn��������$g�����z��Z��̛�&�?�g Tw  �?�я��]u�Uq��ggP������5�\��Q:;;�H�hѢhoo��(\SSS���+;�
���uuu��kii�����     ��� @�X�|yl߾=;#ݍ7�����ΠM�:5�����5�������>�`vF�_|qv�������     �k3p ����?��O�3ҍ=:>��OegPc�=�����{��N��	$)똵��);�
6|��8qbvF�6o�7n��      *��;  Ԑ���U䈸ꪫ�o}kv5�SN��~����ؘ�RS�=��@�x <��Q��s�F}�?���555���Ǽy�     �
T�WM  ��=���bŊ쌊��|&F���A�9rd|�ߌ�C�f�ԜC�e'������lٲ��6,.����*TsssvB�����     �� @���~��PN<��������ׯ_v
Uj�С���=F���R��˭��֦���*����㢋.��(�SO=�7o��      *��;  Ԙ�˗��O?��Q�>����g?��A2dH����}�;6;�fn��    IDAT����ŋc������;wn���egPa����W�^��kii�N      *��;  Ԙ���������Q1��ַ�{�������'����g�qFvJM3p/����X�dIvF�F�&L�Π������     �
e�  5��{��쌊�},�O���A7n\��?����0p��כ����� �K.�$;�p�?�x<���     @�2p ����w�qGvF��իW|��_�/�0;�
v���Ƿ���>|xvJ)��|��سgOvF��Ν��@�3gN���';�p����	     @3p �u�wD{{{vF��ׯ_|�+_�1c�d�P������ַ���N)w�9��vF�N9�8�쳳3�e�����,��      *��;  Ԩ�������QQ�_���c�ȑ�)T���������_�b444d甊�;---�	)�8j�7566�e�]��Q��k��/���     T0w  �a7�|s>|8;���=:���o��ѣ�SH���_��������e甎�;+V������½�-o�N�\q��|����      o��;  ԰�;w���*F��w�F��N!�g�����s���N)-w""�=.��(�駟cǎ�� Y/�wvv����3     �
g�  5�_��_\q�G��o}�[q�i�e�P����mq�-�ęg���Rj��RY�9�q����_�~1u���­Z�*v�ޝ�     T8w  �q;v�;�3;�"�5*���).���
p�	'�_��_��?��8��sJ���=:;;�3��W��;vdg����f̘�����(\Yh     ���;  ������Z�k4hP|�ߌ+��2;�t���ǭ��������B��ί��쌅fg�sΉ1c�dg���8ttt��u     ��� @	�ڵ+n���쌊���_��������e�Ѝ�n�����O?=;��p����*LY�:755e'����!f̘��Q��z(^~���     �
� @I��?�s���egT���������+_�J0 ;�n0a��[��菢��o+����G}4�mۖ�Q�2^�&bڴi��ؘ�Q��>�     ;�� @I�߿?���oegT�+��"n��8�쳳S8N����O~�q��7�Yg���ë0p��uuuł�3
7a5jTv+������x���3     �*a�  %���8֯_��Q�ƌ7�|���Uh֬Yq�m�Ż��n�*�����@e��\WWWʱs����;f͚��Q��˗Ǿ}��3     �*��~  (���������fgT�����������c����9����>;���o���?�'F�����0p��<���u��������_��(\`     ���;  ��ʕ+�����Ψ�&M����.�W��N:)>����w��ݸ�˲sx���ٓ�@�jmm�N(�\Ç�Π e|��СC�dɒ�     ��Xg  @	}�k_�ÇggT������'?��/�\pAvѿ���?w�qG�����A�ٻwov��W����cΜ9����>f͚��Q�%K�ā�3     �*b   %����w��쌪3~����w�����⤓N��)����x���?����`466f'q�y-7n���~:;�p����	`���1dȐ���     ��1p ������ذaCvFթ���w��q�w�G?��0`@vR)466Ƶ�^?�я��믏�f'�&�ٳ';�
��ښ�P�I�&�r�\6e|�����lٲ�     ����   r=z4�����q��7G�^��s�N�~�������|g|�{ߋ������쬚3t��x�{�����_�~����/��G��|�;�r���o3o޼��?��Q�����={v��G?�N������W\��Q�E���Ç�3     �*c�  %�~����~�{���S�ր��믏k��6����=n��رcGvV�;�����}o����n444d�t�իW�����DWW�+_7m�4w�5�<�L���?���>;;�P����5좋.��N:);�p---�	     @2p ������MMMq�)�d�T�O<1���ڸ����{����u��egU�N8!�Ν�x�;⢋.�����ns�����W��+�������'�2p������n�>y��8p`�ٳ';���ܜ�P��{���?��     T���    סC��_�Btvvf�Ԅ>}��;�����?�A\s�51x��쬊U__�&M��~��q����?�����kj�q�w�ƍ��j���zZZZ~ぐZ׻w�5kVv=���.fϞ��Q��Ƒ#G�3     �*�;  �W��[n�%���씚2nܸ���?7�pC<����p��x��J?��իW\z����s�̉�C�f'��ݻwǷ���W���^p߷o_v�瞋'�|2�;��B577�O�����ĉ��O��(\KKKv     P�� �����w�S�L���??;�����'f͚�f͊�G�ƪU�bѢE��C�֭[��
1bĈ�2eJ\~��1u��4hPvRa��o�޽{_��\p�����R����_�������g�Ѝ����
���+W���      ���;  G����˿��}�{��*]�^�zŔ)Sbʔ)��/Ɗ+b�ʕ��#��/��\�=F�'N��/�8�L�cǎ�NJ�f͚�z������.�yCZZZ�c�X���g����!f̘����N�͙3';�p,��G�fg      U��  x�s�=��_���SJc�ȑ񶷽-����ED��ݻ�'�x�����رcGr�k�����O>9�8�?~|L�81&N�Æ�NKw�С���]]]��}��0�������3;�*�}��x��G��/�N)Tss��{9��s��SO��(\KKKv     P�� �_��,�N�W]uUvJ):4fΜ3g�|�����[�l�͛7��͛c۶m��/�Ν;c������ޣM}����O>9F�#F���O>9Ǝ��~z�;6���ף��Z}�ߌ�[����S��{���N������n�>}��8������)t�������ܹ3֬Y��     T1w  �7�����cܸq1~�����]��0aBL�0�U����-v��{��}���޽{c�޽q�Сؿ=z4"">���_�~ѧO�W����!c��1`��8p`�x�1x��<xp1?���#������߯���9��ϏO|�Q__��R�~������c����)t�2�[ZZ�S     ��  �������O:n��2dHv�cȐ!�>U�����74�s�~�]�v�#�<�'O�N)TSS��{7n\�;6;�p---�	     @�+��+  ��l۶->��đ#G�S��|��_��{�}�A��pM�y�嗳�2e�Μ93�3x�����
��/ƺu�3     �*g�  ��5k��׿����K�.�;�����`Meڷo_vUf����{ت��1�N�����TƁ��y󢫫+;     �r�  �ou�m��=�ܓ�o۶mq�M7Ӱo��=XT���ڲ�2{�쉕+Wfg����Z2f̘7n\vF����     @�3p  ^ח���x衇�3�butt�_��_��/���LCCC�p�	=XU�v�ڕ�@*�hv֬YѧO����[����=�쳱~���     ��  ����#>��Ć�S�"}��_�G}��~̠A�z����޽;;�*�p��hoo��(Ԁb����������͛7/;     ��  �r�����?��غukv
T�������c�q쁚��;�c����|����577g'pF��Ǐ��(\�i     ��  �������㥗^�N���e˖�җ�t\?v���\S\p�x�q<;{���իWv�h�ܹQWW��Q�͛7ǦM��3     �a�  �-[��'>�8x�`v
�ڳgO|������׏4hP7Uw���ŋK��=��I�&egp��xy�����N      j��;  p�����?��8p�@v
����o�1�l�r����#G�Ğ={�3�R�e˖eg��c�j6|��8qbvF��ϟ��      �w  ฬ]�6>���SJ����X�bś�즚����]]]�T������555E}�?«���QWW��Q�6��͛�3     ���1  อ^�:�����ȝR����'?�ɛ�8C�톚�k׮��ܒ%Kb�����6lX\x���Ae��_�O     ��e�  �)k׮5r�4,X����-���]{{{,^�8;�pMMM�	�C���.�(;�P]]]�     @�3p  ޴_����ݛ�=fŊ�W�W����-���ݻwg'P�8��;wn���eg�:�̙������u��Ŷm۲3     �S�W\  ��v����>/��Bv
t��k�Ƨ>��8|�p�}�aÆu�Ǫ.���/_{����(Ԉ#������u477g'���      =��  �6O?�t\w�u��SOe�@�y������������q�x���������-��(\���dРAq饗fg���3Z[[�3     �d�  t��;wƇ>��x衇�S�M[�~}����߻}�^__��֏Yv�ޝ�@�(���s�f'�[̞=;z�ꕝQ��k�Ǝ;�3     �d�  t�ğ����r�H�X�~}|����{�v��8p`醐mmm�	Ԉ�+W�����ѣc�������������y     @O1p  zD{{{|�s�����������8&k֬�n��G��C�푏[�v�ڕ�@�8z�h,\�0;�p����	��O<1�L���Q����X�`Av     P�� ������rK|��-ݥ]�עE��c�X�ٳ��>��;�ye�=w���^�W\}����(�ʕ+c����     @�2p  zܪU����<��S�)�[�v�m��q����<Æ�я_����c߾}�ԐիWǎ;�3
u�i�řg�����ijj�N(\0     �c�  ��矏|���,;~Cggg|��_���ۿ�����|#F����Qiv��]]]�Ԑ���X�`AvF᚛���Oc�ԩ�����E�eg      5��  (̡C����||�_�d�@D�����������~a�s�ȑ�}�J�}���jP�H�W�3fD߾}�3
��C��/���     �0w  �pw�}w\s�5�f͚�J�^��|�#���Z��-����_�N�=��c�m۶�B�u�Yq��gg����A,     �e�  �ضm[|�#�o|���ё�C	-^�8���0���?��#
���\p�'tuu��J%�3gNvѷoߘ6mZvF�������      j��;  ����3n����Ї>[�l�Ρ$:::�k_�Z|򓟌�{��4><��fڹsgv5��פ�x5�M�6-�3
�lٲطo_v     P�� �t�?�x\}���o|#��۳s�a۷o�믿>��_�5���Rz��C�M�ܙ^|���j����c�֭���0aB�r�)��W���@	     P<w  �"tttĭ���{��b����9Ԡĵ�^k׮M�8餓���|�߱cGv5���5;�p�g��N(�>}�Č3�3
u�СX�tiv     P�{E  �h�7o��|�#q�M7E[[[v5���-n���������55r���.�ӓ�xU����+ɔ)Sb����Z�xq8p ;     (w  ��tuu�=��W_}u�ۿ�[=z4;�*u�=�Ļ����{�S^1|����=z4v�ڕ�A۸qc�����(�\P�f*A0(�$     @w  �b����_��_�{��?~tuue'Q%v����ԧ⦛n��_~9;�W�=:;�p۷o��
=���5;�Puuu1{���R�իW̚5+;�P��˗gg      %a�  T�-[�č7����cݺu�9T�#G��m�����vΫ*������N��x]��W�+��ɓc�����Z�hQ>|8;     (	w  �j�Y�&�����g?O?�tv���+�ϟW_}u����m�߿?;�5�r�)�	�{��(�g�y&�z��B]|��1lذ��ijj�N(\      ��  U���+ZZZ�k��?��?�'�x";�d�֭���q�7�֭[�s^���s�6­���ٳggg�J�;߻wo<����     @��  U���3/^������Ї>+W��N�`۶m��n�)���X�fMv�R__#G���(��;Eiii�����B��x�2^�_�`A9r$;     (���   o֚5k�����^zi��}�iӦE}��ykզM����n̛7/:::�s����ã��!;�p۶m�N�$���x�'b�ĉ�)��<yr<8^z��Rhnn�N(\��     �g�  ԌU�VŪU�b����_���?��?���gg�M֮]��zk,Y��j/4�r�)�	)�{��J����T�^�zŬY�����N�yuuu1{���B���ŪU��3     ��q�  �9;v��|�;����=���/���볓8N����`�������`,^��j���F��N(\{{{�ڵ+;�iii�����B��x���??F���Q�����ѣG�3     ��q�  �Y����+��8���o}k��-o��Çg��:v����{o�y睱u���nS���>�lU?�@�ٱcG<��q��g�fʔ)1`��ػwovJM+�---�	     @	�  ���O�O<_���bҤI�ַ�5���c����i�����X�ti�}�ݱlٲ����N�ve�oٲ%;�jii)���O�>1cƌ���~��R��̙��P��;w�ڵk�3     �2p  J���3V�Z�V���|�+q��ǜ9sbƌ1lذ�Rڸqc��'?�{�7��ڲsz�駟��P�g�y&;�jmm�O|�ѫW���477���	&��!�y��Egggv     PB�  @i9r$�,YK�,����?~|̜93f̘&L�����Ě���6l�ŋ����O=�TvRaN;��������-y䑸�˲S
3mڴhll�d�Ԥ����µ��f'      %e�  �ot�~��X�~}��?�c2$�O��'O�I�&��ѣ��Z{{{<��#q���ǒ%K��_�N*ܰa���O��(ܖ-[�(����R����ӦM����g�Ԥ9s�d'�^�u��eg      %e�  �*����?�i���?���#FĤI�^�2v�ب��K��l۶m�U�V�ҥKc��奿*\���.��g����O}*��铝R���f�p�Yg�駟��Q�y��EWWWv     PR�   o���������/""&L���ǿ���SO-�轳�3�~��X�n]�^�:y�ضm[vVE)�����^��_~9;��ڻwo�X�"�O���R�3fD߾}�����)5���9;�p---�	     @��  ��_~9|��x��_�������g��{n�;6N;�3fL�1�������y��شiSlܸ1֭[�ׯ/����S��[�l�N��ZZZJ5poll��S����ߟ�RS�6p��gcÆ�     @��  t����ǚ5kb͚5���}���1cƼ��SN��Ç����㤓N��C�V� �СC�k׮x����g���{.�n��7o��[��ѣG��N/�o޼9;��[�hQ�x���А�R���&�nt�i�řg���Q�_�[     @w  �v���ظqclܸ�U��w��1t��1bD6,'�x�|�߿�+]__��������""��룳�3���b�޽q������#G����_��ݻw�K/�j�Γ    IDAT�w�]�vE[[[���Ů]�\c�e�����N�����˗/�ٳgg��+��>}�đ#G�Sj�ܹs�
��Ғ�      ���;  @����ؾ}{l߾=;�һw�8��S�3
�iӦ�����R�O<�Ę2eJ,]�4;�&477g'jӦMN     ��g   @�;�Ӣw��=c�Z�Z Ez��������jjj�N�	�G�����gg��v     ��  @7n\vB�^z�صkWvġC�Jw�|���ѫW�쌪7w�����     ���   zX�6m�N�W�m�;hР���K�3�^�.�_�>�nݚ�     `�   =��r-]�4��ۗ�Q����섪6bĈ�8qbvF���      P��  ���y��	�3p�������ŋ�3
5gΜ���G�k�ܹQWW��Q����hmm��      �w   �Q����SN9%;�p�T��]�:th\t�E�U���);�P�?�xl۶-;      "�  �G�q�������7n�΀_���ƞ={�3
��ܜ�P��^xavF���      P���
;   lܸq�	�۲eK8p ;~EGGG,Z�(;�P���QWW��Qu���K�`Rggg̟??;     ��y�   �q�aÆ�xUe�R=|��8qbvF�)���5k�Ď;�3      ^a�   =�s��N(ܓO>�� �jŊ��֖�Q����߬A�ŤI��3
U�?     ��g�   =h����	�[�~}v�����X�`AvF��Νuuu�UcΜ9ѫW���tvv��3      ~��;   ��Q�F����3
���O=�Tv���]�5jT)�9^e�x�bŊؽ{wv     ��0p  �r��f'n�֭�o߾�xMk֬�;vdg���);�*0 &O���Q��=�     Tw   �!e����Of'�o��������(�[��섪0k֬�ӧOvFa:::bѢE�      ���   z�9眓�P����g'��*���1c�ĸq�3*^sssvB�|��سgOv     �o0p  �r��f'���N�����Ƕm۲3
U����jll��/�<;�Pe{�     ��   ��'�tRvF�:::bÆ�𺺺����5;�P��̙3�o߾��ioo�ŋgg      �*w   ��Ǐ�N(܆���������z��q�b�ر����);�PK�.�}��eg      �*w   ��~vB�{��x�֯_[�n��(T�F�oT�~�b�����*�     @u1p  �0q�����Sm�6�5puS�N�N8!;�0��K�fg      �&w   �fuuuq�y�eg����N�cR������G��Ψ8e�/^�8<��     ��  ���3&��Q��;wƶm۲3��lڴ)~�_dg�+��N�(�{���3gfg�lv      ���   ��ĉ�
�z;ժlc�9s�d'T�K/�4��Q�������˳3      ~+w   �f�~vB�y��8.��w_vB�.���2dHvF�hjj�N(ԢE����=;     �2p  �nv�d'���j���Ɔ�3
S__�f��Ψ���q�Wdg�l�X      T'w   �F}�����:+;�P��틍7fg�q+��lW�_�\'�tRvFa���+V���      x]�   Ѝ�=���ݻwvF�V�^����p��͛]]]����ˢ�����̙��P����Ǒ#G�3      ^��;   t�K.�$;�p�<�Hv�)/��B�[�.;�01}���t�g��N(T�ީ      �^�   Ѝ.�����SZ[[�
U�����ώSO=5;�0mmm�]     Tw   �&q�dg�����SOeg��6o޼�����(̌3���!;#M�����q����     �7��   ��E]}����(Ԛ5k�&�	;wk�fg������8�KMMM�	�jii�N      x��  ���q,���g'@�)��l#�_=zt�u�Y��ٱcG<���      o��;   tw�n��Ϗ�����̚5+����ǃs���N(Tkkk�~]     կ|�`  @8��c	��ڵkWlڴ);�M[[[�\�2;�0C����;/;�p�f��N(Լy�      ���;   t�K.��t��z�����΀n��Ғ�P��3gf'���q�fg��矏'�x";     ����w   �!S�L�N(��?�� �n��q�ȑ�m�>mڴ�ӧOvFaZZZ<�     Tw   �e�vuu�S����[�_��sN�|����)ۿ����     @m0p  �7�sΉѣGggjӦM�s����eO�>=;����1mڴ��<��3��SOeg      3w   x�f͚��P�2]��|-Z���(̌3�
q���ǐ!C�3
S�5     ��a�   o��ٳ�
�|����1(կ�)S�D�~��3z\Y�����ښ�      p\�  �M>|x�?>;�P�իWgg@�*���}�ƥ�^����fΜ��P��7�/~��     ��b�   o9s���.;�P?�p���gg@�Z�xq8p ;�0�>�9rd�u�Y��)�     @�1p  �7�+��N(���˳��:t(�.]��Q��3g���:����u����	      ���   �S����K.��(\�F��[��`����Z�P���_�>�nݚ�     p��  �8͙3'��铝Q��7Ƌ/����X�lY�۷/;�0�:�۷o\z���)Ӄ     @m2p  ���;��;�	�s��2ioo�x ;�0�:p��ˢ_�~���������     �7��   �ða���.��(ܲe˲�Pe��=q��:thvF������y��b۶m�      o��;   �+��2������^z)}���(�C=/��rvF!���cڴi�ݮN��Ld      ��\��  @7����������q����(TGGG,Z�(;�0ӧO�N�Vg�uV�5*;�����`���     �7��   �ј1cb	��[�pav�(�U�S��ԻS��z��իcǎ�      oZ�Z   �ꪫ�
w���X�rev�X�re�޽;;���'fgt�Z�H�۔�A     ���  �1����+��2;�p�/�����H���,��(L�\=?��.��(�ѣG��     P3�  �\r�%1f̘��NRve��]+WϧL���X�re���eg      tw   8������P�Ç���˳3 �ڵkcǎ��8��scȐ!�oZ�\�#��      P��  �6lX\q���[�|y<x0;RuvvFkkkvF!������/��x�j���FtttĢE��3      ���;   �A��{�}����(ܼy��"��Jv�_?;vl�r�)��X�|y�ٳ';     ���  �P__��{���Q�Ē%K�3�"�[�.�mۖ�Q�iӦE}}������ӳ
S�/     �r��W�   �@�f͊Q�Fegn�q�С��]]]�<8�=����V��ߨ���X�xqv     @�2p  �7�]�zWvB����g�	PQ�2p��ޑx߾}��/��(Ē%Kb����      ���   ^ǩ��S�L��(��ݻcŊ�PQ6l��7o��(D��'O�}����(D��      ���   ^�{��ި�/�o��͛����Pq�ϟ��P���??��q̪u��<˖-��      �v�{u   ���!C��o{vF���/;*RY�٨����w�(������fg      t;w   �-���D߾}�3
�e˖X�n]vT�͛7ǦM��3
Qmc�ѣGǘ1c�3
��ښ�      �#�  �5�p�	�w�+;#�]wݕ� ���%;�ӧO�����7l�̙�	�ؿ,_�<;     �G�  �kx׻����(�ѣG��{��΀�6o޼�B6,�>���7��.���F{{{v     @�0p  �Wѻw�x�{ޓ��bٲe�cǎ��h�>�l�_�>;��2ohh�I�&eg�,�       ���;   �����*F����⮻��N��P��q��'M�����=nϞ=�r���     �c�   ��W�^�G�G�)v��K�.�΀�0o޼������q]tQ�x����Z��o�����ȑ#�      =��   ~�����8�Ӳ3R�s�=��ё�U��_�u��eg��^�z�e�]���O���P���s      P^�   �444ğ�ɟdg������el\���G�cǎ���q�v�Gy$;     �G�  ���w�;F����bժU�y����*---��ٙ���*�:��3�
1��R�z     ���   �Cccc\{��i~��f'@�ٹsg�Y�&;�Ǎ1"�<����T��Kkkkv     @�3p  ��p��Ɛ!C�3R�����dg@Ujii�N(D�^q�ݻwL�<9;��m߾=}���     �g�   1x���k�3��y�q�����J,(�??S�N�NxU]tQ���?;�ǵ��Dgggv     @�3p  ����?��hll��H���?�я�3�j����ʕ+�3zܤI�*�ߓ�zY����      �  (�3�8#���weg�iii������je���'.�����0mڴ�����ǓO>��     Pw   J�ӟ�t���;;#��ߞ� Uo�q�ȑ�Wic�N:)ƍ�����͛]]]�      �0p  �Ԯ��ʊ�H\��<�x���z{�~8;��M�>=;�WL�>=���3z\�!      ���  (�~���7ܐ���{��^vԌ2��G���vZv�+*�|Ox�g��?�yv     @a�  (�|�q��'gg�y��bѢE�P3-Z����q�rŽ��>.���7o޼�     �B�  PJcƌ����:;#�w�������΀�q���X�lYvF�����^xa80;�ǵ��f'      ��  �ҩ���O����А�����-~�ӟfg@�iii�N�q�^zi���/;�b��=i�ƍ���Ogg      ��  ��y�;��_~yvF��o�=>��5gɒ%q��������&M��(���L      �:w   Je����},;#աC��;��΀�t�СX�dIvF��>}z��:th�s�9�Ehmm�N      (��;   �Q__7�tS466f�����㥗^�΀�U�����q��G}}m���O>[�n��      (\m�
   ������_������#����eg@M[�|y�۷/;�G�;6N>��ϟ=�/B�      x5�   ��g�����3��u�]���w��U��ǿ����p	� J		��4S��Y׵˓Vm����n��(�Zi��ljim覬UVE��Y�vj��5h���b���A�Sa0����lCM��!������zI�������x ��sOOO��h�|>6oޜ:�䚚��ܷ��&ٽGJ�P�����      I�  P�����G�����)I�ڵkSg@U��ӷS��o��Ƙ:uj�{��^x���     ��e�  @�{����[oM���3�<G�M�Ua۶m��k���(��������^����#��      o��  ���[��[����3��իW�΀�144mmm�3JjҤIq�M7��}������=G���p���     x+�   T�ٳg��?555�S�[�~���a�U�)�#=6�����K���=Gڮ]��ĉ�3      �1p  �"�7.����.Ə�:%����X�fM��:;w'O��(���/Y�$Ǝ;��i���     ��b�  @ũ����|�+1gΜ�)���(>�:����p�����(������~�]�x1���Rg      $e�  @���?����;RgdB>��U�V�΀�U�q�=:�.]:b������ۣ��/u     @R�   T����}q����Ȍ���q����P�v��ǎK�QR#5:�4iR̛7oD�J��!     ��0p  �b�z뭱r�ʨ��K��	����f͚�P�
�B�����(���755Emm��u�bӦM�3      ���  ��̜93���oŸq�R�d�ڵk���ө3��577�N(�n�!�N�Z���Ԑ>��{Ο�      a�  @�4iR<���1eʔ�)��ꫯ������@DtvvFwwwꌒ���������g$�R.�K�      �	�   ��1c������ǻ����)���SO���`�������N(�R��>gΜ���kKz����|lٲ%u     @&�  P�F����7bѢE�S2���+~���� ~A�������7jjjJv��n��d�΂���8{�l�     �L0p  �,�����?��~{��y��bhh(u�����J�Q2S�L�o��d�ojj*ٵ����9u     @f�  Pvjkk�G��éS2���%�oߞ:x�>b.�)�G��e˖���Y000[�nM�     ��   ��Q�F�ʕ+��~��R�d�������Rg obÆ�J����$�]�`A�7�$�΂���L�     ��   ��ѣG�ʕ+���S�d��ի���'u�&:L�Q2˖-�Q�F��+V�(�5�$�˥N      �w   ���ѣ��G�����L��IG����I���<f7n\̟?���-���Y���?��OSg      d��;   �w�UW�c�=f�����oE>�O���\.
�BꌒY�|yQ�7f̘X�paQ��%7n�g7     �/1p   �&N������}�{_��joo�͛7�� ކ���طo_ꌒ)��}ɒ%Q___�kfI%��     �N�  �Y�f͊U�V�ҥKS�d֙3g���F��2T�y���q�UW�z���E�V֜:u*v�ؑ:      s�  Ȥ�˗�?��?ǬY�R�d�7���8q�D��2lذ!
�Bꌒ����E��z�>>KZ[[chh(u     @��  �9w�yg<�����А:%�v���<�L��2?~<:;;Sg�L�F��ƍ�[n��(�ʢJ>�     �J�  �555q���W���=zt�L�������S���U�X����=1jԨ�\+kz{{c׮]�3      2��  �L�0aB�\�2>��ϧN)O<�D����� ޡ\.��é3Jb��1~��+�N���Y���R���      W��  ��,X���w��`ꔲ�k׮���:��|�w]]],]��S��J>�     �J�  ���>�������1cFꔲ����<��T�ȹ���^?q�Ę;wn�j�������/��      �,w   �7n\|��_��z(F��:�l����m����� ����5.^��:�$�����˗Gmme��e.��B��:      �*�_�   ȴ[n�%�~���Ї>�:����'?�6�� ��ԩS�cǎ�%q�M7ŤI������,���     ���  �SWW�����wb֬Y�s�Jwww<��c�3�"�Աsmmm,[����JO�Ϫ#G��޽{Sg      d��;   #b�ܹ�z�����c��ѩs��ŋ�_�j�N����-��|ꌒx���O�:5fϞ]�lذaC
��      �f�  @I�=:����<֮]��rKꜲ������ٙ:(�������H�QMMM��u���QSSS�lhnnN�      �y�   �̼y�bժU���1jԨ�9ei˖-���O�� J(�˥N(�ٳg�5�\sٯ[�lY	j�;t�P8p ���    IDATu     @��  Pt&L�/|��v�ڸ��S甭Ç��?��éS�ڴiS�?>uF����Dcc�e��=�yO	jҫ�72      ��;   ESSS��G�?�A|�3������Ie�����W�W��ߟ:(����غukꌒ�܁��ɓc���%�I���9u     @Y���  (����Ǘ���X�paꔊ�r��طo_�`��r���?�:��/_~Y�_�lY��Ԕ�&�DWWW�     ��`�  ��6mZ�w�}�|�"G�)�ۿ�[�_�>u0��n�1nܸ�)E5k֬�>}z���+o��˖-+qQ�\.u     @٨M   @y?~|�s�=�� >�я����?����Sg #lpp0���Sg�Dcc��~n��[ZZR'      �w   .�رc㮻����q�=��رcS'U��G�ƃ>CCC�S����S'����O�0!�Ν[⚑�gϞ8|�p�     ��1*u    �a�����<>�����ɓS�T�������'O�L�$��s�E444�N)�+V���-]�4jk+�<�\.�:     ���  �&O����'⮻�eVŃ>�J�$���c���������S�jƌ1cƌ���y��-[�l��FN�P�����      e��  �74����'>��������s*V�P��}�k�}���)@�r���GD,_�<��?��-�S��ݻw��a?      �g�  �%����;��;��O~2,X�:�*<��S�~���@Fl۶-���b��ɩS�����-�cƌ��o�y�FFsss�     ��c�  @,\�0����Ї>�s�����㩧�J�d�ŋc�ƍ�},uJQ�X��-��dɒ=z�Ռ����hkkK�     Pv� ��VWW/^L���5kV�q��|$�̙�:�괷��׾��(
�S����r7p�6mZ̚5+>��__�t����~��8q�D�     ��c�  \��|�+1eʔhnn��7��ӧS'�6�����;o�9uN�ڱcG<��C144�:Ƞ���g����\sMꔢjll|Ӂ��e�F������S'      �%w  �����m����v[<������---�q�����O��/����%K��o��o���������S'U�����җ��|>u
�Q��������ԧR���ŋ�?��?~�񺺺���[��ŋ���-u     @Y2p  �ȨQ����o��o�=����:^z�ضm[tttċ/�/^L�XufϞ˗/�+VĊ+���!u�����/|!R� ���\q�������͋�cǎpMiuttD___�     ��d�  Mmmm,Z�(-Zw�}w�={6v���k׮x��ދ���6n��X�xq,Y�$c��驳x?��������]��e������3f�H�R4�gώ���_�spѢE��J'�˥N      ([�  @Ɍ?>>���>����8w�\�۷/^z�K===�+�Gmmm���s�Ƽy��[n�E�ń	R��k9r$��~��o[�P�������?�:�hjjjb���ӟ��u�/X� QQi\�p!6mڔ:     �l�  #f�ر�t��X�t��������q�С�����ɓ'��7iҤ�7o^̝;�Ҡ��n�����i\�����q�}��+���:(3�\����{Z�/�+��g�}�w�      ��  @R�'O����hjjz�����������q���8v�X?~<�;===����UW]3f�x��u�]3f̈w��]1eʔԉ��/���w_����N�О={�ȑ#1s���)E3���}>q��x׻ޕ��4���S'      �5w   �b��űx��7��ɓ'����q�����닾�����S�N]��ٳg����q�ܹ*io}}}\}�՗>&N��~~��WǤI�.���+����������)@�*
����s��\ꔢ�馛^�����&QM�F{{{�     ��f�  ��)S�\�H<��ǹs��̙3q�̙��g�^���bpp�u�����q��EDĨQ�^��c�F���b̘1W��Dy饗�/��/���?u
P�*m�>mڴ�<y�7�,Z�(qQqmݺ5Rg      �5w  �*���G}}}L�81u
n�����/~�uo� x�8]]]1gΜ�)E3o޼��興�=����r��	      e�6u    T�͛7�<`�Usssꄢ�7o^DD�����������@lݺ5u     @�3p  �"��_��cpp0u
Pa*�T�{�7ZZZ"��ń	R�M{{{�?>u     @��:    �Y�P���z*�|���)@�:t�P<x0�Ν�:�(��룾�>uF�mذ!u     @Ep�;   �C/^�G}Ը(�J;Ž����Ƕm�Rg      Tw   x�/��/�G?�Q��
lذ!
�B��D[[[����      ��   .Swww�}����ϦN�đ#Gb�޽�3xN�     (w   �;w�?��?���N��u6�:u*v�ؑ:     �b�  �۴nݺ�������/u
P�r�\
������ָx�b�     ��1*u    d]>��G}4֯_�:�bǏ�_|1/^�:�_�d}     ��r�;   ���Ǐ��w�m�d�1u����Ʈ]�Rg      Tw   x�����O:��ݛ: ""���cxx8u�ǯ     @��  �/�����o~3|�����O�p�óŉ�      �g�   ����+>���������) oȨ:�?/��b�     ��c�   �g����'�'q����) o���5���RgT�6D�PH�     PqF�   �������_�zl޼9u
��u�ԩرcG�v�m�S����     J�	�   T�����뮻�ہ�b\�Vwww�۷/u     @E2p  �*���Ɨ���x衇���/u�eٸqc����U+��E�PH�     P��  �:---����֖:����m۶�ΨZN�     (�Q�   `����ģ�>j
T�\.���SgT�C����Sg      T,w   *ޅ�_��_cժUq�ܹ�9 E�iӦ8w�\�;6uJUٰaC�     ��V�:    Ji������~6�x�	�v���;w.�}���U���9u     @Es�;   ���;�x�hiiI�P2���q�w�Ψ���C���      �h�   T����x��c͚5���S� �T{{{�={6Ə�:�*�r��	      �6u    ���p<��3��O~2�|�I�v�*���زeKꌪỂ      ���  ({���ǁR� ��\.���SgT�������N�     P��  ([�w�'�x"����) �<��sq�����S�T�����	      U��  ���gϞ��w����S ��p�Bl޼9����)�P(Dkkk�     ��`�  @����5k���͛�P(��Ȍ\.g�^B�w�cǎ��      �
�   d��ݻc�ڵNlx����'ON�R�r�\�     ��a�  @&
�غuk�Z�*:;;S� d�ŋ���->��N�8��ñq���      U��  �L�p�B�r�X�fMtuu��(�\���v��'N�H�     P5�  Ȅ���x�g������W^I�Pvv��'N��iӦ�N�(�\.u     @U1p   ��{������ذaC��([��������ԧR�T����hkkK�     PU�  q�|>������ntvv����\����:::��^K�     PU�  1{���'�_��_q����9 �^�����1cFꔊ���R'      Tw   J���?���cݺu�w���9 �P(Dkkk|�3�I�R���|lڴ)u     @�1p  �膇�cǎ�nݺؼys\�p!u@���r�E��s�ř3gRg      Tw   �bhh(v��7n�������K�P������Y�f�N)k�\.u     @U2p  �;�|l߾=������=���S'������>uF��-[���      �J�   \����ؼyslܸ1�o��|>u �$���_�-[����@�     ��d�  �[�^x!:::���#�����é� x�����3gNꔲ���R'      T-w   ^gxx8���i�����;��577�=�ܓ:��ĳ�>�:     �j�  ���_����hhhH�B���k���{�����ؽ{w���
=����O��      ��b�  \�իW��իc�̙���MMM����&MJ�Ư144���>v��{���(
��        � �w�ȑ#�nݺX�n]������_s�΍o�1�̙s�΍�3gFmmm�Ԫt�ر�����������8p�@<x0���R�       �!w  �(
�BtuuEWWW�r�K����ǜ9s��믏�3gƌ3�뮻�c}}}���7<<'N��C�]����gϞM�       pY� �����o߾طo߯|���&��暘1cF\{�1u��_��6mZ444$(φB����j=z4�====��8v�X\�p!u&       @Q�  ���x��W_�_|�M�W__ӧO��S��u�]ӦM��ӧ����cڴiq��FCCC�3f�L___�:u*������7������/N�<'O�����'"�ϧ�       �  @����������|^}}}444\���ꫣ��!Ǝ{�����:"�W>������q�ƽi����_������/\��Ν�����s��Źs��̙3100p�3g��ٳgcxx����        �`�  @�����������S        xjS           @��;           a�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;           �`�          @&�          �	�           d��;          �?�ڱ    � �i�(�`Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap       $?-    IDAT   `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap     b׎    �[OcGq     �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;        ���    IDAT   �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;�v,    0��z;�#          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�       v�X    `���4vG   ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���       ���    IDAT   ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���  �k�    ������8        w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w         b�j   �]� �=Z0 ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��       7���    IDAT   ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H8���  ��޽�ؙ���>�sΙ�w�	��z4iA�/�QĦ
�UB��B �\SJQ�H[�Tĭ�P!�i�E�Ti
�%$Q����,�sfl�q�B��g��ˎ=��\~�#;��k��ޙ��3�zI�g������s~     ��(
�  �CʈX�        ױ�;   �9eD��        �kI)ٶ  �b�       ��*�b=w  �s�       [Np ����       �q��;   �9�        �-'� ��R�W�       0�ʲ4p �=���s�#        �Z��{<w  �sʈ8�;        �%�d�  {HK�#        �Z��3p �=�	�        ��f~~���  ��)��        cj)"��  ��q�;        �ʮ  �'�       0��Z  `�)���"b-w        \�(����   �2"���\�        x���   vV�R�l�m��N        �3�y�Q���;  �1�S��       �A��h���  ��2"�,ˇs�lX__ϝ        �g����N��+sss_�  �2"���O�ٰ���;       `OH)����3�rG   ;���h���1&��h��        v�+W�D�u�3��3�  ��WFD,..^I)]����ŋ��X��       v��R\�t)wƳ9�;   �y��m�~!g��F�Q,//��        ص.\�m��θ��,?��  �y�U��C�ŋcmm-w       ��s�ʕ�|�r�g�^�|���  �����z���3�ZΝ;u]��        �5�������3�ˉ�'O��  ������,��r�<]�u���d�       ��������1��<CJ���  @�����:�4v/�������N       �XW�\��q{DDQ�n   �(�����\!Ϧ�8w�\,//�N       �()��p�B<��1n�����  �<�l�^U����\6�Ν;]���       {m��c�=6i�
>177���  @O��ψ�ꮬ���ӧcuu5w
       �غ|�r�9s&���s�ܬ�Ř�W  ���e�x�ɶm�犹Q]���?�Ν��ms�        ����cii)Ο?]��ιiEQ|4w  �O��/�m�@��[�q���K�"%/�       �����q���I<�}C��?�  ��{�F��o�7刹)��t�R,//�^����;�(��Y        ;��X^^����<��jm�^|衇�"w  ��3Np?u��'"����t]�.]�G}ԉ�       �����8}�t\�ti���]�-�n   �z�	�����|������o���q�w���e��?       �Dj�6������˻b�~���ޓ�  ��Z��4�>��%[�뺸x�b<��q�ܹX[[˝       p�����ܹsq���x��'wݸ=�Ծ�e/���  @^ŵ�v���/}鉸� ~[�߿?��ZY��`0��o�=n��m��w����F�3       ����;�3wƞ�R�+W����r�u�-��.VWW���ϥ���`0�����O��CYB  ��ѻ����˗?]��SJ/��m4�����q��Ÿ����n�|H       kkkq�ʕXYY��R�m1���o~�RzO�  `L\k��~��#��w��]����r,//GUU��~cw        ����ʕ+q�ʕh�6wζ)�"�A�z=[I)5��1  ����E/������LMM����w�iG�m�9v����c���        �C]ױ��+++Q�u�mw�q{DD�4s��  ��uW���w_333��^�ޢ(b}}}׾�Ն���ҥKq�ҥ��z�o߾طo_LMMEQ��       �]`}}=VWWcuuuO��7E���Q��3~��_Ȑ  ��g=��,˟��?��*������}C�4�'��e��ӱo߾ؿ��;       pú������Q{��ʟcܾ�����Y  �zց����GgggW˲�WUULOO���ڞ�o�n���Ο?SSS�'���y       �I)�h4���F��IYm,x����og�  �q����躮��eY�5�K������h�v��OJ)���bmm-"��{2bzz:����      `����������<��Zz�^���#"��{�&  c��?�R���'�����FQ��6獿���z�>==SSS1==�~?s!       ��RJQ�u���o��ڿ\Q����s7�4�#�P  0�s�>??���c�NVU����>���X__����N���bee%VVV"�K��~���`s�^�e�J       �F�m��(F���	��W������v�   ��FNp���OD�G�����b߾}1��i�-�����|�]^^���~���������~���o�       쌔��}���msgM��Mč� ��[������  &�����?z�رUU}���(�����^����[n݀�i�i��Sދ��^����\�w'�      ���.��<�}4E]׹�&RY�7�u���w"�Q�  �����{DDJ��"�]�����뺎����MH)m��]�������~�z7��       �/��|�4��;���+�"��M�RJ�;���m�  &�?]LOO�\]���(������v]��4����жm��������׊����6O{��ۍ��       �VW�7�m|n����~��[�+4M�ɏ���!  �p7<p����W�;������~�ƫs������xo��ˆ������﫪�T       [+�m�nׯ��m�;o�+�bs��|�K)}�f  ��M�?T�4?R��wEqC�髇�^��6��O�q�{��{�7'�      0n�>b��7Mm��d�U�����iޢ4  `�������╣G�~����Û�uW?��ＫO}���,7�C���6?.��      �-�1^��o|��y�4�u]�L�����UU���\  ؕnj���L)}[Q�����~���
kC������h���?������UUm��˲4�      ��RJ�u��X��7����cc������u]?<���  ��r���px�رc������C���=�����tx�|ėp7��W�૪��      `�5M����u�5���Mxw(�r�����R��(~x�/  �*��4�R�ޔ��[9���^�z�͡;�m�/2       �]����l�9l�ж����?ٶ   ��-������[���b߾}Q�V^       �gQ�e�۷o[��O���  0�n��������K�       xVu]?0??��;  ��w������woe        �K�u)���;  ��P<�__���^,��[R       ��R�����?��  L�[>��)]�u?�%%        �*]�Տ=�����   &�������o�m����       `�h��O�>���  ��{�QUշGDڊk       0���9����ӹ;  �ɲ%�|���m?��       `W���  ��ْ�{DēO>�]׭n��        �L�������$w  0y�l�~�ԩ�����V]       ���u�������  �dڲ�{D����o�u}b+�	       ��h����O�^��  L�-�GDLMM���R���       `��m{b8�'w  0����࣏>z����,��o��       O)��,˙ӧO_��  L�b�.|�ر�TU�u�u}        ������Z\\��;  ��Vnׅ��xmJ�ޮ�       0��Y0n  �¶�����5M���u}        �k�v�R���;  ��a�����M�ܷ��         ���Ë�#  ��a[������uݓ�}        vV]׿��C}0w  �{l���ԩS�)�7���v�       ���4��p8���  ��R��MΜ9���ʲ|�N�       ��Rj��9���t!w  ��;y�����{�޽;yO        �NJ)����v������  �>�N�셦�c�  ZIDAT/|�7�m{n'�	       ��i��}��  �v���#"fff�VY��ʲ����       �uM�|j~~�`�  `����#"�����(����}       �um�^^ZZzu�  `w�r����ӟ��{�.��C       ��K)�]�����}[  �ݭ�y󙙙?��z���        ����R�4o����  �~Y�Q���|���}m�        �&�u]�������  ����O���Gڶ���       �������� ����������}ID|�,���-        D�F����  �-�Op������3)�צ���-        {]�4_XXX�;�;  ��g,�=��\]�oI)��-        {U�4�۶����r�   {O�;�jKKK���{>S��GD��       `/i�������~�ӟ���  ؛�j�q�̙���s�٢(�\��;       ��n%��O}�SK�[  ��k��gΜ��뮻���ꍹ[        v��mך�9������-  ��6�������O�u�]eUUߔ�       `��n3���s�[   �v����t��w��/��uEQ��       �Uڶu]����'r�   D���="��ٳ|�wֽ^�s�        �mۮ�m;���p<w  ����GD,--��+��M�(w       ��m���h���Ǐ6w  ��&b�q���??p�������(��       nA۶OE񊅅����  �t7�������>PE��       `�4M�D�4_{����[   �e��G�ym����,��[        &A�4u��{�G�r�   \�D�#"�;��EQ<X��m�[        �Y]����XDt�[   �M�;�V=��C�n�����9��       `�������Gø  � ;p���_��u�4�s�        ��T����÷�  �QEr�ȑ����       �[�u�h4���Ǐ�?w  �ͨrl�����=p��zQ�\Ů�       ܌�mW���w~~�c�[   n֮�9r��^�CeYr�        줦i�P�塹��K�[   nŮ�GD��U�:�����^��-        ;�����o��  �|�ʁ�S������z�o�       �]ڶ횦y������  �|U���ٳg���w?^��EQ��       �Jm�>�0� w  �V��'�o���=/���-        [a4�r�ʫO�:���  `�쉁{D���l�i�?ߘ�       �Vu]׵m�����gr�   l�=3p�033�ceY�JY�U�       ���4ͅ�x����B�  �������/i����~�e�[        �KJ)F��Gߜ�  `;�Ɂ�����wWU���(���       0�ڶ]m�歋����  `���a��Ç���z���E�[        �6�>q�ҥ�?��#k�[   v�?�8|��o��s�;       �[۶�m������o�n  �Ie�1����CM�|1w       �7��b4��^h�  �EN+��#G��l����eYV�[       ���m�'�~����?��   �똝�}i۶������       �^]ץ�i޿���[   r3pG���EQ�Z�׻=w       ��4M�HD�y~~�S�[   Ɓ���)�=��UU��,�2w       0ٚ��ܶ��ߗ�  `��߄��������L�       `�ں�߷���O""��  7��ȑ#o(���z��s�        �/�u]?����unn�\�  �qe��<=z�G���Ų,���       ��������N�<���-   ���}>|�]�~��ʲ���       ����k��m'N��p�  �Ia�u�Ç�����PY���1       @M�\�F�8y����  0iܷ������W�����(z�{       ���4͓u]��'ޝ�  `R�o������TU�O˲��       �G]�RJ?����s�   L:��W:t�����TU�?w       �5�>�Rz����r�   ��;�СCo��z?������       ܼ�R4M����yǉ'>��  `�1p�����o-������r�        ϭ뺮��������}&w  �ne������+��{OUU�TE��       �rmۮ4M�����?v�}����  ����Cy���wVU��^��1       �����i�G����'O�7w  �^b�>f�9�(~���*����       {E۶km�~���}nn�L�  ����}L<xpPUջ���g�^�%�{       `7�.�m{�m�w������  ���'�k^�Z]]���,�AUU/��       �����{u]��ɓ'/��  �K�'�ѣG�?Y��lUU��=       0)����u��)��_��Gr�   �L���ѣo*��_EqoUU�s�       �8I)E�4SJ���y�����   xv�ġC�^W��ʲ|m�׻=w       �R��m���#EQ����  &���.t�ȑWD�O�e�Ʋ,��,�2w       l����i>�4�����~�������   �5�_y�Сﯪ���8���^�;       ���Rj��\�u�iqq�s7  �5������;��{GJ��eY�����r7      ���.u]w�뺓)��[YY��S�N���  `���q|qD�P��sQ˲|qY��\       �M�u]۶�RJÔ��,..�/"��]   l?Cf��[�������]EQ��,˿Y�����G      �����엺�����'ڶ�o'O��x�.   �Z�9]5zsY�����)��EeY���       �]�5m�^H)�EJ�]�}�ĉ��  ��a��-{�k^�U+++oL)�[�+�����,�FY�Ӆ#�      ����RJi��'#�/��F��m��C'O�<��  ��f�̶���}e]ׯ/��p|������;#�UUME�˜      �MJ)E�uMJi���)�sEQ|1��ٶm����~��Gsw  0���fvv�ow]w�뺗��^w�e��(nO)�Vž��*˲�R�GD��8�z��"�TED
�      ��(�H)u�w]�E���uD�)���XI)].�b����/��Δe�Ţ(>�u݃����e�O   `��QO-�evmu    IEND�B`�PK
     ˡ�Z����J  J  /   images/1251016d-b52c-4e05-b483-3027638d0c75.png�PNG

   IHDR   d   �   �|�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��]	p��~w�O6		�����5��P�0i���֪E���
�Z;����^���Q�B	�%2�.�}���9�dw�G����[���@���|��������>�{�d�� F������҅��۷�ڦM�_'''w���im�X�x5m�YjX�UUUy�.]�\QQ����<�;v,j1���x���|�G��Сy<��|���b�Z�vF��9������?>�m����5��ā���Ƞ���цaЉ'�ܹs�����!55�n��6Lл&&$�}�ҥ\2	�a�F:&Ҕ�Q�B���n����3��p�������r������.2�p�\f)c)d9�r��h�(�\���%ƨ��cFH���
�,_�.��]=��r�eK6�7,|����S��$�! �=�	1r�t��OT'ڰ�K,�X>a���ܩ>V�FMMi���u�U���d��H߇/����(Y�ci, �q�\�f��>!�7������yV�����N�ϝx�,]XҮ>Mo�y,`Y��w�=��۱�&B���������T���q���jN����������[�nMii����˩��T(�f�	E�>���$>#K+**"N!��p�ڰa�̼��N��x_���±�=jԨ�:uz	J�׍IRy�XX��0�p>$3�������W���gN��s觟zS�^��i�[����X���?=�4�q,C�Ә�ʄ,�����,o�l"3A0�Zk<!B0pؾ���ɓ郞���ӿlNsM2�˛Wj�Bdf.�M &11�Z�j%���3���v��Ἕ4�ot9�����gV�^��Q_>hҤI������\�k�D!��	%ƅ1��p�ǃ�G]�t��q��o�.�w۽�~չs�:����X�8������A�4J�}֏��}��@i������d�6����.]�T�gtVv�x�A)))W�
��iٲ� ��c#�.�����E�pX�?rܸq���Nz��g�Iƒ%Khڴi�m۶>�4�����EN$�T��0&�o�ڵt����υ�$Y�C��ŰH����̙3��N�Jo���5Ǖo���i��,����4��,��)�M��uWء}�2�n)��"�ٛ�8���mۖ�22z��EG�!.�%��$rf���S�N�j�`&�g#�!ҧO:t�PO(v�ƍT_@�,�`�C�%�[�|���a7�I1�j�8|�w/^�bK����X�<�v����}�>�57��?��G��ÎM	J��ġcǎX���Ç��c&E*qCP2nĀ ̾H�A�P�ҹw���EbO΁��UZFm��O�OƉH�����/��,2g�k���X��ƽH����j2� X�X�jԖj����WPVV�4N��@����������D���}�î���w��A�Sp=� R�����.RZUȽFr��a�|����[j �Df!9?�����l)�n���5�dZF砠�A ���dG���?���"����ᆥ��{�A �qr?�,H(((�O�\�L��W(����8�����w���+\W�@-�	�={V�	|O�%�=�ڷo�X�6(mq�s�F'���D�bCp%A�	?�*B�a�2�"e�1@��W�9�d �w�!�/��h�kٴiΑ�n�:/bT}�ka2�yr����l%���Z]�-1��ŬG|C�UW=�	F9�o[�X�P'"����j�e��I,+ȬG^���
�ib�xauJ�%W��=[鴣3�ew�$�<����Y�j�8D<P����>�v_&GY[����|V�-��A�GP��>W�� U8��]�ߑ��M#gi���}{�-�s[��5�3�3:MO�u<~fj�tg�)��� ���@�NS�/�v�-*�}_�GU�aM���İ������"���m?�l��'�6/83.���{jF�a�Ѿ��Ǿ?�E���i�W]/)�d)f�w��i2c�B2+�b���"F�t;y؃�&٩�ԑ�͞�#�W0���a$��l���}9����j	���?���I0G����Y>��\���#����믲�>��}��%-ƙF)兔WJ,�6�9�ƃz���ے,I�ʸ`���K	��Z�)��O<䭎�ώ�ؗS=��i��'&��?`ْ�!���'Ҟ�?��Ezh�����d>:�����dZ��,[Y8;����U^��^������$������9�NwP��<�	���Y��>�ԇ��wV[B�JUU#�pIAB[dZ�5�K���<f��h��)�]ik_?�XvN����f��&�����Y�����^��v#Y1�'Q��g\(nZ�#��eP �5��[��fOi�ވK2�հ���_�Qssp���i�0�e�	i����]ra���mi����/U�nt��'sɴ���t��d�jð،��q-�8�˸`d��)/��,�÷&�b���b��l	��:˟�tVg�v7���Y�!���X~�2�%��%K��t{{�9I�T	�CQ\5?B�$A�K'".��rs����n(!2�����	d�X���C��b$t�A����j/�9g	4��

.O�Ŋ&栆3D�$��4�匀��z!�lD��f'n��Q���Q�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�c%��Y���?��{����_5ZXVYl���+����g�]T���Џ"�����z�Y�����EV��<|~g%�X�h�f|�M	u,J�	� !*�XLn��9�^G���}���������S�K���%
ð�9�:mV��4Q���vL��w�B'��e,A�Dkv�^�����&D1hB�&D1hB�&D1hBC�		��TS�D�����J	��hj�p8D4M�����fh29c�3f����9ڪU���w�����ۜ���=��ۢE�h���*6l� ,b��ᄶ�h�9gΜ[�E��@�����<� m g͚%:^����x�b=z4}��W�r�Jф��K1�j�~+�Q	���(n
X�l�V|@~~>͟?_��ɓ'Ӛ5kB=e�ٺz Jk�n�&�J��Ѩ�@����n�'O��K%`hˊ�={���P�>(�Y�_�^����$���*��׏^�uaa��ܪht��
���g�ޣ�(ڸv��U�lr_�?.��O�0���}A���@:c�;6�y��$�J�l1�޸�!��
�g�baA K�� [�b�ѣG����ۗ�@��͛E�` Y�=��#���_�DA~w��Q	��ѤM�G�A'N��e�~��w��/�4x˖-��~��$l�ȑ���T�:�>).bb�Ν;E�Fv5d��u�X���.��ر�fΜ)����5$bU������rϞ=������(��矧ٳg�l
�z�͛G�=�� �L����p����A�8/���1M�]Q�d?p- �``�t���Q�̝;W�X��/2��8��uC`9M�]Q{�R�r0�e��l��A��x�gKP>�W��B�ׅc@�޽{�������?�V@&�F(٘������n �<�n��v�*�pQȮ�,,|����>��e�6��L�"�2FZ�\���Ͻ ��M�	qT	��a + L�>]��p�B�T����Q����c��"x����H�ہ�X�
�
@ 1�/_^�c(�� !@v�X�BdhM�]�N�tQ[�n��P�c[^^� �ZOl�y��HΕ���$���]��C�I����SC`�������g�	i �$4U������&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB�&D1hB� �Z�ljDEIF ��$)X�S�V(Ū� ����k�E����*�X��7wR�� ˊc�^~�g=�Ƶ�����<��2)�J Lsuc������*׀�n�������pYkY�����X��e��NʏX��:�Xӽ�!������fǒ�b��J2��vU+d������|�����    IEND�B`�PK 
     ˡ�Z�`�* *                  cirkitFile.jsonPK 
     ˡ�Z                        =* jsons/PK 
     ˡ�Z1٭<7  <7               a* jsons/user_defined.jsonPK 
     ˡ�Z                        �a images/PK 
     ˡ�Z��7��$ �$ /             �a images/e575fc9c-d7f1-4841-924b-9061a1257de8.pngPK 
     ˡ�Z�C��R  R  /             ͆ images/b905cced-8669-4310-a345-cc026e3fb08c.pngPK 
     ˡ�Z`$[ [ /             l� images/dd9bac2c-35cc-4be2-808f-eb026b88f611.pngPK 
     ˡ�Z�+�sz;  z;  /             �
 images/a657ee5f-a898-4bcf-bee9-a045b7cf922a.pngPK 
     ˡ�Z�v %� %� /             ��
 images/dfc5a72c-0224-4495-b3b7-0d06b4ba9157.pngPK 
     ˡ�Zp�"^��  ��  /             M� images/f159b6d4-7cee-4dce-98d3-76d280a06797.pngPK 
     ˡ�Z��n GV GV /             ;, images/5a738b76-89aa-4728-b8e5-f09c859dbb14.pngPK 
     ˡ�Z����C   C   /             ς images/ba153158-cccd-4fb1-9320-38bebad1b7f9.pngPK 
     ˡ�ZM8��! �! /             _� images/53de2a41-b288-4dfc-9a43-3e5c75810bf2.pngPK 
     ˡ�Z,�ln/  n/  /             ��0 images/6590c6c2-4084-4043-8677-a67706af7572.pngPK 
     ˡ�ZI�)�V�  V�  /             C�0 images/f2dbd413-946a-4dd4-beb8-9b389826ae17.pngPK 
     ˡ�Z,*��  �  /             �1 images/685e2fcc-e73c-46e4-a7b3-171ef11b9715.pngPK 
     ˡ�Z>zG�  G�  /             �1 images/7485d96b-ebc9-4409-ad2f-5f0bda14de1d.pngPK 
     ˡ�Z��)��7  �7  /             �u2 images/544a1249-aa5b-4970-8b42-188baf88f36b.pngPK 
     ˡ�Z~��ٮ ٮ /             ȭ2 images/2cd57c9b-7217-4a6b-8577-1769ce4bee7a.pngPK 
     ˡ�Z����J  J  /             �\5 images/1251016d-b52c-4e05-b483-3027638d0c75.pngPK      �  �n5   